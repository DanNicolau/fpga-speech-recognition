`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EErsftIDJVF0m0AzARUB1bTNfa1D65PKFzXVCO3IcVnfdNzarCrieLdbzQivIMAadZGQICQFGhS1
QckM881Qig==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oVVLyVCgNzQviLS1eG+3q0tFr/JK9RCUE5+xAA69a5PzCR+NN1kdZCFY3Hih5lupWCZCqlSR2yxj
T/gFuX/P5PwLJG5+6QmvoI5i4SAxY/rHrl8XM8Kicu6z19CTYp1SPiJ9834l0f0lOlXlTmn836kA
Wgmrcs24F99177fCyOw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kW4owDNqb8AMzEcxlafWfz8koQuLn9mxd/TVVOMuiv8YQ3rvx8K/DGu+WboW7BU9KyEVtBG1MjQH
gJKixZB+7AY25kT/0NwJhM5YyjG4KdEl5DSZuDhsBJip1w/5m+kP4N5/vcsnGSfB2gcc5U+hEZN2
tOLv961hH8596MgBAeOrfvnWa5SH9SROtve5GcJIcP2+J4rtDHR6wFKwG2xp/9kU818nQ53uY3x/
7USyyE73h57I6tiR1+FD47Z14CKQGy+J0+yoYnuxOAdrlqmEtQAPiwIuHmV0R7zwgIucScma6/i1
zxERzOQ0UeBZqrcJuNAcQN3PnQ03sEWGfc4Qwg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iAL6wKTA9iQaAsMi/04OqmErqGG219F3T4DtEhjCOkAVV5xns/q62D9v80Yu9LkL7GOPStNaimH0
0fLZZNbLN9aXY+LXsOjLmXKIRD1NJHFD/6y4EmfJhRxv4wTaSxMi35TYjtTPOpBQ9f3kiGqvET6q
oTK12b3zP6bRyeM2ZbhHWjG88vLFxPuV0/g08KIWxnwsizoJce9xWIbPH46yn/atycdYeI6hNlt4
AsWLZjzzPTaNgwoNSmXe6Z/iHwOsFgDluZ4wunNLVxH5Ru3KpxGf9jGPoEfbj76tqe2kxC3Whmb2
TOD3EfgrtAPEX3iiwhkJ68FGwrBXobVCgJLrLQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AYk0GVXSV/oBWSOxjuGlD2oLlqIfBX5t16vozwXg1+siZJZSMUHEbzptzgNoTGyAuDaMihDY3BLO
EtrWbX/36HzF6OYvwf5POdt/VXMiD/WmbkoqBGEm8hBrg/s//Xc8uwTP0aCjxNObZuBko/Q25mgQ
30NgIumW8FqCkhPd5zaKXjVEqWRkZbVy3s9drUMCg7SmsRWiURkSk2U7gJHgxqNeqEvn/U3HMsD5
przVbreKAnJv/RzsnAueSJ7se+zz3ea7TcdOm8FG4lJPtFHb6jvhIcFQ6qftny2xQ/73EGrSBx8k
emkzKeZp3UgSKQV+dZEMJkjg6+hPhExCSG3ddw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z2aYnMPHx9JY2YhtHwU80KMSOWZwPC6TzLQf1GQQ4Vnr361DuLoPMu0MbOnkBR90QGDH/qF7P5Cr
Ly2yiYO0/eJzmgzCpSyJ27rzee68zFBRRDPmlOAN8FHZvnbWm8t3N4kjdk2vzG0NcvKGeDmWVBg8
WX1YKAu49GjIv50pk7s=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZhLzhPI8pgMrQMSYddC1+njODiKwQHec1wBB4U5W8/l4gRoB3jhisEMfFb5EoL+ePeazVA8YvpBO
fy15vYUdxOsCKx+vVBouvB0iJLQJ7MJ2yB0Atezf8W/dnulTtecMT4xYThtmLmUoLpjc/XY+sv5+
kYuBtkUrJcr6xJNsQtV8JIkAU/9rh0McphkltAYVfKvFQQ4iPL6Vn52nStdWLo/EzZRGxkA2w3hx
RxGGI0fCa662AzFgfo3+9jW4FVA/MfRfrEnMa/qSzvX29NQHmhsMx87TbESpFUhf8rcOf4pNxnvZ
Kz+Rm+SekS5sOFDAnkaGJ2fOU9v6YhYC3w3/eA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
NW4pcXfCDnY7e8k9fHdc6LAwfVsGJvenMY/dzHa3l7e+U7QmEIbgbOTODRZKY/v7qBjw16A5CEGc
HlzdUvX2icSI5EZaUDvJCMukOfxrq4qNPwdI5pdxKyyjT5f0bMgLU8WQt+WktBnP6jYkVatkyreY
+UQs690Ym7ZU1+9qxo12s9VLLx6b6+mO0WiMaF7BJAKKi2+HFX0Y2KH3ZMi9qNih43gpjC4LhWdk
9G5lXKmc0P7YJL9GQO2QBMvqF7pBE+PESRPQp8VurByWi9UKP/J9EDq2lVmOAh7zBu8v87u0Qhjz
WEgzZ5XtP0OaTEf80PEjXwk/U+dHLiG5rh0k1BhapUqA62urdZE/V9SVjo8ZxUYMoUTkbpv4zfq5
wmykcRzdDBE3ai01Zxwgb31h2Fs1mG0P6Q5M1wDd8GE93IHIgC4rF3yNKzEK1GM5LUZbywzL2LN5
Cbvb4d+arwmvEQKwZO6o96FsLGPtGrxfO+jf2z1jLR3bTCoSJH4E45FEDD1PX/xdcZCQhX1wH9jo
m4cnVg5lMJFUMoD00RJWi2jLk/39jDKnqeEvFDA+1ZMlBVP/LOdSNs30ncmflGlp6WVDxoGJdh23
hY5ES9Cybw3ozSaj8aQ1M6F5GX57fLxLm+OjR7ci72Lm/5SNYJ9tqC6SU+bNYic7ZorImgHC4ljP
JUYVyzvguzRU0Dv/fx252VagQ49WL8V7aU+HISIxRTVsbhej/EPNQsSEhrdqC9njRtD2NsXsHJMd
XS8EW56hohlsirTbgP8BDzESLd8bKi/h9KpwPgzMeum8j98PQkRLjp7JlO4w8dZAdD5WIIKC7HFf
xCsP4qwfVVfmOWiZ+oHIrY1vyOuEq6YAOXpgDSK2YO+xFWWO9zkkiwDmmQTraHD1ptF/Hk08Wfa9
8w25RAwGxumXHReGFOoKv9/U2xGYN92KazY/YaIxgiXeI3CQrbYrLkjP9MYI3bJGPMnrckjZg1UY
w5mrXkOP3BxCRad8w1qQg/imiCQVBBCXzCdNxBocY3QqfpMZx90ZbsRc1jZJ1Ax+O/7ehuSiNXlG
4ezTRnSNdzuBVAkE5tOsn5HP2YAOu4O71ABU2qhcXpSUZvSPTyotdnTTmxLgVMnogRxyidV2RKuG
2JzewqYMktk1AFHZeXjLlI01XU3YY91NVaML73/FuROJPuyjXQg9/3nRrX9upZg0YVUzFjD5WorQ
FQj1FDax7kF6NmIldsbiINr668gUYi4qLtzM9ttCj1cjfOebPSflOtatyksCF6PV47PEc7Z5EuXl
an/JLNUiissGSVjDiSxrCs2P7jzAQp+QxrLDw6nHd4AvgeUFcDFnPIuX+BeN/wdQgQhN//yxMTXo
7HGlLK7JzkLWkEjlImEp0k6DLg9fsxrLNk0+Txkn0EQwTl4DZlMAWEYqQswhqahEcaJLvWq8P4Bq
8qX7iPuHtFF5iq6BoXfEQ4CB6dgx7O0wcYAvFHlMWugJ4E4U+pgJwLrGgA6dh9cQNh0SNoS4+u4p
0xWsT5jpvcleVbJ08TkdP3/pAzr+sorrgZ+yC2tuCvJW+TCqXgz+y2Dyjz1VOgYsn0Tv8KQzD4dI
gp+mDInhnYXxzcYiXCch9fCXAjJ6BQzxgLE1QDKvpnM7Q4v25dx0edzOSOTqx4A6vU7BMF2t92IC
Belo4DlTlzWL5IXaO2vsdpVPJOd9O3m/edKpgrtrVmlKHHohrwhxgANQr8twwa8LDpOf3MXylLbe
wBlj0yCvkNEMxfm0OR/sivs3yJx1M9ggGXuK4uqbExfuBk8ZI7cCxtZI7nRdKmr4Ssv5rgn2SHxe
m5FKRw76EProB9t1kHy0MM8khcQxQi2cWtcmyh9sUAGMmX8CmnykuAhxQW1To0k3C4U0Dd4jsBqI
yWC3WsoEdu/icqpEl+BLYeja1GVWYs576CayVAHAyNxhxHeC2UDWcmWIJwt7HwMocXu77s5EAQd6
1BIo+W6/8WRLNH64Cq2edvHFdqLHZjM81sEkuv0d9HC15QqOI/XXGi/Uw+AgzfltTaqmhhZ1dmqX
XRtcy3nqpE9Pgk6UPvZ22z1CMu79iF0PDTVqooV+uQ+Gouik2ajHch7/hGbhMpGLOGR/mzMv12eb
J/udxWJw785QKQerPPMvAq195mhxEMnWC3MlQnFqn3nrEB7RIjBTgmNOBm0JGTKiysnTOVlEvm6w
aVSyJZXgqef1KTDSvSWV9kk9Lea8M4T3I8GwWdQqQlOSabT5HYSKvSTPRVhtApSJn7FfRxhkEy4T
I2T05qYD0sbQPL6L05i5DNAokJTy8PHQKstzlgja+X5OgnBceCDAxyS/I0fTFymHElOvsGhPdTFB
itjnC9vUpczOyqdGXjlwoTpY2o9iHPGcYsvS+B+yHR3siYnd7dyMYnNBa8q5UTDWZcqd29nXpJ9/
PWQb3rniG6AdxcYV4GK3uh3q+p1FhvVy/i4x0iSpJrR+LdSbH7R84QpQZ0t6PkDxZsvhGxvBeriH
S/gEfpoo1zLdUWt9xO+GIi8UPtZ0A9xOC8EhjHvQIlQuIsoCst3cegAMRHyfIq11eOz1M+ugE6X4
bjQgWFkqPw8bw7DTm9CBh5eHo8wqxImpBqSlFW0V3hc2RFjIFSSMvPeyNRr/WSg9nsQXLSn7r4/A
aG69V4KB3V97GPPgBr3/TsY+LtgE3p118p0cA57Tm+3C88QgeO0yqBUsH0P3P9zq8b1E05dBId+N
7LT4io/SlP86RA3sDmELEdn9HEdiqst8eFlFJ1sqQj2MRACxLRzN1lB3TZEtaYtkMg8H69XQ1QZX
iPJkk3YRdPzUXiaoU5lt4XFiTxf62xkJvCwnZgMKK3l/0aKhbXkD65G5sPU6c4C7Z4qPxyASgeMJ
3enhkPNmeP4u+hTUMuUF255pFJMt3tphqv5OMlV7Q1LgwEhmXyjdTihc0UnfKl7p2kuDbqdVor4T
sOvgI9T1/1bzn0NbOPFmw7q5xkcrhpXahLdXRp8t5VWg03ohZfFKyKmakit7K+qUtAYqJSJlYQvB
fQqcMGuzlmjT7YEJ0S/5rfzSTGJFJZRSTnB7GeJS0aOGY7JGa1eCF8C9mJD9TfCn/fcMDG+af5/Y
eWa+0W1pi/3NtrFehNY8sgh5W2knAceybZowJ24zqGpCNVYzSDB0KilCSYvyZ2uFGllH96VCIDim
Y3ileDJ7I/C+bDpyk3lpK5cTzb7rckKHzhQ1bC14gVrKYl4NPpVyE3jOx2CLDiKC/qdj45bwDR1/
JiukfSY33LrVTK6J3KSNwvJOrQnqpT7l6gOuaRWn5HYbxQpIcB1vW7g/xLxcR4Ll/4Qyzt1Bs005
r137vJPRBf4D8gStfdiE53oYeFDSVErMrw/IvHnlJC06E9pPGvApr8hughoVUlme7crtKE2bRPtG
nejHIIqm/nnIeDL8UIOKIWJaaPEdtDc1Ax9XnUf0w3+OcJyrN/bRYK1Y+tVzp/EUybqE5eKscbSe
RizgBqQVz9mGP8+hFQSoSS0pEQxpPBoW3JIdQPmh98mokDaaQCdE92jxkn49JCR8ItyfdKJKHwX5
d+e6c1xVP0vPgyvQZYTMxi2UB/vsNr70BoLAn3Kq/9bur3eVtVqCYOuTaCrjefsykNmYvksdErM+
mWLrO9aeUAphIGK+ymqxfDpaHQwlOgwFuHAYQOuwtAl8Hx3zu1EnSCy4tEtcYjdFLJnJeK0XsZdS
F55xRSmu8W6O9jQqpN8rZXGuhfzQOyJQ1FXBYiSEtkJX5oZSYyj4o66EFMfiVRAdTW0f8WC0Ez9P
GN/N6AdSQELJX4jkA8u9thJF+ErGKiA3KzAPGlcJhlibdJ047yB2n6fWTAyUPwcLeJAJ/4YPPkfQ
qdgHZBnxY+ZH301oQbN5S6WKYFgEmAMtVX5XWhvPB7kLj8HC4JvyzQqCDrqp2KkzqTo4HJaud7xW
+aCHZ4ESZPjRy17U48fDgM2zlAS/s9z8115u/L9GNjK//mCZ2gUEHrYB4T7GHwLprrBEDDRxwfrX
eBC8TlZNkPFUQ/pMUvYgkaT8GMee2DZKR/Wv2aJ9a+oCp/FyuOd74B5uFsOVz2fhGf4fScCdQ1fB
suUbbmCxGRw0zgv01k2aq1zERLtzlllC4TY6OdUIi02h7M6ZEGlPVhedJokrzcPmbijIIY0gjYD0
tmmNBrVpOjgmNmUF/g+Ycz1OYDC+yVTWhrBo8+Hu9JIEADiLMRovYEK5IKrEtCoFKn6tBHC+Xw65
WgusgHTbp24jDMBystaWqiCokH0cvAADArlJKzE/DgrnQVEYiWogaWa+FErq+wIe/R01dQTJyAmR
yeiaCwOF6M3uZksq6GisJes5s93si2o3kuK8nprIHKqI/RyF5jLbbUrvccay7CXJy9znFy0BhZqU
dullzahCnnhT8rvCCfqazR8FwK07ncvwmvXRZSmQkU+8W8TTsvyo9toBeQ/A5NLiFqETTYvX/8be
9VDCKCqSwYhG1XCNpai5NWIdPgGHEZS5iu0XiYvKrkJAZHUJ/BLlCgbokxhYXsKEjkAenKs5devq
jL47SOKv2vxZKxAtXNC0p4oQ4KV1hustPXktUSi0ERsVuhhedzBTbRVtvfeRAXAqEfDdFJbphfmr
lBuU1rfEb8jTWYQAOxu9wkVooA24WpvkdNLL2LpR9GkJqlEDEJn0rSvcHRu6CuYzF/cd+26EUYHc
7kN9KfAECpbRaZtjIAN8SogV8tJ5iTkDzzKQAuqoG6wl0SjSap/hSd+w1X3ombOajP/hw0Tvy9oF
HklPJkXBq+YZGosYp9nIfxz5WDtDxIi9n1fwSQ+AQtqkSTeor3afY9xgoivfrxBqsZlMl0oIX9gw
QUKd/CXwrA2UxJKfoDiF4B3fbW3aekzS/q99yniCax7mpDM+60loqGvyqFEJvxqHQ3IIQK7C/Fty
T4iYqRcZRPJriKcbCwH3jhW+A9KodbDg+HU1oivDrki/XRNj9mC1BLtSNDUWVvwFNBeXUC0TN5cN
/Tafq7lPzhRwnXgVo/hn7F2zLgctlWYez2tkMyLHtSCHixmVKCaW89301Vb6O9A5ln5WhyS70ADc
uJrDvtj2l36lWG3XuUSznDiJHu8p1TWFVGKrFapnuDF4U8y1VVfqG41b0WCOa/55ZFjpKRTKTsEM
XOZkHpdUN9Gwo7SOwoEAsTAA+BGWF91YImSL2ZLG8slhF9Ps29zujI7see4l7lf56wE0LPFcZJ5o
lystFOfdkxEJhVJnooQhYKYBiDgMG4JxOVol+oxBx29t1wA07UaEgzraiOSISuq0108Y0YC8bLh8
GnqU4XoHF6wsk+mdltbQtOc9eXJo9pHbBCuGTrODjGFWmWODB0wbYM7uWoNOt1rUR8li0oKre8pP
ZmNciz4gXXsAqkV8iUv4on6JP/uY1Su9tzk6ZUT0m2VSBc6xmvky9JGlUbqi/BI6I6Bq6qXM+4Ib
5JHBs8bPy4nNv5/8rT0BVvCDKs29PJRpNEnh619bPJEo2ADg0gSkD1fWQxWn44xDh3tN/hDeoeUj
MhgHkAkjb58idmY3JFj+IOT6Zz5O2A/w1m0YnsrMOhLo1CBBNn0oWPz4auBs4oIU5H4FS+tcqCr0
9ldUMuSW2M54TONm0jMluiB5qBQK/V+4dguxdTF/MCIwLE8AwM0YhuoHghAy9yRalXefwJYNCnCp
XE5YuRYHi969IDla+61BYC7l3lv5e104IVz1vULDxCZ6vmpsA5UenkiTMxO4cCqzV2m8sH3tYy2F
X1/gR5+zI8I1PstqnNU+6L6Cy+6EhxX9svOCUm14HrYalBqd6L7Qh3+yEzqUk7reHdd2QQ5p3FjH
RyQCaZISBEpq3cGEUhbsM/C/JTQlF1wbmNqbUR81AopqzayBglL4dOGGg7y/xgzx2V4zWaZCTrwo
WNRA/+H87kuAGGd6gh0gP2kCFcLPTAzSTiYZ/j8hbPLWiTWYfjVqWopu/FCHdDxc0C7IcB9ULHGP
zdFqQCJe9yNBfFVsxfVBRJn8vZ5Gy2wd8jESUeHQizCSphj24y8tBqUoPVTFhWIYAvXkqVVJkaEy
3xfn8IV43Ti8Uojn0Jppi2x7UG8GrEb14aQBrpKFRO4ldNJebYpb3Xvbo41qyuwTJ+rXbICazbch
gk1i9MwYNHufgVC+b0ld7onIbYH5uLYm1eiJ2GGLsKhBz0TbxQf5K7UfR3DdszYy2PwI9H0sTLRV
yjthOxkWIS+7jehNYsxc7xe3g6IsQL2SAuzLL7kob/xOKpqdHl7FYx9c1rfZp/a1WGAOzfvWZJ0v
1MjdBs7qHrVwe3O5z0qR9czAbwjd9DgzGv6FSXMag3oSVv0fTYiwNzbQZi9dYzKxfD6ZXrFJ5oaC
zlw5DvayOoWPxGjU028BACCVsliaKngAgyAA8pRdL2C1jkp+JQbcYSQi6Staw9GB9IaDoN0PSGuU
7+C/h0pxYq8RMDVN5+xbXdj1Ok/ctR6dxXPH89CttekLttnH3DOZhLQLv8KvSykkrP1snNUCxqFq
E2nunHNzPbCG5LoVUBj/7W2VKoiJTDYR2qSaxLmuMw7vCGZZZhljk8vf9HVGN1+SeBPz5gWsZCvg
zrxFJQOjw1HgVtXK9JgHNvFrdOqHwktLXnMNV5EZnOmqvDyoIjAWo/Tsr9o3gs+xsTi3+Lh0h7Z4
ZX5llTbE9QcPHQzd5gyBxfqTAQIB07hAhzvjR1kRGlgkMq3cdH4i9Rnmq2j3S6iOBGwxpRLk5Keu
cyDWWlhexCkjgYbi6dHlD28ZrJkCPQzkh1Sw1zi9ewwGi4aEC29+97Gesg792RYIvERRGn+IJZtp
YoKBrAMLgYAm/RqY7UGYwudF0Tzx2CvQwI7gVPdXsaI2YekFIDc8tuWgkoRzuHoaWE3b3Hk/jxk5
YFecb5r62TO/h1i3Mqooy+JH9Ed4JZI+G4UpHpM164iVkNyt6qtuDVJy7Ym2zygtLL69T6xdv7HE
eXSEM3cDDoclYMiBUVAWi4SrfVZDnYaK5dp9IdH4MStL5yzQezy4qMjT/SNkfXyPIzfsBEMcQy3z
FExFYWx5FqPbAeS1VMYdLiwceNhX1KkIRNQCoJK9ikmtq+8wcZqSP6LdZJf1elWfdnS/xlBjUbZn
wREBV4J5Qi+TbdHbZrQaVmtfiwCKqOSw1BwhGfiD3W0XgLZSVbfUON19ljzcLlQ03CXaZuwqUgJI
imkhj52ymahd+5wmIxnYgzt0o0UxmNjeddfctNRBMeGfIn7Z+NnGTcHOwbarZtrfF/sy/v/SsNJG
aAOYo5jonXApQNGZAL3afEuy/PKKmounR9kh8cZuKuQQ3r4UGgkjE8LS8FyF3MI1D9yDwMIBMrs4
m8AXyAaiMk3auCOtv66hacPdclRXh5NWfgEPG743AMwvElH6KLbwfQn1V4H5O0/O+waTNaaYucnE
sKcfbiwpDVK0NNg6ul0JAQUg+uogFpYL1YeZqFvJz3GDv7DBWKmN8fYaYbyaWv03acJ+SjOkUAUD
kLhxDh9g0YLyCK5Yp575RgiqVAjymeEepXfImxlm+wJm6JRHgxGEC98N10AQV7l6lnUye6trTn8G
fWoPNBvgBWyTbjuNb2aTB/aFXFL/GKgoELy/+TEyT+ystjOhueiaPySJk5ImdhdfM6jEzxxxPK/H
6qDLHSwu9wd/AQLUDJ740GOsu7Q0/IhTu4Ylqa5WNa0bOpbx3tH43jxvi/OTxNh2aq4yyCcwlGYY
bRrBGhk3VYmgAz6/mMu9OAnGq2ONa1M2FirifRlNwAWgOWTdeyvH98Vx9E174Xb5h9AAubPRaQOn
XUnnQ3LNrgE3bvrObyPAbWCK8UCVvj1Th4OtbA7/eavlzd3f6aFGgmoVW1NWfb777/I3biwTHtpD
6nxLLiGHB0MChX2Rm6/DpFlGZzc78apZkEKaWCqA45BJAbz1gZvP58fiv+YyIUi1p8KkTKj4iSgh
LOafNRDzqPnueGZW3mzygkB3J/PvQSttmva4lTwAcvxQmj2NC559mNAgxAObbH5nc18VnXVAcEIQ
5OXHNfEYTP8J4Z8QSR767N7CwyMYbPFrtUTT5kx2Lntox7AbRnsQqnNVq7RBahB0A6LKRyX38L//
4HrOTYaaCoJRXxBmI8x9RFFIdV/PBtG+lg+u7UG1M3EN/tn19wSP8e71obmUcCE8Ubj5n4E0+ces
sOnwt4EJqk0qbg4KgwwpaDLly+HXEWcBQ9QxIqrqD/l63sjtiSCvExsoc9ZP5vlImOIOytYxoUF8
7tSjewjdq9+vDu09F7WD4UavWhMNXSuZKSliGGeJPZy256tZEJFb5NsXm+f4jxqlEY7JMBSzMaTj
BQ93iOoS6N/yVswuD6Fs3Mhjql9ExpAUSivqndcdOW3WyKyENn0kf+OizfrBgOslMci7/4qsOVdK
j6VLqd0na3+tsiRzI4EV2H8DHnttl+Zx/gNsxEnKOpjTVP9DdFkNjpvIr3MuavD38bpiFfERtF6T
obNuoKkxhSyPAerJo0I1xIC0z8Zxe1OXMwf7LrTtfnm2XGP1eDsLF+quOLMh8aUxlZgCtztL83dM
Bn6s3estKGCUfiw6FNOqH5lDoWLMd4oM3ZfXg5SY+KwzM6rQbGvgygoFWHPKiIvlA60et3ze1RPw
Apbuj6qpoDo7omeLjPvOo0atXCoNPZjzzxDo3S0HwKIMY1V006Uq0Ribga3joIGh5CrpQuNgqlQ0
5yLFYTGZfRx/ZNbIvc/muUQXGAc47O0Cmlot78fWR3L0OIdcAXbXd4zcqlC9kJH4jfq3GRAUBJgt
p0b+UH7NLXyLgx2iPHi3qld7rxsaYM/Er+9C4crIeW4RURxqIVX+PF5pAlZTsitEc01H3USwWneR
96oV6EoQt5jIkjQYa0IxUEoReowDf2MWMialcldMMM/cbb12Bg4wSF+lvJXhzdUfQE9BV+Z5XSmf
sjhZMfxvN/SBk+txvES2MOHh0VXDNVKx9tAkM23mIjhKHgbn2FodkAoLg/JZKmM0Lq6wi90FYkfq
hqMOzeEZIiWVrJEbS4WFiaZ3d5FZQtVRTDKh5oohv2np6qQViA2Q3w5jxioLZkktDylcy0lKDWm/
+tqJpU04QMALHUg3W+pD4fIQ58MoH78aCbLwS65KLejByZ5OxKtP6e0KJnDLriEBX3JBMpwH49Si
eox0CNYcg/tpjq4//Zq7GrYVsT8Ihun2KwE6VksXp5HFihz3pQBZd+iIGJucRYReLmQPnl1R/dpX
Ktp8eLn7fmBinFdBJe6Bt12zK6c3lvhNOTjgv/g+Sm1neiBNTs1L9/U8evQ8bFQ8eq/wUtu4OikD
KtgUhIigeQpPA2qwxlw0q2bM/JWxvlUUpUpIAJaGVLCE+8cifsqCPBCofatL0GjxCcLD8l1nubmk
QACqA8nJh63EUXk3Yl/Cdyx+Mnndq50JXi7y0HMvdhiLO0GFvhnjaBxDMx2MGEoPLVzj6a8xb1uz
N0LzTuZK0V4zySqS+Ns2iSTbStH8gqvHitW5W45sLCr5E0JMQTc+sUxCn5VdExN2SmkVPyVQHkKr
pPAWE/tCZ4YNEh8U18HlZf9Ztc3dKqK95CQWK3gBgW0AmlvZo3de9dflC0TKW0CT0IZrUV9xBh+Y
20Gtmxek+kRX+hWtrNOGdtzcdHouSD3Qms87Co+fi9T+LAUhX6AsInWbd9kIyikto9meqeOB20j9
TmhZX+CyeoP5xnComfPj/rYZkhlet39ac0/PClehLPhfiZ77pNf+Zi0cqEM0dz+u0hec/ZGME8c3
qBxvhVZY/rALn8BqYIZT+02a2EstGmKofTAm3Mb4jIGB7UnKk4PSYnaTP9ppaJCk9/TliQSx5Sez
+0YBFx/Fm/aIT9PubXOsb/VB4bCHJs9ansWlqEHY8Ncmn/RME0TyPVT5EmqajciN4AUBDMDPmPVI
jWZ5ZCB2cbGlrDKfKwgPM58y1X2AkZ0tHB1Ok8tHwPD+IRJxKPtFx9+A5oD+QSMDiDXyXq8XLHDN
aUguh3dI7orYkDL1RUzSTX2Umd4kAbZ7WPqyqaXos4bPIs4tiSHArlLmgavcFbmdsSu1RuAhRHPz
QITV9GbY+trh0YTErdMIs53cRqRHnbu06BK/fVkjkaxfEaYD6fsl6m0LRJDjudAMZO4QRqPJFEO4
ALsWAHhhnOjUIfVAN68X2qc5whSmFpPljv0z1D2aERDCpbNZYwBwVmM4DOYfP32TqhtE6YE19gAI
qnUpFo1azLIkPqo23nYgN+np+aHH1ytMKhL3KXH924J65AX7ejF7+nX1JMRFspSsKxG33ar/I2wf
yDTWk3S7nDNOFMkk8YX+pnW/hRtSMWJ8gIPC13nNsxuFzre+baC4qB2VHwjhil9CQmvV7ItT09a2
iiz19eTBN37XalmktAQPUstk+xtMGYy0T+zbAZ2TN4llzWKZFoln0QCbreQnPRgMQ6x47sllO7Zd
rJYRVD+QzFIgQc2hh8dhqfTyoj8BeHKeqn6Bt9AZtmnx5gQnPmCnBAj0pp85MfMCBikEb2E++vu2
KhV1VGdXFRCVtVHgiL8/CwJ+qibhe6+JLxJRR752fWrbbaNY8l0X81603ojO2agH7Me75L4QlJIF
nTMk7P/rTfk1ZuHRzRZvS/O99INYPluIHjGOUT3ZTbj77b1maqBoWr5oOUgbMY7n36YwaxZ4+ktZ
IzDkvFM06BAY55w/ZFtJblgh4w3h3Dn3wq2v7HWSLkPS3dOPFL4jVNPtqSnsIdWXQONuQHb/5/L9
lRzfeYUfbXsVxPDE11hKxuXtGoLC9hzdJa1JQsA4XYMBr29tt/KDs0KDHdxBnA0DVxl+EHK+qNkl
16XY9KijRshK2BMHlYxEEv+BZr3ur6GrzgPi6kASVazNR4GCgaz3Li8S5iDPmcAlZDn4TlEiLHBs
2EvGBMk3abZBGzWggx7RUqTcmuOMLVsjwL3B1BXJqcfVZQWHVlgTnXs3ZHkYo3TzUWWPppKjCyZK
0PyJQu58Xa7mUtY/5z6ZWsPPZ/dUa8RGm9ORwvNBat6bwp4iG0ts1PgvJJHGmtcx1aWgYflt/U1b
wSL828a2XTriCCsiw0C1nWwbBlOFM2wv49H/mZRZ6MTR76Ec70d9BO2EnX20HSfJSkxx7nOMc4nv
jy/H5xIGt2kYqa2nMsheRf+8zg+C5AcxwhFgcl5KqdgG1KEXZwF2oR1RzOYPzXGcBNMvZMl5XwvZ
yBrEhZg4Vl2jzQfYOLw8vVAKlkijs5xcW3Y6Oq0Eii1Xu37yVn+T6FKzvxpFmyG1M/HfpliPfXw3
XVXs1tWOiaNCga9r7LDuYDL9o9zFAZd53zU1/t1HbHVzLcVk/tpIKdCfwXMeqtpiJckdb9JxELRU
TbiAnOGxao8qw77RaCFrBoQUX0UqjSuycKOPbTv48GAhSvWKnV9frwxCeiLa9FHDxEIWoQkcB6S8
eN8UN9HZmIoRJX2QU3E1lKg+frbfiedbOUNO7Jzf0G1UKUqg+GmREqbcsk/1S+qr3MaDIDPkJgg7
nVcSJ1uDHjGF7jNtBy4hvBqoAuSY11nBimPx9SjWFPONOtFAl3S3ro4gRUuQoX97EWT/7X7SJ5II
s0AYmP8WHbOlu1c1JedszfBd6axd3uKGUYWYqIIGxilU65KPVG/8JyHVLNw8ZQ7Dutfll27Qw6pD
YNROrPB7EyDYldrJgMtmPZszo2TLnLdGGYRBZcHuu+aqD9wAFaeIvFWgT4ITXjS1W6iDJUOs/NCz
Fp+PsUu6BfJp1/yyyieAznuSJ5h1xhmPU9PVNFiphkgrE1efq6a/wbFSscI0xT6TwXDrRwO3k9u4
ZQd5dtJSoM90wPQ2WIsAVNHwCIqB3EYXgom3xUCRASovD3jlLYMkyBu39v0iT3Tjx48OIZSFw39q
llEpucnhFv+5ZtxuaJqHg17etuT2yU+dvO3+/YuGYj2TpaWpMXZLewUYZfSsN6BxFHtustDulKmB
gXpOk4AYMdz6StnpYMWvS/SZ6Xjr5Yd+5dtngtb4txpS2TbsEorq8PPKo5dZI0uZ6bQ2yeyB15pz
w3W/yrNI15DkzVlIuJXDLocS5CRzrCMLB6mmUjqPLVj8o7k6XFOK81ONcm9x/G6U9qOc5WYpILQz
hdb/2WfrMhtvqFiHSF3zh84g8fatV8StG/Jhq6vHRqnMOzceGymPV702ikhxoewB3AmJwHc2UeWu
+X9fARIv5rdbDLZfgxNqxgUq3ogawiDxKKUGz0wapBkjdE1H9lhGVCaXvnqewy5EGn9k0UIhbZ0r
MAIFJ19YJiwB/GMYDydFyFcEQrTN1jNtrRS0XfTENOPjEcskO0wWJ47GfsYUi21tvwuGXtEm7kH6
WFiqTbnsuuO5412Y5Yh2uzVg3QEmMivgQcbhQys/Ni8X0l9WiSvTF2LfWrnguuKysQYemoyd7jGZ
QwOUnRrWKcEogaRg5UQQM9YyfaBA2iJql7UDRRfeaGgj1ch3VN85P8liPywmRRs3oesEuX2YVCzl
Fz6rO85lw6a0pHAqPQCfpdcRtgaClH8vSfrO4VTFn4m4uCiHuyYUbsrxrpTVlQ8BsrH7WTRWpbtL
9JYxsnq7sCZZycsMuFdUilot3bxWGDgMuAKrvws00JrlThJoORQmV6KcVp4YRBeSqZUAhN7oRjU4
wnxpacV0hVCCTNUcYvkgMRNHi9rLcVau6D7QD0FmRC/cBsE525VRawz9CBzBX7gXxhasWr7qVC8b
cqxuN/PZXa0fUSsPIPN2ke7WM0t77CPv3L93v4KW8+DsnKmzpCjnXNkppJlZ4XwWrOY/3YrZyfBn
O37PxeRL+Kb2TUxqCOihOewjAJzKdmrAPV6dho6j0tS00p3c4p3Ef4tj37FfbjzgV5dIy3wC/kMA
GPUyB97egYMKTt3VoTd+gKnEwGWIfoW08+yzXYpVzclYF9yji0LZcJKYoGtL7a6tCqMFinX3RcEk
qrWRGdFtqzGEMet1w+KB69JriWKdEAwrqgnA0XSoLErjASxjS/+HJLaAitK4RYkiSw7G1DAHt489
ZyRGnCom6E3Pev+wY7qaVUXmr1bRrK9MHVBDBK+QSNRqag9pcOponKb6W9M4H+/CovXeWjweuihF
9erQia4jWTW0Qbm6uSAk0wL3W8Mrgj6fs7PHCWuZ/0NiTOgs9RG+QA3B7JtqoMwgIoZljIDzUTOR
ZLLvg67sPJvPNddroodLJA7ejF/8oN/2b6xDaebbxwavM6aY77l1F/RxS17hbmJY3sXDyP4W9SHL
Y5o5TsSSJqNKvJGUHuksOJY6HudGArL6Okdi6uSYH5q31T0rhVNv9EpO2W01Us2St06ys69NeI5l
wrJ6qGPK/1ZKZ0otRR02UvBGrg9y/1c5uCZ5pHCNv0Hno5l8rRMcvT4f9wd0DKWrbG6AGTtFHkEH
AJrGM8vsy9nCBPYSA0NyPxEbuIbFh9Ygwye7V74XVScguTTy22Pnw7KIQmE17oZ98ElpB6vGMkjJ
yYjYJCNgYxr1LETlMWF163tXmLFf0jTe5r3e+RXbkpo2Y+uGfGWztwdxqwyIF0GHToYu2deS0gEA
b96GmUnHVAYV9KbPI3mT9ZoO04ABCjcZdxCLoFSnQYRPs7wHYnS6y1HtSNsXRK+cQhvbGxnPxJW1
nQZOtCY0oO9btpTPfCC116bh3dJ1Qj2sKDevAcstXzv90j0MzRvPC8vzcB1bbZycNwd9AuISqMrP
Q89hRZeB3FxiXbt0tuinUQx98SdAfsy5s2FcIwPbEjERzaoBtow8EqtMElxnBnt/1770f+PLmUf0
rCOHSsel4JLrlCPLVuk//Lm/GxUUf80pyWAXOSX6ZMKpwsEX//WmC1B2XFtghfMom4YBdmobSpPT
grr0xqWiLz84rgH26mKr95T20CKp0hBCVO01Iqh0uc3tUXU4tb86ChY4rISvfqVmgBmjnRSXo9ax
0Cx6Ho7CvzzXnj9W6iApntRNPzcDXgRGeYHL77b/r+vyzCY2HmVTeFwjE53tDJC29MquGhSqoXjV
zZEjRqeXR75cfI+xbhnztLPTQ2zAjwsT29A35aOU33Rb8s+6lCKl1Gl4XQFcS2fBQMm1zlCLBP1o
gpovZ11UA3EYtvUcFLQGEQJqI6dEuODV/1zGMhGarmeAKHak2Fk+lLTSytPnbP2fhii3dFKuW21F
lrmPH4mb/i+izB95+ks4poSPsQNYFkMk5uv1/wuFOnR1CSVl6vetx+7KD3YdI8x767a8j3k2jFIL
woERs4mZEsx3LXXsPJlfWJS7dQ/y9pgB3er/rpZHZCyILRv9gFR3DpYHzhQWxA/w3tSmI50DBPHJ
CIwOQSOeB2WWEkhDtw0TfqGwg5Cj5cQ1ShXSnY0SvfmL3F33NTlaHh++DczvIg/QHCa+MLD/2voJ
Li8WvThJoORzCXTzqGeFBg10x8zF19O7/2Oc7O2RRncM/Hdbacagc7day8xAE/a/HGeSsaxemLuA
KVCelkAxJ2pvdMc0PsD85EXgHxJy4X0V3KQhQnTJ+/AT+08zIhnvo770MnT75p1ghSUcYQIBcvCv
5fHIAjvlpNngHHmeVldIb1gq1lLv9QyOVFMW7a3t6ZWRKB93ALktUWjth1hWWaBxS68YzoggRq8N
G4KoaHTQhb/5XKijAykdYcbGU7M43HSiVZD+iUMV+O3+pf8FGO8IlsFH/Oc315yZk3MpOcTQGIs6
6FakBf1ShxihUASJRlrSjVSExcBsfMJ3QBoQv37IUfG6GRGdpWPSX4nw+WDwURbkaa5vwHP8NaWp
7p9vJdY5W620vfHquiSBU5K/WS/yGmozR/bGTWQRbhs5i0/9IMP6Ba5nP2RRz6Lx6lmzpElYyHZd
RUheQKz6N/aPEnep0t+/vIzDtUHt5AcWH1rQmbtvrZLFLrBN9l5N90x4h15umgrUx9CmvTy9lDib
fie0Ku7oUkLUiC+r4dG5A6s440KjoRBzp09PMcdIJ89a85iJzJThhLaxG9z41T8WadXCWt5djyzm
Pq4La/Z0GkqDzGbFgEcDXpUrXSO52hKpflZAAQBoyM6XAX0w0DuxvwiXs6DX7KY/CzfdQRL5tKeP
8TpMBpDZPClEgg3mYVdCe/2Brwf3dhlV0cj+ab3ujF0PC0lWULbSRLZO7qo2J87obhUmzayixYb9
cGHsejQ86fnzqZdovfo+NlEaC+HLPrJcrcUpqRTQNltpytQBhADKtamkOKtPBnkBNmywnMkALblx
Yn53VUNbNftxULTAUml0RLRw7U9Fi0AmSIJO8ZjY9nrHsue7ThL68smbQDRAfdQ+mmNCE2YEXRZJ
EkrzRGjuBs7QNa+Y2t8/D1SPfsP9OGSJgqyhGTbv5K24QZK437Bs7VwdTDy5/DJkUWR8MNXmxKL6
ER7wkgjQvnYiZYEu7Z+11HkElDTxGcredahJaUZ01uCYuG+IkEjA3yu3qwH2Qs8JXscnxJYAN8zs
lZn2H/i6KXyYtlsAoC/ErAYdRZTSQREUg2XPHnYV2XGukalG6vcUJlQJ7niuunOPd1RwBnug1Pcw
jp3H+FE6JIs0aZSEaJ4bfgjjGfaLd+7TPPGh3io/bADN6WltrPRf65kOhNVW92VIl32UVV9WREUG
e/BKETjWJNnYW7Gw2aryhtqE5QGabe1zoON8fb9vkQRJuXhy2hHo+gk+Z59/PP+Ga3C9zedd70w6
Skwbq4DWIfWRU/iiA5GIs/gaVyFFJxvb9sv7aibl9v4C8nNqfLa1nk6YjPDR/4F1ixV9MlnY0zG7
YH9I+a3f7SibnTt/nPvcwCLiHzrh1lnPHS1DvQigz4jVvj0lBE63SQkwfFCvs+THDkqRwrL0QhZ0
SCi7ZXRS3A8L74/+OtZMWvNkE1ponKmEfAQwod78MuWABixfKhi0x9nw6mRT4Shs961LQ19hw/vA
p+xP26KB0VFVdaHlxbj0x9jD4SyvYRYV6k30tGE3Xm/hFNHsL3+huheric8ozarzoHa5EN1lQNxF
iK+4RUwClkVgTkOnxdiiPaF/YWGArNGs2fZHWKqZLnH7DIUhDVVhqFiWudGnhlU1vApYBSc9SDcD
02dHrZzZ2LsmZ2aqo3XWO0lLegqaa1UK1FH+C6/XR0pqqwSoYBcSK7om1rHm5rRgNQOz9shKoh+R
4RaRrgGROIcFu8/6KsvOUjW6Z+YygMt5KQOWtY8ZFgH92PRHZT/ONXmi/4+3xZgiRPdhRxuCStp8
nRv2/cBorSQwOMR9yxx577DxKHXVY8JYyw9ECCoZ8/wc25CtC21ltPpn/366gu+Q8Tkg5QYNQQQe
FL7SLhKyE7Xn5GPoUjNU2iRhZZ2sHV1NrO2orEEvkkLBChQTD9hVC5yJ3fa89a520dNe0zMGZIi6
JYW48hMaaf7Wh4CThy7Mwn1fRHGcWPTxDv8+UfO/f/1mtQuJgbMGR/FkGGz+7qZocWddTMrWCn+S
HjnxYVa5cHBcpNJHJ5KZNpD0WNTNucxkYOizkbT1ib5ts4RXlFICjbNLq0y1gcyPHW2WkQ8B2xW/
BlcwJ0m4Q9V/REUrm2QvgC2V5qxkzoIFfFr+9TjfW5Jy1ZuRMrmhBo1eQB6W9Wu6XVkPjxbMqW5m
/BYh8E7V6xu9vTk/2+1slVgvZ98nxTzMQSlC7yJjSEd7BE7WeUK+tdY4j1T+XDTqEkvCyvHMRbgV
6g39LtiyhXjnjLZzS3+ALb4ra4RGda4ZzBQUNvCdfZZN4i9kpdHyEc6UizlHpgH9TO0wmfdLXATt
WxxqXosCde2aGpqvVTS/VubWJ+xcPzr+04934BG69Y2xskrJG0gCvrRin/g4CzQmwYEkFberPBJ9
5nfmSHQvk9yiaBB5mqwNX4klIw602M9ChlHypNGrc2a8Oz9oD4t0olLCb8Et/RpI2sp4poTUOIrS
VnN2Irfd0oSJTkav+OV3wbdYdTAfDNqEUJsw62G4cO4cWBCzWnaOel4vJgLRQ9LTVFbogZXE3156
5oRmvqebtPg8xM6PKS4BcZyurenjDK0z/qrAcAbdZjiaFOBiYzLDJbttRD6t++BK4+0d8AxnnKJ7
Tam6uszH6Kkh1Spnhqtgksi8wp28V7vDfH+IdgBVyxhe1S+7nWFxwzzzBkVQPNDWM9k1qrBmHn8h
kKSeHZkVH7TKKM2b5J/QgY8LTsP1FlQP+5721NT0slvr5pPnm3gf9DCWX4Q5bUpc86dNHKzkeB73
d1e1Ja+bojlEiuhRdORCjOCI5IsET1JH74Vx9zfzFXZUq1aGMgd7IBB2zbDHZ1wmlGoZSTqtiwz6
y9FsffQIqaNsfCyYRmXYXAq5P+WlfiMJEWtSfyoFNRu69l6tlaLDOnnWBhoBpS8rqz/fcS+32HV0
LHzQZGK4ObA2+09yOJk54HoAA7H1Jl2r4R4XrtvbP4FRVs7cE0DbesusJVifoAr75AicxxRum7jW
MoeMkUG+YLDoiAhzbj+WCyre/USdeGK7C6gf5eKYCwCG7qQrVXM5SxTZ5F3Coc7KyaNKTRd8T92Z
fJWHK1oWb3F3TYgToQwfelqm3HCjTg1E12TA6bElkSpnbVhwh5F4EeCG7/OYBWfV50SPp6WCxGIE
JRyjPsIIzU71f67n9aa1yZgh4dm/UGXE+wWaM5SxtBjI2v0Tt1hzLChrc4n5V5x88NKhCgsSHF/G
i9rFnaG3vsSskVazNIUqbeiPIWeim+IGP5SvmC841m6X8iH7v3XakrV+uA/jBbUIEyfVTK9NN1m7
UnNOfkRDG4z6aw19KJXU9gHqBOrxjwHzx1GscczRgHPuKGB3MVqV9AcgqXKhN7h5Bc6N+KCIC5yd
kt7dEyItrN8a+D9v6jOUHBWFs7EFJOTg/ee+n0b2ET2E2YLhr1Pnq+YqSeBRNiBuuIE0HwsHWvdS
oNDJOek4ZykptYqNHO+SlbgnFtnilIFbYEvwKCRZVo974Xx0hYuiGy9RZrvcBLUD2oq3seQ25GQw
h7CVrOjrNXwc6J6LKxKENgY4siNpPdJtYcWI9Lu6DMKU2zUwGnTDgUSbLhXP5NJGmep3MPCaIXQ3
D6wXgz2vZbM6OJ57vTZ/Rjxpo3Itpexi2yqjK4Mr3HhAguVHozeir3JnD8yEQOhlMYIVBpQuvBRR
bvEp9eYxYc9Y09nT/7yUCx/xqGjUsg8ZbtE6Sg9zKypct8+vW0Cg/snYkWX9fXV08vhjfDD3c3SV
NNGn3B2Pn6rHx7WR0XlkjV3l9M8KI//cwsN+to+9M31zpx7nIMn2X96UbyO+0n2oad/iD38yb8A+
0Orn2tNG2lKWRBTj29H8tZ83uGN8L/zB3g9VkDNJCUHgMnOaNb2qfhkU5Iqca2axJM7hn8KRaCSf
muST7j0Co43e3F5Ka9HyNcGKK/E6CzjElYUEtVBP43e9pRHaERy/ZNab8VZOwjMzfv8AN+GW3EeH
9DTNfODYBiky8KGYPU8cpoUJJ/ox/Npxp6M/NJCppStp1OT91rE5SIWyHSsq/XNdIJvZPC8PzRj0
HrP30ji1RFp8TtcRkciWiz0OyD0feoyjFXoWt2JdzU9Z0KmfzMe54+Qyf5EHsCg7VZ7rsMIVxSKk
D6Fvvs07fFK7YSCx59kfrX+yAPmL89jaky1KT56JyW6sMI9v+xKL2LANtvbScwb5LNhHgfTVQmjn
kUlcwgHi0A0do83oQBeJyTtc9ipsmmDHYdCp9yCah4i3NXPVhbsEV6mdE5IMWjK/cwIN0E/Z1Dkv
YKXBVlDMXZbjTHwSP8jCbW/DVOJpkv6aSVMbb15yLXxN8WlMRluccxI8Q0dL0HkgSh3QHY0mN/PV
Os88qjNhqGflLyGGNNnU6kYW68UmJ6JSi4Ch3Dm4nsg12P56ewOdxGjShc5IW4JzcuVV70psYTjg
AdJqkShrGfdagHeUYKL0G8/HH/kAk1khfSn7AyUsIElYSCuvrdDmAsUL1wLefoNDdt/esZx/Wmb5
Lr2ua09bz91Cx7m8RVCbclzZOa45vqkHJeAupomOZLrUS7tJ298ssBUUgqPg43rD+Jjp4negkGQM
4U2DiGbzYFYIztqrtUvSMLnlNV+0n2vLBgRj550y/W8gklqPGSV7jVRCq8SPXJ65oPtHqa4xxlk4
5oJD5bvja53K+i1o+1NCzuGg+AYRPyoKHc1ewiBhbi9VrCAV+EPP/SSrMgC57Qlw95UYKBHZ+HbE
ZZGoCww38IElDL9U5Bn+QD3AH+cC7BwXZXNuhk3jdy9NINp/m4jZm+q4DxD2rbInNamWrLDMoh3L
RNCZeoqkVm/uKCA1qsuC447Ma9j6i+N44suXo+kU1iSHiksmtsmLRwNJOiLYBB+qfG+6hew3WR1S
Hj6skPlY/gVQ0/u2x+eRfWpjBCIItgvbH9QGGnxNvzkg8ol1SlpWiougfixLRrOuk9X864hg8uCS
KtwRgNxg4SNm3SlQHRIeQL8Z6Ay+UbXsMiD06xld2V2rp2P1aCpDh9EbQ9lRRunpqYztQd0XrHmr
Oi2AQE0CvqhgebZwQYeQEn3OkmKHKCqRR+l2QgTPXi37lJWYI11nhj+VNIqANJ5VQQZoIrqzHLjY
Zn4XFRdeaFaOmMOjXMsvJHvv8ekscKnGdwHkEgyIPPluC+spBB9DO0pL6snZcnOl4uAwL6LSKLEj
VMCtc7wwW6vT8/as9liMf2Zxlm0E/drmFaS+RxaPLHjLfPvYnvjd9LssflicRCSuGd+OouEwJypV
WzmQxIADUjzcVcPZuNveiQeUsKw0ipdHZoxCHKEPZxhR0opDr+3xRhGHkyJRacvYdEOcjni2M53M
suApdqHs3CJXs24u7lW8edBiTK402rc8VtJGv2cFpGuWaFMLW3IyZOSPLUJmYzEMn6oRTyOPdDpY
eeGXaxA9BFgRCXN+FXgm3Y3Wro9Ci46FQapM2acYYcOPEy5s8ti3Koh3KMjuBglRsV330mv/jtzO
ni2lPqwKDP6a3hBhOQNFHox5UK1w9EJJyvPo+0GLu8abLsqNG6GMgWZxST+JD+Pvgn6Q9Na0T1qg
rXhRk9NJimz2j2UCvseM661HEfsO1lMUGupjXaEDqw3OsFlATOZl09GoGNajaQ2togpf+GJgwwQV
wPVaFeBrbTVsWc/jiMfXqmQuQs694VXE4XWFkpQ8AudSOZAIf0mleZtluGA4+gARX6EArWkHZ/dt
TRchpxM3ksVObWXeKJ3JozTChB2GTUMXfaiUJpPByI3hkHoGssdltO5oLXlLtN/zo1jzmMKLJbP8
nVCR++0Xr+pa8V4QCBdAmc2nNS3jaM7Dk0JJPUBR8ybXh4Naclylm5qy4qlerp2b3+bsrGGmRaM6
+kM6YrtVmk6NASEZUD6gc/rz/cuuON1ClkHEhYB4HiKJuytMnf8AeavSTd5rh15aJ9feFNG9eULL
lvj1BBQYBTGmRNBE9U/ul7ImRiH3Kj6o1g6aZOnAN6anAoUiI8RdNcD7Z/YKr+gL3xjxYkE+hnTR
I0h0EmJ4UsIIK/UDQ39cZWk0AJgfp2inV84kbCA2WqAB7WyZ9r+o3qB8EXxK49+Ci9IegIhnXPMw
h7L5gwrbdrWKQ7/R8OIrHsclQB62YSpugIDkh91l82N+xlzAieyL+8Wjy/wlf8wq3h+LDqTv4w2b
V7EuoCee0qK3nJtEkxxXDXwZBTNtJ+qSS4fJttukKApGAaPHSX3XIYZpzYUWFfE0QsBXGBkeHMr3
PHJ2zmSfdc9hJBJsWurMUqWQaFZH3dmdQiWCiMjV0vh7+QePgL65ZMo0MG6W3CFcI38LNCEHH0mu
pXwJaJnX9von+0QDW4dPpFSymLaoWw70U31bdbuHiAiuArfv+UgBnQ2aU8dAgI3dXu/+CVoVqAHd
/4ZFIx/0YqsiMFCx3iETr/oixtdVbcs/x2jpI3k68lcvrBYUsGg0OH122Knz/WkbZu6GjaUv8K+5
cVrJSo5/3zVSzFDg4LxGMp64G7sXwJu0TVJpGH8ByTNoQIeBABhzrUZJqRpsKJNNq8XCAFawO3gj
V6+zj70SI4vMgzqSVsfabQCq6vjPFzfBs6AEWVx+S3g8u9cta7SVZsJYuhr64ODLADYsrq935EOv
xNWq3zcQYyvceijB4RXQLOH4Jqb7EGvOHEpGVUbvTPHTM/TK2qrKQMlTt8ktLn4zVc/Nu7Nd1l+R
3ZMlFTe9dI6HzECIXw8XNzKddig/LQDt/upjldQTg68f8nS1mXuQEICg+LK9ZnWMXVh/qlw3/0vp
IROu2nquaNq4s615w+xqbjYRbWOQmyqc4oLIz06YQQlA7hWjNxkR6pLkOFtSUOiL0MbD8FmfVchk
ezyxzxzBTVNlI1gTEE9SrDRJMGqmP6GE3GRKg7BiiX5YRM2tXu4wXbQ+aC0Yn5BJNZeATeE0wkhz
5QSMqz1Jagcvbo/Bgy3ThSi4ylViLewdPQT1isuZ/7FKckphyeYQT6BHnMrG6wFjZTwk0x+fq2sf
8B7eotxjd5Opu5fLE0/KbpW1yDeLeNu16BODehYpMtgJV/aiRz9t11G82q+Yfga1tFg1grWW2nMj
XvzIscI4n/7FCcjPh0Szc1N5uO8SVFR+10NBSIl46xsWtuRbiA+VYa/k6IkFvVfwAeW9Ud4Mu3nd
2EhYemMyESQwO2lqyQOy1v5ZLwgryxvrnI4ywf7+ysrU3LUzYuatIss3qLrfR96AHyqeGDAknZ0G
GLzNhMdCkYFwW80HekkiWdPY8CoRFjw8sBHIuu/7nW0eU7swq5dsDPi4iVSYqgAkiRnCe3bQ2hCA
djRzGSD3HiHN1BrDYOFpQI00WR9VbhFxKod2RfUMNkNb2aokQoFJR72D8Uk9x4D80aCP53ihBAw1
5ojaUFPlsbqFFGXmDIzRpONAIaste2CkruT/lhecf1pbWXGbO9JwaAZZCfIM4lU04eysfdkCzhty
V0UqfsFUh+OQTdP+tiTbAR+nbSYRL5C2B9vDdVOi4ag25wXxdxLbaITHcdeRXps13tupzdVvEg4E
YzsYU0dMS9NtQDg9Y3RS0wPvG6NxKNYqkeH5yoaOZAAhE4YXYdNjqQU8/JzMECwskp6iAnLYC+cg
ASlbVIA1lkxpFHHit4AKK7a7qCnkd4VtjENNjao1+FC9FmANd7eN/4p4r3SXrFGr0zH7lIitLjTB
bdXesQ5p2LToIKUTN3NnjHti9CgymieJwztps7uOizBsYXerb0Qd1t28U8C38CQpS439kEDQyGjw
aSbvNqY58DdTdd98IxkFUWiwMhYxW7u4pPDgIdxmb8HacOIN773R95yKThkQn9UlJim797mRmNrN
M/2CxW8yXKAEsGTRH/fAvsXBofOwJqnG0RJwApzCoPA+cxwFBpjkz1LpPAUIAzr/2jFXhNCrGG6B
bCc2iWHzdUvcB2B2BiXFb8GIfpdYzV8ZKlxDd6V16VQNMt2NwXG/VAnDsFmSpvBP5u6IrQBOp7E8
TQ51nld3gdUTitw3/FfyrtatPtX9QTU7ElFdn48RJe0ua4eNr94fPSu4KFp0Dlpxg+efg73euyMb
9orwgjGfQv7lWzBO+SjAg6UIMtQusGJiO1VXTB1g8QT4pE18p99oCe3geWQlOVBatXUE3s2TFEjH
5t980uxgVMxCM9jstHGDDzZPCnxT/yaaosrDsuMxfj9JXI2rMcqIGKKsoMXMkg/Um9dIm0W8eddE
9B8JzlkLm5xEO+xAJKgCbJ0hKirnIIlK6+DhIqo0TJ2gEF0tDT3eB7bgBNRQ/6OHERWFnS6tk26R
vPsHJzFeSRJYRE91dDktYGIKqT/acShHFEr/gyMAXa3aMUdWwksLhgkyx+DMBN4nMf3+2w5Ws474
mNP9TgiNcTRo8zKaR7ocQ/JW21KTE+GFh7jK4PJ182mZLvuAywDanlspzwpKvjxpCUybucYXj51d
ox4TKOP22LH5ohhTVNnq72PuHP4bWSZX7JZTNvAbbeBlHR2ik1scOZ9bjbg6XEFEx+mXp1YGgNe9
rvdZyf40CxYOZUe7wWTZZOT5trEHiM9m5iSdlLErGymYww6C7e+xj8U7d8wd4hBsu+lOREkTVcZw
JiVczYCiGOPT8QWAzQ37F/I/lv/zNynMGVlhPkLPSaaAVaQvHI9cYPeCoW+/m+fKScnSiBH10Tow
XYbVm2s/MP1wPN1jl1ReENc692oyrkIE1dJRTneLh/0c3dkJdlu7kvK5k9EdVI4eJAPB3v6R9knB
IF/PU+Ju8wVJBhH1Q5jdApDi1C7Eh0pktL2z5z2pERuRIYjlK1Mgd2/xFVtYVJQK3GXP+O7s5aAB
xuaYIKvORShmEj19t8wE87bwpOnq2tqBnNGzZG5CXDamnwKbkTLk2kOTiFv8uZEA9X5+HlrRvtdP
F+n2gwW3oFvsO8HH7Ku2cj0lEEsRbWPLcX1aRflDg5WGhvPKeIjOf/cKbLe0GR6uCVxm3U1AQICx
gskYo/kRqw7Vk1jixbONX0kX59IIh9Q6WQd4OltdsoNLn2G60th70B9wf/hyCTXwkEMJULAtxXNy
8Pqa020hrZwQB7Dxj5woh/oB6QFLP7i5+PAa6qz/Bl/lytQbxX8wf/PHQHbKiyjdQHu4semdUWh5
8gQlK4HpgPuKVaujc1LnBBPKnUA0pyZiBbpWoq9+gmt/fGgSt2csuFSbiUmcf7X4YWKonZoMO3xU
iIQF5SDLJamC2BdrZ20Z1C5IGtELaxysLG4Tk0VePXAduzaGQaXXAylexzplZr7panLhd31hsKPo
dUet5bT7L2RDEGGekk88+LF1GOAb7b2Q+5k6TtSWTcC3bmYb67y2WfLMhtZHgeQRmjGLO8FDgHHA
JBclsk6jZhUGM10+KgOL1zXTu6gbUiVjxoaPGDOMLGWZNYTGKT5SfOM0Wm+y2wsgxpoAZSskmVyp
kcS7QABnCg90lYAr5fANy+0JOru6+6S+MVtEqPcaZcpSUAf0Tt0XvAbpp1wir7GfNQZbVvUD8u+h
R5nrPQiPt5Q1h0gp/aW8goEJ5489U5zPYH1gUfWy1POzTxTuG6FJpvq+OXvCuVQjEaMbA/Zv1YKY
jSKz/v2KeOGxd9mBHw5KTNDnFi3/MIUYgl14d2JeBaSp/BlWd2bKFV4EOuQu3g9nNQvAViKzyZp2
CQbaKWTG7CNYblOZYwnXVQOOBp14OL/cvvyvEcIrLIZJT/hyvIv25OG0t9E0sqtQdASmn5H/d7u4
dtm4awxj7sjHuy+TkkWNS0lnFbRkUFRcZZ9vVwJdgdpA2cKL18F0KdySzz9pebtQHAbT6nsjEn9y
vHUi3tPIUOGRh/vqxDmO4M1cdemVRoIH1Idf3CcVt7PNNc8KsvEA9h+Es5LzVs6JbkOv8YESeqaE
fanbO82BlfkpKjfUQ7OojSNg4Mdyba17whIbvzLyq8/Bvv941q+McZf9FlLiKb0b2QifFGHSe48w
Z0BjEoqfI4R4XhBRqACnW+wQR7zPzVJ5z7Uln7qWCy7FaPTGkD1M5Ghek/HGDKQwPkcvuP3yPfjO
uYPKc6LxWF19d3QtYl5VGRrhdCg3Xk8rbhKb7NFYrXi7nZOZoXerjxHA/kpESJ2LzIW2ls8hfeG/
XnRYEPRx5ucv+FOaajtCS+rGIrKhSnEGc/EloXsgAjNOEwBtqPn9FjDaLm9vnUAS6f6AMTXWHuAj
g9AFUAIGccSgVis4TtkfAYQy9dKJpEnlh5B7MOEYslbD9Kdt8R0cre6bqrEArc5Kgylen7o18MZM
2VuVa+KapuOQ3XjNwkrOhU23UANmlBQwpQqDK+ucytoKJ11mP599xZZkdkSI8I97yONLzQiY/wx1
LLOfrd6Gc7PzugFKvDJ+DmmIZvaorRYkjPCKjzKS1pp94mSmMs5P/TDV+XDYyU8MjFV8boN9cWAG
I73rKhXvAkBVytAzO4trRjWgLRkEfjh81SE2ixHRGVpJgcyf7AmGg/q5PXWct+O/vGcFIQlcP0Lg
sEFe/WUb3b7x2gVm87sLATTZE2MTOn6pWDCbzNp4w4TBgFUIMIag0U7AxXvanp84fUeS/evRW/U4
1fNiErqYbA2rKE+1VCdzJJ0TZJgxyVa443+YYs2mOoHm2dH0fnCQ4tjpmhahhrqfA6p/+bxE/EK7
N3UE1gWUnCol/0DGHIsjHChqTm6FWtAIey0HED6j/mQgwjpVoIzDZhdo0EYLpDIJf3NJmZFdtC3v
qZDoLefMYUQUz9Qbsy1hIHKvLhTaDU7Xm4ev0lUwPDVz/wzLFvaa8BFsqpz0Vq3Ek0VXIq7bDtwv
njMVw8pDIDDrqF+KvKft7qeeZsjVjQgRWTAaxsewjc+0W266O82PyFlO/Vq011rH7eEwLgkxpqK2
3tWuVaiNOiac+WnIXh+nOCRcyoCTxrwOAtPPetF5bPOvmJ9uLiajtkhOh6OhF8R3z/rNwbedqh7Q
B4DuHII1vQ9F8vPchVZ3UGbq9pXK9QzdsJoKtX1mu9PKPnZAGl/w41Td6GauCQeIBLg//CafH+Jc
YIiqC2V3qjE5APnVsuuGrx7udm3Zk76QnQhxnPkjEPnWfZDROS3hk8Z+hBUzPwRmLzocd6S6kVJx
04rJOb7s3iI8BIe3l0TecAqiew6P9NMEd4xbHDIK1aB1myKDOoE32xSfTpatzlHBxV99dhxoH7dl
xa1Q3qPITCzHSRrLyd6ZZYX0ha/MIfpd/B5IeuMCyWNBICddfo4SOQBJbs1XOG17AtS+dL6OiMfB
zMWtIHuN3hfKrH8yhtlLOHy0m//VomtwA9V624BuKNyRw8spX7QVgBFg4OCWow0x6ZFrX3CZnOtZ
qq4jNg/HRU1NTGVJME3zDh43m0AVIj+WCW90HnRYkHSXTP8w1Elm2BwOLmaCqkt32oW8sc270zIS
v71BKJ/V4bvV7HmHH5E6IFbBoWMRJAhjuqIMG2p3k3APib7dzN7+YdYPTxcJSTgitRpUwURd7beC
sve9zycSftv8oA5aPdGrZ9DgT1dkikoTrbEYDDA5ZY9z/WFjDA+kFPBjnHzuW/2SYUtEqVqshQbu
nSaPC2GTp+9wznzL8Y/nNVcJJHNqkHSwrw1ao+OYEbAd6lBHexHVDBdRCSTzCvjTCQe+U/izjT7S
NFxKO+jkLnLkD0cHIOUJ6O4dKx3mmcV1hcqy6G37UleIEtyIadx4jV2ckNdxkIkQ8ZY+YwvgL/xc
COItnW0tv688wpWy03KJpAw0YdaklRZhyDXbhj9UQdTWQa9NrNuzRhw4qqDpTUJWijhsfItohFY+
H34PeBqZbKnAvjHE8DJydv9sXcQwlJdvpicbPKXZ922kI1Jfla5LFs9UbkmUzAkdyQQgZEbPj2+7
nOtbhNqhgcUPT9OPEzZJgsIekRZzob6KVzjzCZFYeYq7KzOfJkBcGzzfyuZpKoSGez8b8rSR6XZ2
HynRVJa6MerMXKdI8ygCJgQdXGVKNqwyqnF7xY7liLI0era6i/nw/i4mKxNo74B+sHabPAU3MGLD
pesnSC3cBFV077r9+7bcdGA8szhir6Ltg/ca6nkXkH5I7bi2XDIoqpop0AdeG+WojZpCCpF/z9z3
vYPgcdPdlQiYeTWG9pw00TVwdjNbcbmXHA5aHsRyXpMY1zlnwRVsbPKFsxqmxRrElHhm9js/boMh
IrvxbNiItWBf/xmuYO3bQkLPseiZNUxETcRL8UPbXRd6m1HLgfVv2ddRFIbVa16Iz3hBUT8pLmzO
226ylrhcUXfV1l25ioVRhvYIzVDaOFA0QIUc/QdL/llddBnYCmDw3OK4X9A1YOk1bT4/FOb7+IAW
VTpfN9sMEWyH5cA90JndCsr+OGu4y83Lv3hZvR0r7ux+2jcZJGoC+83rbdXHOdLQ9OXt7s2JX5RY
3ZqLfCnPMX16b4sl4U4uXBg0qUUsBHw+ncuWlPApUunXqXETkB8mXbVYNE+he+gNOqHbPevlGuAN
YmwGC0jEtedwvu7NI7Vz/IKj1omvIM4FtX3cy3lptuWKb6b/a00BRMsjYxZZxgh+52MrheA+WCrg
AGLi5Khkt4XYe7ochAGQx84LzfD5+q1JnqY2g3emRLNzrl9mE98MxlVbNUuHQukfTOCFNe5Gg8bR
UUmQdC/nMt1Zrc+/sDsUl3sDepAAPpeHTuv/dakT8dv4K6C8KA1AM0XPU/cwd7qYmszNjgbSvilD
QUnLDFFWV4M8pcugqJQ6eW1s+oy7pcoslnUwZxAj+Y3AylpgKBr3a4quLDi4Cc7eDQzxIPtE3qB6
ftu+ADrdGB9EJ23K2mIkUsx0WDxYY5QJF3pX8lB5lwFTeK2ubuksYOJ0YMrO2kZJNsjhjebJOdn1
Zkx0OvZZG1xUxnks8fQs4ENpRFpOSu0dJnp/JnkljUs7OMYGP2O8SsBjjJNEmwWtC0tCVmYwGSbv
ZQ5rxM1Cgb9CW4/JVFQZxY5ytL4boIpT7lQVqKgeapcfHDLS58VuK1xpWg+VjgA6uksBfeMZ4J2j
rV24CmI/Oo9AQrCSDvGvWB7WKalKMt8h4RK0+PuI+yM9EnhNBFPp+/3DvFK4p/cv8Bbo2HKaJbMo
eHEBfGYQhPh2VWwZkz5ckXMijAziIEVjmfXuV3L3cvSKwyf01hDisHroDAtBNur6Ji8Lxru/t74M
cY0zwJ1VFfI51K+POx/AFyB3S4JOfZTT2iRO4XgKWlD69YyI36nkBTDZeGWdOi0/Og2Q1kXuMn6Q
splzqenk/UeicjkVAzmbgHqjOl9NLUbHp2tH1dNPZGSrOcCcSiFDgHZLeBVPKUHeQALftpsf8CAl
vq2uRLRI7PJsOvifMsL43zb/JBcT8COD2j9YhVQ/no11wKkmBFQxcETfgTrDio0RYzP94mtT3ha5
gm9oPmF1iZwd6QXB5+gOaGLubQxjrkcAEct+C3M8xyevvNlHgsYR745F/HlHRglsn6ziJt0aS5PP
OY74VzO7zEQi0bzrDA6RXjatbpNWnM0g+whWM3prG4mpJIJRUK1I8co3Khai2pXzf38ZHdMKeisW
4CwQcSOBlGNuIPp6BOlaYqC21HjysSYIvr9XjneH4kekD76OAkmkvaGRpO30ucSrj/J7UYd9IS+j
U+Pm7bRkqP0zoE62jGjLOps8+1Hcv6SsvsgzXWQCKgp+/XLjK4n6VDwIJflyWQOf6cuiHhDYNwGh
+sGwMxivQm/47HardNjNbL4ECSgKsKzEMVRk4bDlT0Pv+KEaTB7xbEJzvkgAabQyi7jUcQ4SZhzd
1u1mklH2rO5NUMX7sXfYEhccb/VThANWmFOfSGj3X7xDbZuPtjNZ2Y7w33yjeVUhdJFBXnB6PpSm
O4pfI/mKWFNFgtqshoAEYUC+WELnXpHiAU/S+x2D1aeSMvHI9qvR/LkwwL5oF/++JhO8qiE0Lu8w
KvmpuTR3ePqbznzBd/E88tlYzCV2e/IK3jIi93g+fCfroJJUNQiPKQf0CTWB8qIBf2fLt3HRCIDQ
+H3EmXZojbn9DFpAAZX6F4CA6gdbIikF9/e/ScABVyoiSKlYX0/64+r0fx28H9ohtoOVGxB8fEtu
RHR0+ZynHFWPQEx6znJdWLTPDBnTZwmdibts8o5t/w8hS4y/HUdLFiVm/3HeOwiftK50EEKjvxEg
NrMqV3UsnQOPB4UPPpiJ40PSynVcOfH3rhC4Buc0OVDT68Q2XgOv/xXjZIfkxKEtxUlAPCdzfkWs
uh8Qn6eY6Fsda+GwM9CPF88ygmWStGcZD8ELgBRe+6Fg0b9wbFaGEFMIkNEdfXx6o1x6Uli6GBB5
w/X/XQJEBYmo3cc+7hY+SBDPh251RV5K7+ayVL9TQ7pVURg5Lr+gOK7R4aiSQdRx7Pk8Oek8mCtm
424L5XZ7NMQO+l56PtdQmUb3gu5Q2ZL4dNFwBzy3hSwu/b21vaWi4WvFLY657mb7Y6ynVxXvMuFI
pDXYrqbjG+zQnxpMf94fLNdd7TK7zhTu9rZeoJGP9ZFzLTJugnEGqECyfocJEumwdSQPSjr4BPS3
a/xex/Iujbq+GZQjUhGdJtYlKaF+HWqwJZozo/ZafSoPqgflqaSIFB7vjHnF51EqEhkfn9PgwNJ+
dJxKhhX5Zoqja/KJNqtpMV/wDPAEa3jWFFC8GA6nGU5y8qIEaE8owNqHQB1nMSSa1YW0yHgOGxnJ
djKnGj9WJXAsmRndWfPgCZdVNFGJCsfEtTdgxwFPxYpJssmxOnnp/V4hwNEmSimqgx3pW4BNkvFn
NJNXd5hQaRkv+iCb+AxZEAeMe5RmzMutQ7zZiwj60gKU8jHIKWWfU7MK2Iv38hImXf2kihkkSGTr
c2Eppym61v77Bu0Mp7huV62M8lQi5Pb3AwV1kXzT2tgiLHpvQtBMNFjuD88ItTjd7iT7CVapfLyG
0Y1LxdImT/lThqDmD9f8CN6yhEbwTujQYBXHgMpJQYFjiHedZOYzhYvqKrLDXSruZUcWtY2ohCC2
Q1x2nbtaCVEgCivvtP1H0/IPh9Fubwg3QfVL3aQc9dJe3eCFS8pr7dN5O7qri7RIVsaTebX8DokK
M5IOIRaP1xgGD66ReN4a5jfEXCsx/Wl2QX4RBDq1l+kAHFIXeqzJza+xECotWzbjqJoXZ15tFNkF
zzlystFAfDmXi0CCQJB+KrTjHjYb3u9G6ykR86EogXGEUfdZv948BaZZdT7ch51DbjiurfReD4fO
XGmbcGK9VFfjYOTmflcqImKOr50hZTY7YH2Twp4GnrIm5OYh3/27FSVG8yefeCy3E4iRnMcxXqU1
ofhMZXnnyz9WGJZbglkKdabdbu8pEWPe0ZGNcu+E5H59PUciO3LpSzaxxRRC3kA1vKK7SmjnUyY/
mna8RuxIq1QvL4VNxpCOKFxzA8Tvg+fTwYEjrs9l3u3tlbUpprZMtZniDu8MUW2XfAdVl18Gxvu6
RmQN+M1vO2mrZZp8meGL7AuRGnS49L9b8Y2FxrQ1U2R4FJz/6urtQRbbKnbiFMuc1CLgy23SBmkI
N5GzkWcyLuykCilBr22WIzVq68Z7JN13YkAA7Muiew7pJM1FV4JxHxKjGsfpyOurfkrzzSuWdH+3
IiaFtxvotLfnHc1EUBlJghI7eXaO9IEfI8vXwRnzKul4a2Ql07kLvCtVlL5IUqNCxYjb/9N6wvGV
az1nFmSSwSA0wkEfUYvMrU79kSyU4ghqwezBfzHWgB/Wo/aFdEIbcDtwjKkHHpFfcEI/OFZvv3xz
sMGwnOqH+WZ4IM3XD893r9YaLRZUBV9amwX49klDIjIA2GwTwIZCClCcSaOjTFjBS5szNSDhJoFG
wfJcbThHa5gTjHd6WlENyOQKQgencxWdyUOfaCf8FOQwemcFUhbb4+c3miCj10SbOEbz3oetl+BK
8DXuv5xSUbBhR5BmSaMTdkwMNqCLOaagKUwPRtvBkrCUloi5SizgOw3Y8mKRVpsL5BNeEAPnbFbK
y2h6szjKZ3fjqVqdRUMe7n061LUvKOVrAnB9dIiekOUzBmjz1JXz24fKn5gTHuwf9NLOmzgXQTDH
dcf3l3OhnmoXiG6B78DG8OXNoCEHYh7QYVJRecoBQ7/D/SNHicpSr5EuDvmvHtMfP+FF/uBLxtC5
cya+D6QH8eX+qGRAxEowlbYsLY/TCxEOwQpGwHiTNAARxqok+osBaFCM4NemFdWMaKzCA3BcFZWJ
zrx1m9O2rOESioP9aK83xns8WMI6nHQa+ZSSLTW5VD/od5LFSDuZz8SdY1I+NqHtTjgcCeL/p+Oa
087YmdEfLIB0GXYdjvR+Rc1/sQsXbwuX8boQg4a0wlPeU6uoERiNyZvx2TeDmf+Ky0OlgQGsPlau
uML/RH6AdyyRH0K0Debu+0Wcvwt+32Leb/01ohx1akL/bM64TzukH9iSYf4KCU5X509xYaRnX2ZZ
NK76yaRsqs66ZiB7YuuyuDqy9Ua4sPUGcL+IEAp8SCj8AaRU4+3d4MIU0I7H1RKF64+8d4tSbmnD
J/KcaDqoiozd3qufGZMQktcByyUR+mheGdN9sPGHQUCwh6MroqwWGJ1bUEC9E7ZiC1SaDb4UpE+b
jTXSCU4LUKV3HOy1cIMeqwBAB84Ke9BCet6EbgMeiK85LnL/N+xQ4rSaquUg2PzNP5GQqxZ9tmo/
VkfKyzyBLi22hL0kWH+JG6rXfZpoDJMVPk5p2U7Jt9mvN+jTsOzcZiTFzupzdMGz/nHpM03RfnHh
f0qWjWVOCET5KCRfA7HpWSYoCHmKdkPHz1OpnsJPbS3bIVpI0VFve+fN0F/5qrfbsIuHIuojXt6i
tv67pr1VAKmOJauj9LIL1xdub6fGFEWtXwSgyU2fhJ6ZQQu6IUzwnftewZCND1sSL/K1ul3hzd5u
JEbcpxVK6lyiw4e7vRNSSjp5uv3Q/Sq5ehdVgOrJMZLWgu/Vw0hs/HNDzOx3HMw3giRYUGx62FGj
+a3BDEX17qfRuSXkIchSB9jMgYMaK748t+sRFhj0ZlVtm6YuS1tdHfHf3cbCyuAwLBFhw38GmQuC
OmI5EQ5q0sTXHlFsImb8JC3sRDgpAETB5JdCkDGeFNKAly7h1zDqIvLrZ+n63NIab7oa/fF55gJB
zFFAL/vDQdfBsY6gQAjxnyMzAoJ+B/O7ICPVgMIxaoS8FKLdfoJypGKU9fyUUcSySe8nE0lqK6Rv
grcAIy3Gb/B0dHOtvFzAbBQ91l9x8+uWOArQDcaN/8WcEjfHhiCODJfMDlhRXTtrYeDGyDWTOImn
9/rAK05Mw9Tb/YWN3Sz/HHGbMHGo7pChenTxora1cU0oS9w35LAmgXg1/rCmRZruyv/HApvzMbvB
S8RG9PlSeX17qktO6nHkpWYMVchXIi1oadsqTgwp7G7HHvdST6arVZ3CXGWNZ+7nJ1L19vW4tmN7
6Ho7wIQbsAFA9xvC93yv8dsex8oXXShgFy8Fd0gNjeqIqWWulLvuAbC2HNSgD4HAutB3mWPNR82/
TvroB98xUVTv+UEJBF0OUZF6PP513x+icjvdwPjaRlRwP38BHyVONy2UcDbPEuUzv8QjltUlsRd3
szD+kKb4+rM4gBjHKzyzPMsS1lB3JeOtfLrzoTQsNcKJxBzQZcDez5mDdMV9IRiZLm76wdmU0FY5
th44GfZSoY1VSzxvwbxQktaIIblvXR5LGWtYUqvgcym1ZnT5+XNbb7m3CRlsfiAAdWVx2hU+DnIn
NNdmVuVTIN0vXTvQo+X9ufU+Oma/Txfx8XNKu1AO90hbtplD34T59NW66z7WmrhcQCoGMtW1C6lj
xJ3WCA9jYZaZ1YYUb7zQFlgFccaSB8d39jA/dlm2C7za4FnRApTa2hq1XrRtGLPwY7ojC0tIUkvX
q2ke5mCBRkOMub14nGuivYTPrqm3+LALHgi8ZRdj2ul6iDKLOtdCnbsp8bRM+JxG4LK6SIzNFEYZ
DWtWB1PuKdD94tKP7lBdmL0+m8dKQjVBcbnqTQqtQT/FW1kkFbp9dHmPjEo3tYHdQiQuHstBWjE/
cq4KFthP3O/n5RELdYwPnw/LAca6FMNsV/27mjvYBp8tqphGi7tRNmBZkKWeu8NHs4CXjiC0Y2iC
7UVbwR9V5AgXjQGkE/6uoHoJVgp8yUJQTQUfkvl5I53EIbG1Tn38vDMlXjWv0prLEps3gqJ6oyJa
PIrwlEmTOktJpryomrEqrLEUTU+nGiZOk5gs+/n5Wn28q4y/HM8dv37bU4yvPgCcRuukUuubHfmY
aCJUs3d4VMze3pVWu3aWEX7y1vp3N6f/1tMne7CA5ibjz5Crkk9ZhUcLcO/max8q3T+tll2fX8AY
nm0deG0L5nkXtPfyyGP79+uF6jTHlypeNpJEIJKLTlD4n4T3nVUWP9Pm34HZRKWmNANuaUjQoy5j
TzPweQQNRUMYLcPM0WzY8adMTXYfjxEMUjCryqCxg4xdgoxwLVw/NgiTmwftvyALBMxedymgT24B
1Nw4ypNJlcqW6KtkKPcc5LeSoZSVGfF7zZeagj8XIdbI2zB2sCCY13sU+8iZUhSpHXXRvwA8AJ2Q
mm5L2kRE/dmtUib9Mw0joA1olVFHScL0XIvvmr/pem3kWAW73UMEsKBgFj8lxjj+j0or0zsaYdBL
foddG16ZI6q1qjkFr2RwlyERvhN1PfN/rIORYylh90XPCb1nrQsBOccpIocCAZArXgwr2AwPkmnD
VQKcKK7jQUqtwsLyalouGYq1uiOP0Okhk7Agw9uWOVJ/fmGuWx90frAs+6C5pXrzBYmRRC9IAdAn
8vU5K+emVzH1IUuQqe1UWnH6T2sJMG0PmDTThnnGwS+0l8xgpR5OEa6tcupQRoTA0gM+aWAmaX7L
a8iV95tO8AioCoVHQIzl/zKi6C1cAGLBljuGN1CjtMcq5bhYhuU1FSaOPmQQNJFT4THt891Xpiw7
Ob/2Wfbkmug+ON+tsz7VLc2770TcNDhu1Xcjz1ls4cK2O/cwEMFPXwF+SeDk1RTAmHBR5uL+bmwz
afBb0Do7wJYmuAZbmR4DD/hirBoG2DQcOiFjAVCINPayEBJSj/Yo1iK9YIEDlaGXxhfWBaK5xhLW
dwg1V70CBpyPFbM7bHk1//9wVZsyHbZyRnHQmuTWvlhuv072U7N23b7ZH+5xlg/UfLb3tJVEULUi
h0ffU27mcBf8OxooRyCNAUfJXiVQjs0SaLH6pdhAseMND1YyDauf4LHkeWRMj4mSniMFliJqJ78A
CVvUkiqiVcud0YxbsbaZCQgr+bPHkZD4jc2hc6BRpdJlQqLnjlJVbOmNMVnO5aZuSePisGCEl4Tf
8U7GKNtF+NTnaA3EL62kcGt+TAx7HfCZ8dnIolj40S6rlrPcLG3FrtYWGHCO6D9Fn1ACnsChs4jp
w3YrGrbK+Bcq6X9DzY4jMeXXtFFr99sx9ig41h+wHXevdXH7gcvSIsNq5B8ZD+DydE3rBBmapbZy
yH6wnKEaNFT1BVL3qH66hQdapsDvaw1LDniiSvnpgfEdnlsI32Qe3ul6gME0nKhyWuSTqlX6L6dE
8qPXh4+NbI9b26LmUpcsJHjzjwDkBBZZMdUq1b6PfLTXguXj23pSH17j2VGXWaN4B59p/SesYORy
xMu2611QiTVbkazZPRo+1/fZNAeLC4Uyq7QcWTnvpnZdWYYgwJWYiUDS25UOMyInWrt7dwocsSQe
AR5l0wYH8LhpCVyyt31hLCLe+xbJv//UJJv55FEGi5AQREiouQj6yQNy6iq0Z3TOBj9DoZpq9Nb7
7ecYxCm9SWA9qA9SKTZUSnYefkZVTOnOsDT1C+Xzp+HGFmelFoVl2FuBAgyQCbMWxeDZTv5RiMoy
H7L+ukGo2LJDloyY6KpPHH+LdyxWOWgplLfWx9zosYupS1LKHZMohrp4WI79NtZ7zqCLPCo7PQnf
ko//KOCTxMsOUolkB8gPskm96ShIQ9RFbLlqPkhP1NgSK5YSqzVTyXdf5q0QbQ4mEFluXm8v1Gsb
2FIXFJ/h2uC+av85IStTZ2tsU2Im68F92I7Vwp+JmeLesC4yMb8MeZJKOEU6ZZ1CmEORzP6Z59Js
jk63CuxDGjRAY9i+1+dfPABDgFvph5/fnKs0A/Od4OPyg/j/wT2eSIdX1Ktu49PSvfo9NXXb/fmZ
PLlzGSheJowxG4bsQdePaOG3ThjlDBRfG6ZFc8aWrdXJ7ur16VuHhZoBxNiDewQHZKolx6ctbe/l
+//08lZOon3PE1eZ4vcsad+vBWbq6e8xP/gIhSzhuOod6ClvOBzYVmsSqDmhwP+nKnV986ut6tYd
/asgJ5SSW329H0GaTgGhjHg4O1nA6wxNgL06nFwxyQx65UOaPjwWR+6IeMDT42z8pwGsFm4a1D8d
BQk+4Bf0hTs0Ds1pf4xxD1PyH/YmaeAwUu+bWzWaN6RGfx8ny/Kc/e74FIkTFh5IUhnETzzF9Vbh
f+sL2uSQlMClhbPceYI4xGNfjzALXWUCFB0wmd7IwXvdEq4AVsqYBNf6Du/xPyrgg1EwJPrK/xCA
8n8Uo2dEgbgmFPZy/grjyQBeLfavrOCDGvciFHjiIydqYB1S2IYLP3SXQnOQ4ioHqkYmqdzqWOpr
K3PVWtJujPoH/6lHjRaiqsx806JVm0XPNGT8uhraZh91MOiiCJ4lRFUsgDmgCz/oow82bq6rbU6v
GVw0y6noibG2x63lnsTUGi3GCRs255gEki4dBCrotQ+EqNkVD0xlwmAcXPLrH3Gafq7bQCKtfhRk
98J3VavlCIwjZ/qAUPQ+j70pVaPZS5sIMJYrZSbDr19LC9LQt0/bZOkqh3lXxch/4bImpxsux5xs
o1AqIzA1LZ3XOmniHozHQMz2o6FhfRZtCCX7zGIC3MMzYB66GTfwVSRk7xw+mSmOkyxp1ocq8OPD
iYHr4skh9yQhUynQiUhhf4VF7eN7fPqtGfirl7vp2jdIjo9Xl2DdhNCnmOImSwbCRxPYzHZCGWNe
aPhx2JEnZbiJ3mxYE+VVwEGBt/1XJDucJJt8TH8RTFUr4ippS+4W6dSTJ8FsxqU+ThdyXptMxNRZ
uymkd455WYoBPtMGVq5kYm4fjHyHbcfvGVEONpFgs6cxW7+9/dywW4M085Olf2IFuEOKRyE928nA
jGqKXmh92FamyDuZc0ywtDhVYeN43mm8uikSWD47A0ZBhks1AlrBpV0ETPuPydhFoP2l3FVKBc3z
C5MJCawh0/TMUfesYU5cI6stMBK3YpJ3qlAqxbXfANdARX2uEQ+nV/2OB35QQZ9+EAXld2cYnRlF
kwDkPAj/Lu3A1wgeLvBUilad8E9LfuLZPuThh2jBtCXL+urof5VQWigVqPJfTizmOm2uMkXKkY/B
g+BBU3rw2TCVVTVY2xWjg9bZtJ+t/oOXJKhTgleUWs+nUnj3Gs5WDN2u/y3Hhwb5eTfuV4AMP5Sr
pxUlSvAS8pcISlmL79op1rs9WyCbEzpCaokPM6MVI/QBQpANhICwx0yxvWloyYeMrTGKN1mT+hap
fnPbz0KCnb/OcLOIhz3VyxL24EbJvOkKa8DFUx8xtBp+lW2tFIZ1+zL2yNDVbqRRPQCM3TfSymxF
CEu6pRYCMhuIx2NHa5rFiE0VoXBTDb9kPC3E+TB0vjU2ehufWx7bD8F6/1t8PfSxrB8xoEH5q98G
gOg/oYP6zTsNsFjERDa5WB0vBzsGRGGSPIxMWRhE0cH5EpKygH3ul1Xs9la9Yk74xyfhyE/CtPfK
EVIEW3tJ8MH/kxqZb+S7OxVUW4psNsH3jlaTL38Topvf9IfQCKYZboP9PVYv+4hScNBGEPTYKabG
0qjqpHL+feCoNavpXOCU9d4WQhqqo9DMV27TMxhw9Hem9fFSSy/dPKngu2f6yaC0QrkmmfV51rnl
huo8u53rCwukYEwacp0yseVmZP7T/ckHDSI1E1yXrK7h3K/pX7bgF+/IuCRCnHu473hiDiOwUCsq
meqNuvjXREHEe3GTBiWpwAM7HFoQLG759wEgcNDKEi38OsYkfc7xX8LzexwI3RAY3fZ1dIPy46i1
04wpJXefRuOkRcRhmDsanWopnB2JZQJ4u/sFRDsuH7HpQmp7nnMLql0t49FVJKny2f8EJ+6d/ORI
2a9W/aaPYk//PS6zSaZ4sVuiPYCzSctVkMpct8AVzlkINB6z07MgXnmdjw5JqL375VA04KHykEqz
ENaiGiZbwr7ebwEOeLh+StEgOtfbAxtJFSItfRRR+q+RdH91TG54t7G/X3bDMJ0KR4jc1ylLiGnQ
9MzRE2dijb2n7GqW1kPK7+kRxNrZje3oTkEQTIg+t3BdbXVAIsEP4u4JYseUJcUYL/MZJ+jqn1BZ
4yi6zituiqQ6cu3pgo3F0o7tbI6hFXgiLjrnlwbpRftmSxKF6AGg7aLniPC0yEsR16YWgZCW3S+1
gurvzFL+ITmsmpYcCi2T6JvOFVFSPhXmxyJeK2Mhhys53ArCNJnyGIM/Rz3oASIm7GfTV1Yj1Fd3
HabyEors8YyzixTDzKpsgRh70+OQiVIe5r0FkaYKhPTgapw9rg4++fuGmb6av3O3w8gZu20BDV5n
MoeIaQOmbEpPUbtpJX+f9WXPSc/35BR8+NiQ6Vyam0VtOZzydRIYti0TrUQdzIVMR5jsJ6C27bOX
TJ/2MutR/R79NQi0AXmTxp0quKdyq+8r3955GSaLXUMTWfsqO+mfrE7XW+Yxf400/6JTjhhfecsz
p9LyQGwwX6Sw3T/MUoDCy6MzoBCd4EDqggJWreBwmmUgXvqWvQrEYaQ7cJ0oSbCdQNPOTbTEMVPS
7weipA1+BbX/sspZZNlEmKAsh2mydCXLPOs216fovee62BxuPuoaCOlrNHtr3SFUAoCtuQmaavin
cam+bQK7RcaTJsYuCnfRWXK7Zj8ft8rY3cFP9ZRdY7uCp19cOgi8/nu3GeROOD9dshVlF4UdgCFt
OX3TGAn9HiBr/9FDi7endRhN+LH+cU7r2FlmobRprXKKMjIOXxqucfMMAln+YTZ5YYN71/7z2ZjC
S6hLsMpufJxZM3aH8XJA1ExZR94muTTI/SoHZ0VlgPN0qOrQCNoZArvWksyaMkQfRG7mcSnNXlvm
5CFge8ACmSm89My4Zr3zXXmD6Vd4TbXqEKw0ESaM27LIKEAWQ5qVk83Vf9dd1Y9+D31Cr/wjpDwo
ECHqcP1EV3JpBj8Yh3+pZr5vbFYq3J2z6y1Ack8HfyT7NaO/PUdsErwbSXhjS7Vt+uP36NfJcu3J
drE1M2rxd4wxg/45CSpqPG6yfbVkBWR5JLJhwOthZeefQyhTEekUx0EHhcU8OpZdWOYRw4zNXp7d
gfUNgxPu9CPWufO9DYIHsRNLawsUdCrzJQxsAuNqTzkEUTX1FfcTEhhMlF/POByPhQsbpsKOFXq8
aWgJRT3S4YuMeEngn6f5OEglcj+GXaMVyE1QzXZaDwaI1UeRmqQ2qUQPO2FEPUID5v7YmKt+iarC
BQIV01QxbCp/cqM3Dicx+RAUn4lBUc8P8Va5UQiXp3cbpQiCCO8NvYnO/FoYTKoqWgpN+OXZgJD4
iFHiaEEAUDN6uaQ9Tqa55WDIPx6McDG92UgV5W+t5XLyNFxDUgXio2DCgJTrB80qXAgYzaHic/tb
rAxplurklABo/Mo3P9ChLs1q5BHXj12Gd3/KQ2il1s9ub5qSNUNYas3y6H73EaMvyOyyesJ4Clwj
+PVMLWKKsaX1Fcox393xmR8Xi5Y8L5L2vuuyHQS7W79GM4hS7sSuQcnpPDEmXQ+dITgHgBflDLyf
NtSaW/n1HFrCmOu2YbuBxORWe+5VRIvV1Ry1K6B9MpoGq6fg2UvLN8h9s9kkoxsVCQUx4v62QK9U
xJ/Pt5zIy/agJVyNmaDl48oI5ZLi9TLD9kSF3I6MiIe3jyjD+snBi62jcB0/OzVOPjbo+nl5r/X1
TMW5D9Vkbd8680ali6i+kwOB540VDlE5XlXPT35EQzbEyUCtZI3g307NY349esQrWPwmKmFL3I9U
EsZ1LCX4BCFb5fKxmS0Hd0cJ84MdmIVYmnY1c9CGAoNAtf8J5UoxebHBnwkOlSgkXnw6YZvDgP7W
LrdVNxb2SnIgMreD7KUYiaQygL38AlS/0wN5gHwhxcT/iAiU+BPCzYwjSOZt5bStMUl9g4E+nxSX
x/Ohc4Bk/YmOGT/7qlPjke58LUcNTnRy4W9bGatKKuiWyffn+UqpxocbC5m1uWW4a1SmyfPgDJWf
mCtNRddSypscM05NUo73W9/tFnoKfDFXtd7wqEIHNM8KVAm64ZZLm+wq9OJBQ3dfPLZQLxiRknK8
pHyhEYMWhAPYdt6Ln5k/Ljv9IWF2MjFD1i9UFqM2n5RKgHg11FmN0QTn70WKBBLRafuQAV4JP0mH
fqX94nbVosGNBArXM3kvZN0JPBKJOOKX1Sl8w0OFJrGUTjowmA93Ud6MeCuCjh1+kDM+r3gOb6KW
L2OySdtJBtWa+TDfyd7jXlDAVvvQFVX8FqkYgLMZETzATYaN1udB9YAyxg0YKcoJlYZOFG5o/Y4i
uc3S+r0LiFeP818KXcEZRjdu4PIqE+GOrhnNUgBStX4rSvlS1JVh0y0e5Hx9jpZHCDiMbnlNESx+
WVel88EJpw8rC/Eeq54EvEma0mmv7jy7O9oeU5q2eUt4bB5iUThdK0fqHCJuifg1IPE5CLL+ELn/
2W2A41LBdvaUDHKUlXVMD7pVdZ8yGfh+S6fxksiNvduaQfHvKtNWckNf77fy8+m8b6k+5fvrNKW9
V1SWMKoaVeOKADss5EZtjE+v3e6i5Z+xVShS9oMdqV5qMU7Nkrmx/61pOZgoBtqu1AKIicAbfvVH
w8aZuwZ70Elf0jH2eyOttqh1o0jTO2MJfwGB13qcXE+94Xqke7Cb3enKfn1EQ/+A0jbkS2pcOhba
SeA9SsM8mOq4lcil4JiUa+tcomEZMCjgIMW4paadGm7otuNp8NKAXNJdsvpnMFDBBse1K0Pemr+3
ZMGfC27t0Cpq1tfsjYouvPtm6n0QdrPy2NpUZmgmFuj/dFraePSfiacB6wLdRlbhuaR0JgCjrkNh
7V9NivGO5AcYe/14TWd+ntakfpZ9du5yyYuA9b4jRDXqXryDKnwPF5WC9fGsIXVyEEURRYBG+XPB
HNaGPRcaTWaGIYfLMYcYiLA5QFlSNwWzp0TytS5nKtrJcntH2DWQKP5ASvSxmXt/6Zez8mQFU8WB
u7jk+gTMINyQe071yOCy7v7/BNvo6KGx09JVF9GT7GC4EiGwCQtVYgSjCMuISa/fm1e2QDjwHRRc
KgRzVyFpmU6RovtD+1mbzEw808L9KcC+FEvFHUl+0eE0ZgcqvCQFZboHathp84V6xCtWV+GUHL+C
oYiyfTfpXiK9dhBhjoagZUhWxW8CJxjg4rEGUn1zf0CKueyO2i2I/Vi0f+mDqW8zbJYu5DrQXu5z
eZNcwESaNTQ9nfsZpt7fWYox4fpT+g/AEEEMDW31L5fQMZ2uknaqj83m9KlI0iyxprvUnEwOclze
gccytUjhLs58ohAbRmSIgKyILQA5yRLHKRzD/1pOclUaPN76gMRuBuzCt9AlfaGRdtMzuhAeCb1n
SCzyLYFbwrpRJ0SDgF7uzfl51f691CeiJA22VHvgHpn8bNKwg8SPwySO3qMgILq2Jt4sB7zLlcMx
+drH/EObqqpwoyFOZAQfmA88Amz5WEyHYdmClBcq+odpFb8oJzjVS0FUuSDQSRo0H1hCWeEz96y8
Ie9UQbCbWNXthPWyipNpg8NBOAZ7oR57Jk1ehsGwnqV9+Q32eKpuKRCkiMnSdFdihdxfg+MdHoJD
d3w2eunZgFp7yA7FORTH6cEp0RWBNHudg0eiOzxA1/u/QZumwfYSu7BL+uF1uz52uqLFCEGTXgZB
7QyuMBFCoyGjCk0CdgIPpCu/IAEK/AeAvwvCNlzY9tiCVsjy5hiWveHNoOuksGN2oZcfYJaSNhX2
ZSC0gPXXyl0a9vNpIJIwOPLvZWEAosvkEoVdI4RhttInnj/fTGXNWzFFJyPtiyBb3mfN3riH+Ema
79C6CwppX29hgZbbKHXD8LaSgGe7DnAwmd2iK6KnLP/UVFoEgxYyoLAqJzxhfs5cokTUtP46CSUU
QFLLJ2DfSSyiLmELw+GqRe0KPbZyootOdId/u9ZV6+jiVCUrwJfH7htD+oBiujiulUdGpi9Ts3+I
sNIDsXQ46I6Py6kdz0/Xv8ZsHMwjYdsJBMT7XwQPqNUcuMS5LCnhmBlV82fPEdkkf8I+/1kq8wGp
D1m9rvqrkpk+UvG3LpuEw4aEpOXJoe5R7ISbYit+B43Qjen+m8L1lizDPg6PJvPWdkFHD5P/7itu
RNSkquXZNwtTsN5fAKW56UQICFpmy3k6wUvMMIF/J79WE1BcfzPGRASG5G1GIz8ati+tGog2zuV5
NJKgZRb3M/xRs9kGxhM5phoaRgKgIJubAX04WBDp+lE3AlBpl16EBJTTNjClu2jWCfkNlI6WHfyW
AOe4c3Fj4m3UZs3FpA3CDhzkNxkx5DlfM1c1ijVSd63mGxGIyhL0recfdH3ic6vRtOXa97gh40fW
7c8ocEXebPtM/FcbMHESqPyvYkQUgI6cjDV/XNEa7rlUqBbp3/RamlOlB2bWfS6p6p9ux8ZsuJh5
pLGovYNJPfxrEtS5HmMn+6AQjp/Bg3lvMTYu8p1yLIXX0URi2UXBQXqvkf4qHaNJhMAJnhM9qEh9
Y5rW5Xp2QfU5HJT418bhXE5S1CpAxD2T4B+hltiZ2rKBaWczoOCiwNfx+PsON7K7gBSVS/42sOQn
/qL6Wg1xZ5hMNPNwl0o4e7LvQSel7nKwTQBOvgT1ZODEDVwlTjDJdvZ6ZngLlBK7Twt45svFwtSW
+Mbmof80y3IcT5IRSQ2ndYSe3pWsp8wVPAz7MwN4H5rVwLvMgofV3D6dLq5cJr/2zbm2z12PlzkL
29pILbZXqZMp9dw4REHcRrBdTG8WMmxGP4l1Ce28FTWWd7iOPLsaTU8hJkqfbnzTVWAkcoxeytN1
xVuC37eJoJXWh/kDR/E0EdxXSgYSffqinSWC5vMAEgNhObGqqxDeIwRJamzTcZ8rXZfdgJmw725K
Xvg/Jo0E3HHw0nCWwjiw5aI6A5T+drZi9i4nc+/uUoztBJ9Ls/Rg++BEzQ2NmeqaIbNI8KH+mnoy
oPxhpKgOaFg9JCnLGfVfnUQMQ/c0eq2XK5KdcEwUP/yWFifPNwxKaKt3uOQ+dE61cgPGZC5VVTJX
rU519uKWnFr2tw6bj/CPfQr4ddjioFhNNuryx/z56+ZIfMiWg21c4evqHT6r5Hm19K78WLbbrzdr
qpsurnth4oMtvL65laCBYUjs7U8Rit6Yib/g2F+LhYdLXEgMZna14XBRzcJ+jgw1tCcgc2AWqvTK
9d20EQZzG7cZzXifGtZvoQVZ3BHhLKCpujDYD0XOQjOW8EHaKt/+x3P3w1mdrKNTWOXMEwM+ENsM
buPQeguT9kRGTU9TW7vy+z59UFknqi364MNIXtSEfGL9BdR2liNG9w0KMt/N5P2ZoJcU4FN5EN8R
YqKJ7jnWYFlEKWw04YKsOCIezAsiUKRbBM8UFxFBUERf25zfSnmY8U8ajORftZWHDWuBjCx1uaA5
WQRl/NqNK+OIL5Ozq5gSeAT32yEhbq4a8JPqvmBfdcXFdEVpRzBxuxGrE4gFL/YWkYdj6fDpOg0p
UCrST+FSHt9ht/kRQwE7a9DqAJDdZcOiYSvi0gb347AxWiFIpnp1xNRN/BkQuNvAT34JKYs+enem
khCP5N+8Egkm3ZXLQkQCXKuS4kgctFeW8+Y0Owx/X7AxTZWct/a7ff7OlKHs+bZnGuIbx/PQqnjE
V33tQEZiB8fR2eWlri6YyCbFxJk1EMEwXMk/wxudD3UDy8c8aKEGdvpSzqqWtfQbd1lQlC/5Jaa+
ur+JINkixU5Ial1279WGV7JXMBiHIqVne91e2GMc9wpmMm0KJ8ADBPOw5sTO7gOfHPJtL+1I8/6T
jDaHAij/GkA/qpA5vrpMrTuug2ywMMQBitp/DLYgY3fpF8ld61C4T84p3bnVP4urXjMAHfCzQWLO
CsROXcP+HU8TEZXMCgfxMm1lOD4CPW+nCGpDiRdABtRZUzImhIQdQVLmApwTO7ZUMbJyD+TQegZd
8RVPHFAXhyYT+1QeEnnttEVCPUTuXah6S8soerMWM+hCKtX6vkbsk4ph78hsTgiTDA99dAUNzG6i
kgGELG3cacmMgkJ2sKR7gHnozl+3MA2waf5DtR/SjR6V+Zx55pQw6m/OzXyOEJGKrrjs5F1TmoRU
holktSWwD40ycSHa1h37v4GcF/1zObknDSBdLFgnBoOQLT6zUrnizyZvFj260kFYg1vPk1Bpuj7D
L4ioVUmkDWjq5GTXkCeLqyFm7N4nIZicjESkHrJ1YFXevA+VPvX7Dq6oerxBYchyWA1AEseQzZNy
nElNkDOOHDhjcl68K7ybHrKnvFNUAzDtzLDOshoImLCNG7a5zJLAO0qIZM5NGUs4U+Pd+ixEcFfI
v+7AXBUrSrQzsPPz3o9yPmUbdPyBMklVjoiNypdRiSwvJt50S3IqM7TPG4Zw2KTGV9eETgZAyRUv
W2+/bwPWbHbz8I66V1wW+AaijdUycpJ6QCAFpTwXGz1xmEoanw40vT2skx0LXnA5O/MBN49v1ro4
GaEhK46V1I0l0KueWQdDLGPSYleauSgCWT5qMxjpXMa5YTkUlzWlZJt32WddMDHY3vu8VikJJKv3
Fu666676qsvNrU1RhEyv99rTxs4YvUT2IwUU50VMijt7hXKXelGLBVWd3YxTw8AQIctmPi7K6Yg1
Yc/SCjYSaE1fCnI1kgC+oAdmPvPTcfBFP7SXtBBgsSzovz0WvQ8+x1T7D4Z7Q53ZWzUvRqfy8FYp
jwk803NgIKTHLrxni2BXOb/o+ZlpH45ndyUb/iTaft005WGmrb9ZOgK9UqQiuFiOp80RIl2TqyPT
kaOlv/QcuTtJt66HPVZNOk+e9Chs8YeZTuMz9Uz6AHk6X9MVFRNxrS3KN2nYT0hvgNKkNY1q1I5X
iH2xdosoZAnNR3Ql+ZWIhZyaBYydMxofZrl08vlbIKxx+OOu92ruqMbVJ1tvJNHRCk42ogYr6i4S
3fSBWK07oilP82xoYXSBR05mE/aaNNBkF1oCXmEFT0+NCFdX+xbcsRo1BrNDy3r+tZn9jKEwuTNj
r3zEM9n8QqifhmgFT9HjBlgX18IKv1q++J7VHLXkIgxlevY4PQLIV5nJVHWJkbyFUNu0Mp6WlsxH
0bzqCe3+txm/UhXqD1sYp7ioNpMocS4omb8/XU9vgMXaEH3Nld4hXew/T18alxRFu4ib8kan3hPX
tLlu0GoRK1zjk3OHPB2/zQ335oaQ67qPJkBNHGsQsM9NX8lDGRBLCpcMLtyx3oQfe2Q5qNrKLhZy
sFYR+0i8zpiR1VFJqQs9+iounjF9QOFWUOsX+HS5/1E2EF5oyU+HTNj+TPJXmjIh+Gi5ySAoBrP3
aw6bWVsCF8klju8SobqZNL8mlRreQpMhNaMY4uG0g7XSJU9f1kl34ODH4Nb9xKiefCFE9XJFj4UW
tlwOOksP53Zl5TcRy5QCfswwkqvRz1Y0ptQUGj0Z4/OD1+D2I71aqKNjM+clLg8w7AoirGJOI4rs
++gm5ThIasGSa8nMl5IRp47/btflc4rUPKbwzM4XoIVhZ2QmNGnC6T0ZW5h1R3wCCBFTJyqX8WG+
N7EigpCsdI3RQQVlGA7PuFulxCYbdRQdOWaAfsuMXneGJo+EFETDuo00Lo+Q7JgFhN2+pp22gSmx
8/AnThRn8xh4Aa06WqY9HgHGA4S6zpKpYGGgPGoTdPS87g/IbGkLcoews4wZwHnYcud1QI2GBD5a
7Xx1I5U7C5+nh2e59b4UCF+f+z46iSyPVJ/ADoJTazjRn7t7i2RhvWpkmm/GZRIHKHZm2wYMHfjS
FryIEcHKvRcD0HlNj275cEduy7kZahd1M3T4cbZK+3Oj5aZfPZHDrhZ5hkx6yUSerV+Ji0Zk2K0j
H72nAbtHZ7CnyXgnlhh3z7sqyy5bAuPTDvQr/N+N1nSUqgyGZ0yLFL/yVZRRcjUyivqbb4h5kb3Q
00+dbBugp1M8L2VcZhAG6BAAYhTD6H7vCqzXxUlH7Arjyp6xgK606BWf5Lkqa5WZcztBfFK99o8Q
ptJzNHdcBzEcZGKtjeZ0wgosaruRjKJMTDH9pkhPu3cJ/3eszeBDxVQ2de28UNS00zzMptUW/ZiL
hqJB62VW7NMSexk7utNNTIxHSsOk8ymwp3BCW5y+plLfrfxDFgH7LfOSlJ6wtAIbM6EnTkUjl6Nm
3QjR/TSOx2y9P3OMUIL4XvQDdifvr/4pL2G/+HDmHfarJspYCWAILVGbkhms9N0u/vkVn232nxsk
yumBzeeanVGbLE/vUM2RA/36UrnX6Dj/yrDvcDWCIe45wUPsgGUuqNmoqJYfE+KLd/lkrUhSF6yc
HJOQkeEEx+zoXQxxZJ05YfdHhNDu3sETRPCUDrrxPcazBmsSWHeGBS+XwXo0xU6svs2uGDI71pD1
9omiwLpvT5gKh2lnpRDqzwz74ZHKgDr+PZHjc/mx7WRxKqaCJ6ASDyOtPRou1wshlx3BoF+xG1hp
K1ixzuHTwKVmdKehq28tgbp6y5eH+1J7kEVKBqla1M2OVP0b6RY8IkXAee6vZD4r+4I+s+ynrEpq
r0oA0xnwX+wK5ld6H4g+naB12ktrZkbHekx45YPwMbCnas1bDL586s+uJSys2gsZSaQ89frBHzgV
T0ERz6ZeRnJs7sOSceoYEOP2KmRAs3g1VesHLbpuczevWL1Rb5f9+xDVIrijkqqyAh00QTkKc1YQ
xOEduSB5k3o6IWXU2X6a6ZB1148hGHvqgTyKL0qTOCYZzzZ5J8C5uw7+4NkPdy/P2lywIdqN+nB9
80WxTolDN1uyr+tc9LH7KAusX63WvKN8qZMJoF0SwVQlS3MSNFENimMBuKod7Nw71feTxHIJctGP
cMsUryzifhBpqIHju394B46LUX7cyjY6bm3Xl4xb1+rrZ7X4sfPS5CbLLTs7xrjfnsdpTPS1lTDG
Omo+EqOZNmmxh1RPnSHSIJMsLaXmyRiL5Ec9q6YMST02Q7CqTu+My23+ZA1a9gDXYwkyeWG0MECV
eGBus5sjeVI6BCyKBvvRGKq7+9Alb59Ou7fsMg0R5oUxw7t4LXmSqSabFdgh5j7ABSrwvudVPm+0
GA6/OFZ4RNBqzClX6Xx27mE2waiT+pxvgQ0buAA9b8aYuC85ZziYvWRjYAGAHJ2hkUzvmT5oWmAs
BWjC756BijCYBCTB03JDsNcCKKqem1i/hzootzXcfx62qrqn33jHixtcEF/sKehNwEfYiTXKYzq+
0Xv9aIKlxVbv4rx9ws1RWM47azCaw0boHs12eW1siNl1S+PNbhFqd5Q98Iyg85w5+mPzOCq1Koli
AhiW9RK6ylFkEswF3YfFu0McwzOWBTQ0MAwX5sgpHJ+qs4Vb/qwPa5ljtxO/dPXw1o2yD0cOCkw/
zjxw9Mq4drYmRI6Vojq9KDXYC0n6Uorl5rrbE5b9zk0A7HqFL06m0U5rlaV12kVIK2BhrSOGtAoE
Tr0/1rVFoV5ax2F4VFESWcHEz/a3djCqLCQ2Qn+mP0AuEjyoRPR62Hezi766gAHEd2G6a42VrFy/
WdrkRTErAzl9jVDq1lFtm5kznqQAUKojrABweyPgpZoStK48Z7oSgfjntft/uaZOjClbVN8mqA/D
ZNHfxvnc27R6k3TcGJPeRDrbCjsg8DbOnXoyw7ades4rWtndrYOPUxZraUqXCUThg3QzIkOcCCgQ
LghAszqS2OfuNP4uA41jnPNrcNmyBvgq1RctBV+uy92fMwQ4KLellk5JbIqVoYzLateuuQ+aX4LY
/wR9M9QCtxD+nz5DCRsQLzJ+t9lUea3c8I+SSHqPHriBadz3/xCIGWxxAFkS1bm2GuDwUqhapFE9
3QGy5BYDGtO4Oh6L8pi6hqFxqoTdynUVotWqkEmxmXdSnNOuaDIieeawqnF+Ba7CMErKj32Y+mSt
DwZg9yviAR7kAZPXwX+OJLqGigvyKnnnp3DPn33MibBriflBkWJyRBW4eKpWTFKqol24FbZBWEHL
36ZbmQbVqC2BxHcEu5xGounuTy9thA5FqrloCcny7pQ5wbVb8WyZbFkM9kTttj8IkDipZWLAlnYY
SC8N6toRGaPu4h9h4KCckKG3MxlahIgUa8CoDyKoNqyMvt+gpecnxyCap/4HgA3o5ZwFhu5wirTd
EGco1SXpXNhML1e2Rv/eRj4TRAPPDdhEIAecKh6HASb4yrEKW+XEjJR68jDeg0guTkmhX0LdMaap
710Oachum+fJXLlUnd20gAAo4KTqu0//V6Nsn9SVJrAYdQMnto5qIHqsTEB/zFmJtFqZNIaqOyEt
V8YIBO1EhtLxB4M2JZDt0Dtvi6BxO33EngAO0mwzcYGX7QhRL8ZfFxXV6dHF2NADX3z2ipZVPMkl
weoMCVtpUyu4iM0n1WsFROthXYcDm5f4ufBU+Y+1p4NYa5ZCeeAzMXRf1jCgqOasvjkbc1OY+qF+
b9mbMyYJbSaaEUEce8HrSkvB3oGLRsAN9HHvyhIqtlaaD8o4PPUolZhFMyKFAOdIRefmp2wMU+KD
Rkp6Pg12tAF1nDWVs6ggj3CXAG8wdObJ2aqiD3zLL33nJbVJq5rbFqQdzF584PnWfKEzwZXLI/TM
fB2IzK0fFwh4jXmZ/eduPwU2/AoJtN3bkFThc0uHf2GZBgHKbCV9h4v4MsppuwtuXN+Y/fZWbDWe
yZ0RtB8q1ZIYwFR3Ox6Y1Rj3aMo1wTLm6K1n/4aM5UkbtiZEniqkBatcMy5FMIBSEn7s/DpSKWKf
E+pstDSX/MAJMx21oNxaL39B+IJJ4QNw4jYDV1skzOH21hvwp+ITuxNYUZJB1xal08JdWfoYJUuz
+s1J5sglt7B4+E2LxCTOtW8OeqkstOq7i7P6l59yYLMM0ifrgbDcl0TuSbH/2tHHiRmw/DUMNgHS
DNJ8LGVz1O6vqhUR5fuqpQtktCkDU00f2YFIRby9Qg6swLPrQ2aFDi3IxeHz12xIfbuLRVmhdPI5
sqRWmBnDhhNUTkFeE9XSZL2xvM1vTIruvTeXzK8X5ElbNX7i64i0JkEqTDO6ScAd+TaMyYARuxB5
Fl969llwLXTDLZIySFw8gsflSJ1QC6qpD76A0/WsgJzY4NW9A7X2DpmAW1L79Y24f33/PF96QlFq
+Hgw4/zOUu1XQv5aW6Io+oYy+dP81h+vDK/2TV3/sgH+ilwAL3Jr2pn9VlOxGwRpFXGB1nlF98L8
63tjecLH6ATrky+7thnLdCkx+/VHl0BtFV3KpF8a+TK4YE5F1dtsTWxLWFwvvjDPiglv6KdG/yxL
AbP81ArZL+3XnZ8/bfeK0hqN9Xa6Na59V8ZhmJti3NckXczKF7VJyB+9legwPPj448u+0+DWZB2e
gYRdcRgtD8sphXgq/Ot2CNsRWjaWgyhjXgYveqsX0J6Be27WsaZDmi1ErvLKRn+ZVN65G8DhYqoU
S8X9N5gxry0EI3zepSXft5lnyk8hiqkL66O3ZkRuddNOLptkWvtB6JsJCfTbMan6FzqH920rqmko
eyE6s+j5Bf8EoYBEXzEpgWPezst9uB49sGK2wU01hFTsTLewY+0JxBmR/UpcHoqj/dW3BFDaASEP
kEFT4IqtHGx4Cedj/fu+olq7lEPLzfbjqYZKe7PNt/7nB5PdnUB09WvjQwp6dvgNjJ2UF9kgpjJS
GsMIZfXpwoKcgyIitGq1+7P5z/+hOLXCdebApsOkotspTBYnJEQl7M9h55+ktNTs846Cj9AMu0r1
IZxDTrqkMTCqeLNwvAx5HIq56viCvtQdTq/2Nvvytq05L0zKW6paBzXYPK4jeSiE3rnDsXaCDyJG
ncooDLvt0imDAdSHRCbPxlq/8TTREjp7tRUmpY/vR+yr1VCIIIgIFj8J9fUU/3vCOneZQRMovCln
61yUegV4NRsxwpkgdR18UoP68t6olgJlnf7v0HyRvG8zO9agHnXcFhUCm6eaI47Ev73L0dxJ7myb
RmxlAzs6efj8xz9SzYbXXYCAYbjJAL7WXMpt/6LA5aQadFfTnjP4KO3HEFeM/nYjM5qRrghOALud
Enao0ZTmCS31O/W26kAjvl0nvNPnZrIWsARto6+jAgVtdHCe6UQLJvkQzrbgJB8JgaJoBCPPZStG
En/JmOzDGtIyQz+kxZWO2uVbl1S0/QsfS9bD/LlGGuEsyR7pK9GEf1EM67I/v9m9KVpgTCuiB3Fi
yJgGB9c/PkgBM8skG1wFmguTE/+IZLNgqx/deFebC+HbEDNmocPZpAsseTXujKQ3oSBJGuE7AdEY
sNtERuwHFugiuWefma1oIvvxwqzMnJC0cGF1aYFS2KTyzPvNVhvZEYlNM5xQAQpBE9sGziDMoJuu
YvCqH7BrqORab1pPsFSxGgPtO3zk7rNpngFBQgajR8M8q10efc7AbBW/kn3WuazMNvmbvvuggTxz
RAcX9YhhjHyCsSo5Ff0TI5R0pinkU8GcZVBorpwXLhocYCInSbQQO5mSk94UmSGGpnf/jhT5rvtu
d5bz3OY5RGsiW2YfB2duQm78jo7ss/B/HzOcEu8KwweYJFi3xLAajot0ss1IUwBQbSzKLvSLuE51
iRAXgoNknMLB46Mi9irywsVCIjZjqtaKJBW3d9Ls0X3WmfIPWQDSMEHrl/fhuplNo8jC8+zoQOk5
WKlScJm7SSzQLqKUF6BDpOIn+hjBtDP71oBK6PofX8YYjd97RhrvlWzh2wk3eGLcde681GJkSQLy
DY3VJ7kmbyN4s8D+Z+qo2vYvJ0azQaSgoxprpWX8THCZ3zEPBSljef6qiBPLEFcOusnK+OeqSBjJ
9W0bKaN6Wcrg0onhfBqKrQoF0L0cs5HiIDYDsSvD9qC40lk5QMJig2qCuXxGV7V2Ey+c19mBHOEi
X65Zh4H01CeiSF5Dru5ncag/CwKH0DiPz4mnWjQqrN4Qj4x/gX8rj8WbHLMbiRW0wm0PnHHzfMwE
NA8tsF6X9ekqTT4eHffECKFb+8RGseKi50f76VpQjYbYUJEHr4vAErry4Ux4mDV1ZLdrxJI3Q6YR
npaBVu/pFTACzEVauY45zJfJHUrgm2B6nNocLI07RQvyEfyR5qActEDeJmiyEB+zVi0H15gbqt4s
e1LO+aGVdJg0RwDt3kpZJVOdS/e1WwGQMTARriwpJgDsm4JUv324E6da7Lyr+Jtj9FH8awJl4Eon
z+JSIbGh8t5dKUIGjDHcOBIvVtp5PgzOkyTMeyTVwTm1IgY4Blwk9vLefjqy8JLwQtbkHhyR6dpl
9aCD3bwAd9GL4Xqj5f4ShO/BUkwBSdtSd7/V4Sxg6QeOwKPqKkT3x5o984/DSeHgkJkwH/C+tSSZ
KR0K9MA/9weWxAaqLg2SOXb8SV6850XJB0fwMv981ZkuLMa/Am4jac2KiUZOzXm6DVhzYbUeJI1Q
N3OrUyhSUiZ1pehlYSIlqlw0Tk3ddGHv5cWeMBH7KFMwpxAq3jW1WBqn1BgTbWw35lrqU9E+geS0
9HuuVQXD+XMa5oHcJffmxnLASE+Q/3au4wVf8O/CKISYSVqs55PZHtRO02eEXok08XA2mO4Nu2C6
NlkWeiFHtZlxzCgEgh4ZKb4qQndSqwB8hOcB/8zx+XkumctCGj6BwioZvE8sOI1+heSu5wYkHCQO
f/qQaEmAmgmLjQ2xRjv2uwGsBpEiWqekq06AabgOTxF76LAhH3tZ7x3THeWie3aSdbL2zgeziAs1
ANaixa8Hac5+9V6KCjqm0ELCRIxc6N9ZqBYBqPg0W27TMKo0ThensG+55vFnA+DEtPJnm7jVpxwW
2uyBG3DcxMGrRCst4JH1e4Gf/Jb3GgKQ7KvT46SLG5SLeIxvLYjpnlRwYOshPmwJ/pyO+7ssUUAo
FKVoZYy7o6dyVxsyoNqXQcjBNxBLyUzGvnG24jnvtZ2nq7Oc33Y3JH5NxD+lB4R7WpIX0GkRpqaC
jiQdWTU4Xg4/ha4wzGeGqwIvvr8WWUjgDqPazo9GNGvjrbE3GQeSro3Q0jLIiNezPDNB+EHV/zHA
RGDwVD0euj9XsVyj0B+yu8T/oWh0EbbaLmAekkRy6jNn45fmqdkICywp4Zu89DhqbTcry98fABW9
SJrKWVDpjSl8+mBPCVshDPO2ryG6ydpNA7EywbX8KYIfoNT2HFwZvs9CJqOOorkSdES8Xm1U5Rrm
jIy6xhgsjjZrp8+JS5e1oD/ms6lToROGbegAXkIs4GFB85aqBvF/MiLOed55GjHAgRGN1Tll4RIJ
D7/PEwWDmF/STt89A4qCYWrIKGLBXAxKD+04lW8XiIIqeoRYkFfrUpSXON53lmdHowcyGychbUjH
wMJOW3+m2Amg0IGDCeC0BuyZer0X1FhvDywdXidhkpNGOGhvPtDi8XjHiTyblKV2/O4oo9FKRvSJ
7u/rneOf4Jpqzrm3G7Rml5EFCF6X1x1E6RfNs/tk2P0wXnqG6t6NtA+yOi/9njs72Kipd+rKkQmq
t+g76IGpfXbAc08ka78bMaYMixFhlNgR2XlcNKGiX0cQoO+Dh+HQOak28GXny+Tn81IijeuV1FJZ
ZVCTihXpeIUhfPjS433AIG1AYFvwIXC4HQrDZu5Cph3MP1NjVGF+T1zu18myN5cxai+lthyEV+Tp
wD93YKEKqIRIywxAw1T2x+DcSDJHodKt8i9xYh6tWiEIOoFjGLVkHtOzLtOZA780O50/o4RIUSfY
oDvplm++w3FN7Cc+VOvRm03INJ8v6JbEeyxS9r3lfTduMSITzZ3S5I39/H9EzlZUfr0/JwQrWFbg
eJjFvjhZENGmUZrkrhVbXt+Fkxf4uBAJdSHbqacnJ+lDXZMXLowCt1QMCMkm/TzyTGLLXod+AM7C
vAQj4Qh/oXZpbZEMB9inzldPtoP9VkWRw44yAtlamPbIk4hEEfyX+dWeqDniMxk6PRQWwpOOkfKv
l7aj0a/7497i0qT6MHGjP0CxCm7MGEXYeS0jchvNbfIEQZx1Ejtjpnxc/BpAXQ8wSLaciPT3kVqH
84dhTCbiR6DHc5AjCjxHxxmnvdBe/FTF2IhFw2ft0wIgTbDuBCPquqc8jpShqCCGrG3glSa944zP
fHteuvV4CboHRJ0Q0PNC0hxUFrB4A7st7x3KgYD9wRH4RvdfXvyFXBNkghl1MFi7XscexW1k/gtJ
Dps9OkeIiaXVaoRp6Yu0p2ouAyf7TAtStiszN3naFN8Jjwv5+7406Q7c1PdzZtlIUcq7xVVQOewW
bCeVEIr0aeKd04ffhKuEeteB9oIcmw2fjQkJ4gV9As6bI+dRT83ED0Z+582YQv/yq/Soguqwc1Hf
OAyjEhWvnOzfy7tKINNl+WYw15Q15UK/ybqC1ReVq1SnQzzzcnziZSqXxovliElz4glZk4YeihwT
VMwDsdKa26NuiJJ1ECbfPzM9ZgRAimQMuM3wzwzvmacQvBZqSNbsnWHP0h43ZjSPoWcrt3kPKgJn
Jgtn64GYmIoMTQfjI+MRxJwZo+oXBz6iL+4YcC1phgey7Yd2MDyQfQQXSuGK3qSICQ8ny9jvBGOf
CuH1SSszeUYmuez6d8JISh0fMMkvd8kRA2TUjcbAfQT5dTPmXpBrkbwqaQW23S2d8VjJCehfM1qn
sxPSuSfdIQvJbubqcTRcTTfI1hSU31qpGgU+WZtt/UQ9KqR/OlBQeqzwcTJud7IczwOrBTDglVsq
1XoJ5/jgBj2ETaSkOWWkxK7XV85C2Ranzr9OIEXeR/vnjpYvMLRa2LTmHhA1jJhu2Zon4kFZCbJ/
fSRTmMgW+F17EIWaBIRokEc2VtYhzAg/KUKab7EPCAPBHLb4PGl/J2MUNd7LJvmmf4vEF2iip9c0
QphrvUXlOpoU6LuBslkskHB+6bO/8F+tk51GhRGGeLr2ctQWJRt3eaVtz1EqG2fXm5ToRP+6y0bW
HjejWW2fvCdtSHB/3OjhgDHSBWjoNT1e/biwGKai+E9C8jmHwYMCTIXBTCgasCyp4A1olfHkcbk0
6rgBW8RgVhGG7SeLLjgU+Q0EfKbfa/d/k4QWQdjQMO3War6i5X/ryHzHis/8zYhQ6SxpiGm1vMle
oYG4mVGBy9QWAPYWkPo2jfTN1+JxkvN2AYWA1m6XD6aOkjMH5YWmUzWu6l1iaPOgPZu62bK7qU6C
D2xHt7FoxNqFX2oCwLn+Swuwff9mAoA97Z6q5QszhrFy0oLDHPTFwTeA+mpJFFgJvhrh9gMkdcbS
ro+D+wv199U/fjjzfo39bh5dy8smuI180Qf4lBq7vMF8J+XSnb/QeFafyDcAtNRM82E5g1NnX+zP
AbhXRa//qDmY+VcvTjwo8JOz8kLqeYL7bhttM3UZLW0NoVBZ4UJdtPzPDnWiCGRt0lrlUDQqmtrU
oH2zn3AJ5ZH7WnByCw9MHURI+WNbuipgp9+9GlCfoPsAXUEW0dJrRBtEjOb6KGyHgtUaKvi9d3Aw
Yg7U6ZDHuisRtlnonB2lVQC6uxEXWFWgPQKCaAhECGA71jHfN6QTY10qCPCRsZXT5iJHcBugmZ7r
uFPhlj8pN7/ZXi5NkUITvM1mXuDmx6tnQFJGQHlY0a5M4qR2zpDqHB6vgmV3fRobrPRiU8MlfL+Q
Jdgjb0Yf5XohZ58p+XUCGB8LEPEQVwYHlt5aTeJ8rz1IZpmBk8bRlnIktn41lTBboErddqKprUHN
k4jaTvoSheloaU+FdSsOK0XFkZ2UFDoWb+f4lvdFgmr5Kq15dRqRb9tCsRVvFFtX/rC8/ZE88/mQ
To3tqzmx5vCVerJxvyEdD3CtyqS7/yF/9zRCFOJRI5irlHq+VenQsW9bJj6EhHJ3zkFGY1JKWb0R
J2g9hxhwh15hfZXOOeaeLFc7oauu3KGxSqXgf3ydcHdWZpr+JOg0Gf1RcXIfj0LuR4xWGQc2Ujcl
XPwsLWzgFO17BvrC0oYr7YSQJllwFSiZNXrG8ucq6FpqH5ealHcUXZZQfoYFok+mAZl2IcVOMi/7
kinLhZqd32tOhXMZ3SnzF9SENaGmOD9UWUAZlpLfghKsNbKw7BBhO6m/dZHRZmdFj8v3n3U8ntzx
LNbiixmJ8mMMYCgZQVm7Ee8sP+y5Kp8HoDcxDHfSd3+e3m5RUT76UJqKVv3oHaOptch9FMxmccOY
CbqsQruDUqJQV5FEm5EZ2hcJ6jIH5Zt6LJanLoltba2KhkenwoqU/gvsPotH3/Gg/xrqHpZphznH
/Maa0VYaxpZgghA237G6vdGuuEyiaaYe5fWk86E5yAEuVlXxNgbPysFXdTS0sDrGGK71vlm0/mnQ
DgSJHTnvCy/2pbEz/3ncFNc8e3R4rGzUxnTGPCq3fa7xvxLfaPXHCe7ncDB1FXKIMRLQoKPmsk7b
1hk68jf60DtP3KGefzqQyOwN1fmEc0GGMerKXGHwTjnZ4AxrR1zN26P4d8VwqAPJzxC7UzC6ug6w
tqKBCOajO9pjFoo64ZN4Pts6HaT441uopRiflgzl6n6ExaYutPICtcFmyTWoDYRaSn8GOaPOXhaP
yJ3OAQ5hqbN6nnnhlzIWfaUrpoj4Jk1i73j4YnswIVU6k6XLNNGJkbmrUkW+4oY5uzv+sSr5umHO
H73xm3Vs2h5sXZWCGnA7U+/7yfz/x9TvTJVE0xi6IiNtV4uamNQOS1fDyn+AbRS3OqlY8GribIBY
VvD2NcX/ZOsrlIQgotSRseeoHaFdPiRRtI9/HAxGHel6F9jbnqPBpXanrXP34Y9huFa87zh9zRRj
oAUMZnfISj9WCbhFM6i+7vIsRysSLRocOUaJFkbUW/WHd52uKF8NhbrAGn4piUtaPpqomqmogBPm
wnW8/BqK2LR2pM0ADC2vUKnDvYMMBTLr9eVRlAdhmirbbD9fu7iQWTsOlM8iSEX+plqS+0efQ7FT
hscnrcwk6AhTD8MQSw1ouGAQQoIXgwb4DKOJT5Kygi/4m/idRfEi29pLIIwYJro/jffhRLevOWBt
uTsOWZTwSobJD1Irc3zTOxi9uWnuAszKlSKYvVqPqN3BfowGy9c/mfEaU4kYoVMCoMpE17yvYU64
bw5Q9sfXbM09hMzmeHKtK0hfXa0YHSnP9HeDwhOKA9ukROKr9BIQe0sfuxArOzEUBm5y8po71MyO
44p/NmQrWWlooO6rZAyej0NLEjuzuLGBw1/ib1hE4dh/e4JRwfqgvY8kAR5nAtcZFBXC2eR1EzpD
yaLIEFcoVPBle8mpv7bQs2BzfVrxyjl8L0H039L0q7O3gzGmswumubXC2bXTihYe4eUScwTFZ8MN
wE57CmDmCqitzjTetF0Qzfdxz5t8UNjiqIxaq0xgrpPESwdk9ZoIjKEd21UiuI80oooTijlRWaXq
VgXMuWmAIrujBAGNoe0Y8HyX1IYtz0eV8vD6ntzBzgEKxBE5nGOcWUuXgBIxsM/nOFaHMzw0DcsP
oKOeFgwk0eRucM8F5hlk1S30yn5ncTf8PH/YD7iL59DhQvZ4i3bI4WV8WTwNRPvAOSpDdLfxagJ8
Tv2RmL3lwNu4FtEm2hLHPlOFGxQc/cr/OFxPa5kffdvizRMeQRw4+TA4c5fK4qmr0mO9qjhL/PBF
KFO5/yRAV6wdSmxvzfbVhWxb0zlPVZo4QMM4ScYkSszIUvGk7BHWNnBFi3NJG1SLGzPna1adRP4i
JNiHHpVTklsdPBe1BkJnNfiRe92Y41wz0DACTKU+mcpIav3COGhEFBvN+kRXTJyLbONzmTXQrJiT
z0zdwNcG7GJ+q2vYsrA/QYUm4cJJqhuZYK+MKDDBBQnMEjXsTIj+O4KC4eGZu6MJXlQ6G3+sIuEW
PIlAIBvCErcLpyPkyiE2ods492EB6v+xl8GRIslDNiQw6QDs5onTQO8+VixYJdL9IbT4r6+N+IMP
hN9PBPO9Btr8VJjhn2vXExRura1JcZPN+Mg1W7zBm4kKANKeovSK2LUeeFlW20ZQ7YXdJiQYXU2J
AXfq8kAfnsD6L8vFlIBbOnpSV4B/w9qldxlK5Kr8sAnUguh4magJM5oZVfrUzvseWM5LTi7DPcII
HrE4hLMNE+AyCfJuPPlhlnfJLDq3HaSa4aFNLj8+JmrvYJWcQODdP0HqFgkUXhofnxumNuqi0Y1W
Pvz2nMejGUx1+FLVO4YMEo8NQmKhNv8Urca+K2/atZwjT5sJhJuj+nlYfBya1tztuNIKgRSdTsGG
IhxcKaDhVehHz+sISedohcdC6g2rois2uZWaK5zt+VT/gUWIkGJ1fgijFDYNdyXQXdFj/M184ye6
qhMd5wKAVIBEnY3yPBeLyCjMjg0LugW53lwM83GlfJ9t+gM/oDTnJ3+pRBZ+PgfJGuDgBG4SiDir
R8UQ8o2r7lAFc9RFlqyxSPF/wtvJjiRoOM4/ACDfl9fuoH4JQPU9VrmfupvsA8ecm4sbS5VP88wO
AeiAjI/fJQok5KgvSvk/6ZiAgI9pt48+FF0xUKDhsW2p/oVzg1bF4ZHjqbqk0VSXE7FSHqdctz76
x6SeainqD50zLZkf3CKlPfEroXNu1AMHqOAyM7Nh6zcXT5p+hA5uJmQVx5lgnQqBSNy932hlgyB/
7LV2Du9gxuG7l8tQrtYgOPHcoIWghxHnENZSqNBZT7QesaVKcku5DIUSDDk8dor/gxOCzYa85/ep
txg63ld19e6rpGiaYK5ifDFDn1Zh4z/JKhSO4aXEfgSfBjNePsSxZtfJAosXt5H8c+9CFqAa5ADs
wtgh5/0oF20is/DF4mzkNiNJVB0eI07hYHFZmpc4Rkh3XfoQfkbPRIr5RuBFt6ONOynU6c5pN4iC
wmTw73ihGdh67Qp0tiK2N20vwO7SmY3I8z5SupRCM7tirmYvOB5tHgXizbwupTPZUebUxyfFSyYQ
lYEzm84Z8zT/L1UbIzUNBMdPyDbvMDEo6vFmLHj3HtsxOR2deoqG7ZLDIEn1pdOsSnDZcuUEsT4C
PP8PYGpuQF0y+06ubLmckc5Ke3yCua1d3nJAFPLezcQ2yrVecmw68hyMjJ+L7NzwcAwfZDmFL5rc
/tUQepkmIGWVLlHMcuXdG37GyzSFk/fHLBSx/WJsuyTGFYXe90aikpGDbMDk8aVSBLMXLtmeyY1u
E/x2gHizVZ8TzPiocbyx+3vGJiCU2YQ1jjAfdjOVxq4LArfBzpvOhEXoWXQddc00MEz9HclnVdTc
liSXK6DyWeYxFaIqMMDn7n5dMm7ALTZDFsmeEr/kIq0Qis863tHxLxPCgwKqOar3bgXczVZQtAQX
LDiQntfUejXVg8UUYBjNXGZxUnGjroiRG1hqMEPw7+Br1XN/5I+XuAaTazO55ZM1hSPVmKfdWz2a
nGL0SrLcVIBaY3Wsrsek+tEvDdYXXSQkhDknpdjXh/AM2U+mY7G77xgJV51CY0lcNnUCkrFrTWQg
KNRSYNA6W8c2UgiSRaYA54q2tMe1mquDB6E3Y33YaiIkt82fRUk5pj6dYVQI2L4pPkW9xv11vExn
Vy50knEK+0lQ/kBYXqxvoED9XStHoFOegPaNBLLr4Jqf2ANHnESl8UnJ+T+/Nmyt/OET5pGRfxG8
S/KXK74LlvABdnMs7Hp5MxD3qB+OekbfR7VhkpJFpT3vPwtk1jHLYVh6ZqD/NkdinQ/teRVaW4aN
Ax2vG8auS5NNwUcu9pzCWMfjJZaltysIE3YVYpbdi0Tdo+VE/xrEKgzoj3xxLHUOuEjkdN/P2571
I4QacfuzdL7+XqFry2cpMvLajGpcKaTNGoJ+o+quw4F8c7dlnNdQPqZ15HtLITmh4WYoZqe81uaK
RLuzck3jsWFHv2pG09MXh4pb0uHynrhUmzx35xEGBFP36o5Z6bsOF0UF0k3MU7cKcgzD25K4gGr7
Fwg0ym9Te4O1MgAkeUPFpLImgU6WhwQlAd8VyayylH/jNiw0LUIMQAXHzcqnyuaAFImUzTdVH/ey
p3JghvtVNE6aytvtfvPvf5ulb1HV/gA0d6DXW9kqacXoAD925JybqRR1Wl7AHmA4hup35epJ802p
KNJJGfwcnmaAGffWztDZWwsk2jlvX/vrMFWP7WvH4A0UXx3vOAVLqbP154a6QRPFoGBSX2u8nExv
Q7OSOwunnsa94IvN3TK3PPBsmSyNPlu/a+BWSLkAbUhLMUQPXqNlLg/tY2tZK51T8oIpCjDt+ORv
N2iYVL0Ng7+4XnkwVlWW3SrhGYChysU1LvAcUmvkqzspP43vsNSgpLx5UoTWrR2trpUB5qB/tRuC
7x97A59lTAuFCpFJepLJPpzHD+XLaQ+dt4HqzqdtsdcXfbL3m0V47WHob4op8bLrduQDl+K3cb5h
o8+1hUWCKZ1ZfoKC+llI5qmMGqHgfTuit/v8pz8ewMhhJCQOt6+t8hh+0BzJdzlOStyyA2lEFluE
IH9EFkY4bw0T/J82l/mlKhzyOcaBn9bDgUfG0Pd2zihZ1z5f4JTtNRgY747TylKmf/TqmkcJifjb
LqarwJBxaXRu7lLhOzhSbR9TSvE+lXp7uxsQ6YFpE5GGQSp7Yq+HZ9MjKHrHsC4ZT0WXGf2EzaYT
kAJgKjVq0CTeMYeW+p+uJayZKb45Clmcdoxbd+Gzsmz+25nXzA/5iyhjwpN4yQTR+T4yIcG/hot0
g8rfOa0iF8J4u96BvQBw7hW6qp8RERdBSFvBHPWDRJr2O70sA2DrYZ9f051lRhCrwXrTBbBktZZV
gJRQjZK3djN//lr8sRx4CjqGcWn/PF6FQ+TS+F+VwsMxVOf6tjwTQvwQ1StCymf7QcthJnBtxLCo
5pXU572pBo44XQoJvwjXT9aosp1JhyrrbCBIp7N4YFyOYfOQ4q2DlzraE9yiqRdqAPTlaY0O1Ht/
mT+j02Zpe455NZBywc8g64aUWTzRxYBs3SF0ftOl17mEZqJSXiYN2ymlWSu7dB93YPWP+SMrn45v
yAy/7cDRgYZdTPK/1f0nnOBO5jv7mtq0Tz8sBCd6FXJozdgMTHczNKzZrTGTZ33cVznvPXEIpfQh
5NL0kd9P2c0KZAFZGacu9NAC+zTAufBIkDsaxosy7vK0Bw3JncYUdFU4PA1GwGFqkaANUgklZtq9
5CxwomidEL7v8DIu02vzYY1QfKYerx5zhZzuAUWu5BO7RJlOpFVJK906V1uRpqDmn6Zvuw86Q/y3
epczzbXn1ANHyeCttFFohfEomkhvg06Wk9M8GzUjd4puAWhzOtcmSTkDfjQwdNRcHtbLHIgr0X71
EmhkpSfhZdemFdaKuFZouzptprIpNrsVEWBEJizJVWAP6K/p1ZmB40+hgihugZwm+1Dvg4wI0Nue
YrdUPuvLd//upXE1OXdZ5QeMkdE4kkBMoRx61Skq4P/HeIbhobJQ1CRJSqky/lWyFdGXUOylPtUN
WmgxnILGS6aN7eDQZEoy2aJfxJvm8Dd6SHEoSX3Zdv7DtfJkhud4bBxLjl3VVvGC6NhhIqD/mv92
medmUMnw6Uzaxerq9DcKuCpb6Wg/hOn54MQX2CyVJRffWjoXwJ2eKTHgVL9wxXlj/rEP7np2zU/T
/Y/KmIdzZEhiPUvkZa25iNKyhoKILEJ8Gl2IIRx/pWdO6c9a1eQSvQwnue463u+LixSNH7sVVcHO
OvQoYpKuUu2YxPNTzhEEDbBz8b8Okt01j/hm5vuc3ADlaNIS+guHd5mTBjzY9wvOZCAMZBN5ASlm
WIAfQI7wZjQ0frm334oQ0wxA5V6CfVUUTUvTSl3Mop/qJ6H6jr9pmye0e8CVCagUUI2rwGpT+zgU
FjUy8wIq18/c8IkuxNwsAKfjYd10ymFzICGzbPdyH0lh1akEd/VMgPEHGilty9kOjH+8Tc93puoh
ZfzTGaQyd9xR4ubsjYdgHeWRcXA0QQVXr6RN+OgywA3t8eESYPOSGMxpWpgxj7JWBa0lHMZwQFjn
DPfJs79dCdSGC4D7vukPDc/uNXuGcVg2q0Tg3kZkcfZmyLMoZ77TRcTrK2b9apb7AiaKD5a9I3EH
r53baherqFhnkKhEW7t3lQQ6QXT6bWKrY6giRcn42Auq8VchKmdnICuclaOO8hTW8Q0lbsfw5a2t
U4ZDaepJt0jHCaTN+U6pMB8jnXPdZn7zJZ1KWKm8xi6fmzV4YDBZSkgbmDf1r14mpOys/gz4ft/n
BWYSSITDzrYHpkIua/1vZjC2iNuLJuaR2dXb+i5moPkN8JWQ0a9NiLkqCPuJCSDUuTBQwgH9QgOm
FGqQM++sjhS8JCyWsWJ//JZWMkaJ0NRgwJnVJSxoTdMrnoTTZjIRVEce/Q39eNTwMA9xts+n66nn
14MvEksQbXaY37tyaANte3snMn+NQdaWGBv3ZEg3JIUgqHyjx3vl7vjFvLGqw2v7finSIwx+y8eB
vOjArOxesPdAvXHrCLfFc5OBlqlm5Q86yHKyGvjK8sndzxkmvUtSsgNurGxYV8MuR17e3f9LGio4
zKjU/RGyC/qTCd8GewY1qpOid+ta5FpFSAXnytapTl4sXRCxjjghPlmQygxCUgQlCLOitdDD/Yyd
5wZrX59oyGckov9fH5xiYCbq6ykbg1YZ0Sk8vMXEXo6FUCkmyvtUCK2YJr0LcLoj7VjqFTakoIJo
ChugUf6pToh85p7Jh5xPZImqmTsvXWoDhGWJmtbrwyDHSQsdg/pMsjiLdLxpkn4170XsRrfnhCQ5
TqjXZgxLCW+uZ7Yb1tcdPSjlUULXoApEChu+/VKBqw5f+zZxnVehhFW0FexJxj/K4lNxz+W6Rxk1
jy7TqAxgNECGUKejew3ao3EFu5dQlNptDivpBJCxLJQ3UgUrCmsZ47/zVNX1j0cfyuy7VeWrhzpJ
LhKiU8ZSgO+qDeS1smpkv/efXQqXnx0ZHVbErjfcmy43hxF1Gq437vSQyj+6k8MR7bOwtGco4atA
749i4iwpxpwbzow4dSJdvvAPOG5CQYEPj+CE8hJmRdgpG+aD7YM2wO1rmwWxyLOlEiDCb0ZX6Bnf
mM0LmM4rwFBj09AYlX6Xmv5p0t2pB7CGlinmOibdEgWkBj8FZbZNGBUdn89uVA2ysBoqPMRq1HcG
4ceT+O1V4kh7NBKw5L3KsfWLU9qdODCL+aX5oBFYBdL5iqxu0126L0eCnETsido5GtkmPSbxiL/L
T8rnL0u3X3+2jSJ0zMw1Gq3dOGp6hLORWtuT0qPL8vP8SMyCIZ14dJre4y9IFk1cVzH2srKASzoS
OYZFsNaKiBz8JNx0+Shlq4Hr+LHblfpiKKdrc4yqqbuQrCsQPz9YzHnLjikPLpRx5S9wluPO4fzM
gzVrceukwqUZa06BF7iKvXfX6YfNKX8wq455WEbSmypWLe9Dy2XdOWjFEQjWyxNIOAEkJm+Xyu1L
82xSgCXiOfl5u/oG2zEI22MZHFMoLP52DEASOciZ9wPeYY9t5WCQ0C80h3RCxSHnlNl5BiSy18+J
ePAjBfzUd5snZXLWN53lVgH5Zce9YT9SqwajjfbvWjS9COxl0FvO9dr+LoB3WHJk3emEq9Vg6mKR
lPxEg8qgTRP9Z4fA+7/w5EfiEB/I2F2cWBZ7ggh53e+Nt1QB3axNtihoj7N07FEI8z4uTjzqbl7w
+rgjwgZKXRZv6KHTRzw2X18V8gIg5waK6HWYq6LMh6fGCkZgtzpzWFtmZJ/ZbT0XlfUm5fxuZU7H
RnVYzGObguYezT9l7XZOjkF3IiYUVn7X/9xv1CBZdRVdZ4AVotArEFXXNs7MdOw3EnkkWuMnVEUB
OCWtTiEJTeA1t5gijPVdcDGfx9yEw0xX6d5odqb7pZyVWZ6wm2E9MSvXuSLZVTzY6PTp9saZnvn7
wvNgmRgt3bV7Vc8ag/N/ii2RBz6kNE79c37/eI6IwNan+5KPDBXYiBdddSzkjQ3Ug0ianMbKLcdp
0eoQZSJQZhZ10eKDSaji6bX3PElb8Pq5BrnFLGP5x+sNrjtFHMJB8gjIO4Th8keT6cwY46ow444f
91I0zntzBYB47/VgV+uIFd9jmtJcT8o0dC/N9ZoGkH/2Jup72D0dDEV3OzrX64GF+pZqQo5+z02w
mMabSBUkLo9qZc4+AJ/X9lKHhgFsrQBAB0NWZQyOr/eo3VlmnKXLzxnt4ry047Jpdl7zr2nuCFng
ONHMZvHCCWud7vphH4BS5V7Ux4ne0KjbZOfq7EHOXghVsq6rJnFzZJ+1ALsqyAeF9Dt/hFDdRg4q
hLkQRBhdedXg+RB0fG6aTeUVFppXNddDTJXUORURZ80x6oMJRt1SJ/HdHVdJmXOP3N1wNDt4lfdG
HZihwirxCTpgqOrc7Tfb3u8DoWBlBK5UzadqQQhjGA4p+Gh8QKsqUViUniK7SH/nCjgHwtDVMqMl
z3PGIagmIiKybwd07VQ2k6KknYKhpNtCLbl+vNImpN466OFr8NucuL2kYFLPedBdXHQm50FVr0St
SKGWL+GbGSf+OiRC8mp3T1wpKGMMkaf1KX7eKui7wUMYAdq+T7yyf5xCbPn6sN8SDSIJJ7f7svmv
Xfbyozh/B/fAnPQlZ4gkvZA5hiJdfL6cyY6X+yzuXXfxw1UM7sUX5I4OUcTnG4+EHkUGEcaJza/i
0yV4JKSJtsPwiaNhi/8yTc5ZK3qXI9v70UL1Y67Iva7NYE6n1FlqjzsNn3zMeQBVh8JR9xYEKT7C
3NEmse1OanOV9H7lH593f3nujSGulgAfWAJPzuytHqeBWCMJHQvPM85ZTKzjbsAncehSnQIyKHBm
hWJNXTIwVlIDEqas4PZ/hyHfyT3ewKdoPklkpieAQQKUGDUivEjUN5Q0QI9ImoQ99+8Y0QXAO0G7
GJWOPNI3CfxsKWHEGTgsLLs6Nvq+B7mXVmXHV2k1SUvdZHJudzmWa8GlDJ2b4mERORcpAQJJLCZI
qP27xnZQZ9Jd0jO7PcQBWHOmCYmHPhP+c3V8xFispKvwF2syrkWTJ5eOKwLGHQRW6+l6XHSrz4J0
7MRsSw7q4fkrXNR3U7x5s53NWSjIocMX+lL3enhD3cT6EzOR6a1R251u3i9jakqfLK7FkwBuMpmg
huW4/lHktbF+KHM55GZG5K65gXcMTyd+54OsBn8LXh+lfUUUSPFf/JpyJppawbWCvGACVDRYagiu
EzdP9oqRgnhAfhTs8Gly/BHmfuC7qCqF7Qk2WHy8rb31yFZDTKrhQW8HFYhsIkBfLfv3G0bgia8C
eFcjjfM/3pVY5o5TSb4arjfE0lpBCIHx/Y5NyTdwfPTcqimhDdw0Jw5xyzxdwabcP8Mc7Vh914PS
lM/cA6BLnDahK9ciYjtRhl7As7vj/sely/efiKBq46rJnTor75+gWkwxn1GrqrsFoEmlMjDZFuxS
N1BACTYoFlDacMh4bZxcxeJov/96KPC9KEyqRzT5GFcPu6hTwcf+Ks6F84xMQ3rWCWwWt5wpfiJU
ZMiyX2DHRGAQy5DZF1lny/z9jSgC2NK7kvKHKWwgAAAnIgGakEq029R0AT5AhCDTyFRp9kHEUIyI
sxdYZ4OYgkNGlMBBkWEzeqRGntmwOoimx8njmsCnC12WziN056b7R3gRfE8tf0nhc3PUaEcy9bP3
xCOr8HmVmqjdUKOvhyhAHl8lwQe2elFRTbCGJOotDpsZ6sFkAH/S4zedZE+PJtQ57Psfw7jN5Xnv
a7z2W18a94bzSqpdcCB21fg95OeVu/dBjSlcrTW6vAy9Vx9haKXGSOuZUEGC75hzcCtTSwUDptZt
DMwIdkJccpkYLloLhiM3V6Yjgh2qdxDUPR1sLE8nSk0aLHP49+Q6UdWa/iD+DoABAqf51peL+GZ/
hkHgxbupnOFsFSE/Ag65E6DptKFG3GtGH2XP+mnL0NsxvT9sJIWzSdx50LUVwd1LpIW8NGLw9CVe
QBLtz2Fj4UHkfUn7LSBhxYyah/3s3EdAFcxmezlL1/3Mn0XgJhLwbsnKN+Wiber8fZi/ewo+E2PD
Q6vele3zwQpkIjYwpV5i9x1GuWKTHMDpUWilOdyTSEMeSc4mR20vyOryEec2S5XDKaV5MTiWvc1m
UmjgK/fYCuftLyKnGzSKM4yKwRlH5FpI+NM9EhJauJZM6Pbx9xib5Kb0s1S50rlz6Pl4UrbBGOjN
7DL97G0lMwNoU39mFc/AmYv23OTc8aJ65HarcoOsYd1lE5QKegnYu2Nooa0MFossWItgSt/HMNVw
lmRuBKzRJvxbdKdrX5nUFdISkWTXcXPc4p3S8IKHKs88hRmDGeTvLKqQ5ZkfAoEi5mpEUbin6pOl
51ufUsM2km0GhgJgcBWLFkauQ8di22QTe8NiVW1iKD0IKVHf+36r2vR1GQcrad9c1fy2MdEkQVt3
OTG/UUPxsgFJx3APgR4D2TlwARg3kXXJtuEEikKwyE8xMXAeB/0f24JpYegS1cyz+d7SXnRff6fD
5XxL7PDIscRVb+BMQgBQ9NxQs5OOEa//TqkGZ9xmK/WO6B0S1/xtxeV6GDDiu9q3zMIPdP4OSBlT
AkxRuNoNcstxQy6EiL2XrQH/FUk5dBncxZ1xlZTlHuAkrbDJ33wyQayeByJsyVDfEIRA3DsZP95x
+rvFwMcBklPR70WTnFn3BOSAP4ExoE7zimsePKnTEUHeY7vr8iEcPnWC3HVnqkpojI+fdahMCXhi
TM6v19FHaFzHfXwryj5DVlwbSMaNPYkMZgARVU95+KsdmIKFUjug3t1AdmkQOUOS3VCVRUaBNY9e
2GwWp0qEy9CUf/5XNkzupD1QC9UA4pfaXllaGsbdil57pW/aATQ5ROX1iJI+CGQlrX1D5PCGTEUP
Qk/pctCO+rPt1eOUladyxRjNaZG5L4MgJ40ZLW8KpcLAyz1ctjNR/xfzc/YDEBpSu8oq6OU5dbVo
ZYZKo4F3NW4mZNBNxv2sAXw6FvCC4pbb3GBC2dq+CjvbOXhYV962tqxdxZjEVvd2CgHD0PqTU9fV
U/IZdAOoKNGc0VuErMC9ABX8sPeAAjlVHj3FJOPIjShDOKIAtRXT+JX0D5arYS2yDNrfgmqsiz1S
WlG8AWNqxxqUOektLZQeegasWE65ezwZVNSv3AGUL52/4jreOdfd7BbfzeKm18RrGmk2mBpT4va5
cyDPM5t/OnB2D67LKhqWvrXbSzcNUKHGmMH6l8d8hIwYqQe9H65u7MkwZ5qjEVeZdBtp5HnavTOg
tEwpK4Tp5sElJoLXDtIxb/kRYTIsng7zZApYMX93DqGLuyrfnxE7/Ts2KtUb+i02p+4Y3j0rIQms
YgyYvwNxOJsmUL8Tsi9I8Y+Zsko5V1PKetQROOp8rZQbtr7tFoCMIYKqi/9kpSQ0pwalWlV+V8rQ
ktZOKJA5tynR/4x9x6Sb3ZjhJkjjiZccJQfjCbPzYJ0kWmkOdAUHCr5yi73uBan5/AXnfOWSYeVF
Bl9dQXnLIE1PKwQBHzQ8pQRHbwdYGkeUWliL/50/IBcr7LbIQblie9cH5ADWhP26R2DIDiMg7LGh
mhjqgI0e1TDObDbdeQfYy3S+uLyJ2OTGYhfTc1hmuYnP+g+5yjHNG2k943gMtbknW9kb0u1rbdnT
1I2vq2n9uAwLSWsFbmHaee9OLwpVLLigYDZ95W5eZWhuUolGNrLqZxARPHTb9Dh6JbzEumQVHzVb
FnkB4s6sW38hYj5DjLp7ri/Y4ENGHMHvxOtHky8ZNyz/Za+RBG6VUuSvbUuOHpj3SoWxE1lDIsfM
b3K8ju959YHdlxT5A/Ct2UISjEdXE0HWy0HVnDE/uy+p4tUbeemJQHmOOUtng9bBrnOAX9gCe7wX
Pa15dVy09cjF+ZmGKuEoZrCxbS2In1EeuSmrtF6c3zGHUoUlP9rQvZHmsZSxtXwiTHbGmkkijCkK
G1ocrrQqRNijZ3FsRGfkmo8Yf0CHyWzbVgSWwPdn4wYapM6ggv9TU5t6SlNLQ6kvFyDN0vqqZ/XT
S5DaHFFnXOT0Lh2YGBxc3CUBk/F1h+2Uvmd8NvHaMn0WXoN7LfoMc9+a514+Imv4Amko/754q+wz
Jvoq7jfB3PiGtZBjEiSiSfA5l0sO8sK4uYvdshHN2dGaTSH35EoVA3/6UJSJzwwbWcJPIdH8ZR7V
A1iJGGYB0TATDuhtiea5SJL0g6SauDLKg4XNCEhEivTvDrRDMHsPv5IeYAjG4/7ZvPs2BvDQUI5s
6qx7vJcHwZQshguPzCFK1IpOW+6RZLSg7VrN4AEbFEr0YU+XHIs0uRTFZvkchWUGo3gRvVnbOAFX
vDHUXVPttIsEmiGotsHidVd7V7aqXN53VnuxuLsruqmTqlpJrzERskI5LQtl5sbQ+ZSIFWXzae7h
f4Un/b5z5USz1c2uulCMKquEwrRTIZhT3EKD4ftGHpi8YxiWXRSxz9r5mkEqUJ8y8itBX5PmNZfY
b5o0EwHcULZdc6KJU/sdndBlJPldOnjOqYE4FJfNl4e1SwAWGeXmKn2pvSRAVAfW/coUok1n1UAU
y6SO0EpUJQrrPkxms3u38aCZ50Ii7UOTt5GfQAjn2Y/icoYkvew560U2oa0c/0VJilGMqDNB79vN
TBNJsyPfkdcC1vIAaSZibhBZOKRtvW7CTlVpd5fiXPEYKExufUWIBIWqfSihKOVdpbBltXh2BWdG
zGKHmqmhOpi9v4VSEd2v+ppDvBJ1CHu839tn1jMtm75wfT3xECJrsCGfGgfUakvxBkiSU/Q1M4Tk
IZdOHaOjBk8IAOXlzwhawZDVjQlAmDXxpLZTzTm/unEUJDGD0xSuzC9r4xMTDwR7bUm66J3Lt/5A
XPlMpJcDZTnO09wq9e2NQFvOwWRzsIxr/8gOsJ8WM+Rs8Cp+FO1Gb+nXrLZUU3iKTg9KWH86n+Gz
ZNmWM7/MRslpTwd0g6adqlU/VfZy07UYgKO6BPg/v/bOgDSsYwh33P0JszEWHmofgtdXOmxXLLyv
loNt0Zhm70h5nyh/ueSERZ8dAxcAY7qIGj0Lv29MpEm4v/sR7SHlJXHwk39vON+OfC5D5wtMWpTh
fZPQfsDWkVWuAjRoqFBtsdzne+UrLc3J2Jlb6dmHIHMHd1VusYq5W5o3+TaxShA2cQ28Fzblbea5
dd2490piXxgiLAiKZW/NxGrz7KHi56R/t612oz+xY5Bm2ySNxFvZrmKvuPdnCWoxILZgdSfqYzFN
U1ZiZJuBpCGwd+2bPyz1UxNROWOAPaZ7CjVESqzhb/LoXXrNXjtgRa/NDOt+krcWI8V2P9jEB67y
h6ka0Ku0fFn8GTnu3LNZtcPscXjMt6M9FYhsNxu2tKeHAyiqUTYYhi86IQQwDk0F/Bll5PNRj4AO
rrVWTKLA0VQtOMpwsCKst89lr5TY9+a+OaeOxJNI7MM+HrCJipfQV21IDWpOQ2rhMrm8zFHCKLWx
170zhMKN6d84iaFO2SZSK4c3fEHsEj5g7okDIribNDhisa6jlrcLOpbDfBOTbYgHDkkBkZpp13Tw
PtZ5u6Xw8qlPMcD1MpEOT6lWYG5gPQ0+G950yM/QFAvjpJIFH3Pd8lPlF5o4rD5MHwBvlE6OAEki
bdXY/3qnqlkkupiJ2UGd9huOGO2eypXmgq1JB/x5B/CANcMS5TjDoh4R3YK9m2Gpp/7rnp/1DNVr
VsDy+4J/6bh3CM1ceJxrvYASL8zcOAWspufYgZE0lACE6+yCGRrPaYW7ThM8PiFOar03Zj7vdzJK
WApNTHUNh1R7lUpTIKmA48a1wyLN9bp7VvkphZlf1hT6SZeGc5wQt0HjKED6uGyc9+xCC9/oT7O+
NGAADME0hCv+HrBrOOTFH6uj4qWJlO6GQYSAZY8ZDit1bF+rqeLj/ApkmbsnP0zMEZpfx6GcBj/W
HTuQVlhrqEf4MxZcK9vV06GewWNKMpBeagutYKw3XJuNVLUBSEkVZdkE9cYTZ4+nDTJtbrovPp5e
cYjUxT/YytT6h4agJKf+5mNarjIKSiGVUXkR2T/8TJnndbbpVkbW+6zpPEexTDlpNHLzvHLQgwyQ
XNgBP2o1oRIVgpPRTN2xnhMwI3YMwjlGAsYzcirD+K8S5uUPx7rLDi1g75ioYmeZk6d2qu0IE+ue
cFv5XnS9OdEfG+59Dj0FViIPUM3qm+U2Vn2RD+c6ASOdnhxwOVa3yXSVVPahWKuc0k0jtS1lrQ8W
IpowSQhnu9EZJA0KLq7dga9X8mnX37zeM3RcTjvqlJYJKuSTjYxICN8oS7kyKYSovHiF3XG9VJ9O
YNTmhEVtXoeP0j65HmG0fi8waDaHgfvc7gYnkDD+z/pFtmjjW3YzjPbTYZVvQEaa6hWU2eqQIusW
ohXGH9H9cIw8VXD4wCMGrndz5Agagn3jGIr70VS+pnSqOSmWxiPWj3l6G6iTkTOZ5Ix72fvjXxdD
kTYvvESDMZYlgaAfYdfVe49O9bmjQ5qUZ/uEiavFUx49qoOITRvt2ew7PLbzLIG+MTRyRX5NktGi
45uPYuYB+wUc5yXCEA+fCWeIfRkUwFETIqc9VR8F9e81cEbF+yGEPpMBZTzXTU5MPtble5U1Z4St
G3836h8D+SGzrolThoH7v3nusYseolgZcJctB5etb6Xgm551h91SaoD1baq91+LvClCKf4b4jOg9
6TJkm6SjLwQtliKhmF1fYJBtvkrEzVuRNSlcRni+FhXJVbdxAUeY9lV6cATedd3z7ZkUmHwec08K
ntih7ynMQJvsCk8MMdBwB0AR42+KGW/JF3HTjC6tPG+3BAROLjBrbqFfEThnNr7QC/YcCh5ZA0df
m26Qy5Hy/saKfb2sLT1pMJ49ZEU11dvMQpWufeSeDnxPO4ApZU4vcpbKyUgVKo8o1dsCSEB8HC08
ZFrYuXKehYGgkwgC0RokU3ZnEpBEwUCOQH9ulz8b9AWs3hTHMzSalQRZfNHxXTG6L4iCea9GsWLx
iajXDNVu+hRC3Ua1zJcIEB4zrllE+0uqIMUj57arRRHC/EoVabkbIija8/0ar13czholvH3+vC/+
1na58QfhghZGsPxHGr4KXkudD7S8zZ91/I9NHjqr2meyHaLfCrHS16kR/IjYj9YSmlgtaL5H/sME
Jk8P1p7wMpGX1Egeg/Z4UipBAG2RxHSEEgmvQXagjCrwuGf/4yEWqYEU6bF4EOjg7tIQUQT0kKUz
tju4qwWqpLI5NUc8qCJyWkCB2rPStcGmRNz1gkhAznam4J91FmpHqe5udxKe+tBPMgziCNgyDDBU
pB2ZAp70+c1tdqF25eHXqirnm8fX9LMOnOCaQy09W2AaJ1djHUqKJKNPhAiUSly6KTyOk4E2AZaW
ZjPaRFzpYbb9iSyq/YN71bjr4tXduhHYE5QCG0Ql1AQoQ7tyeOzjJZq4i7N+Llc5gchnxBRLOv6D
IMQ/2m/5VWKuqgRVfTn7cQlup0MWYvp9Bd7hUzXQNwEnBGW/IAUXrmdU1rJSP8Dm4i77yYBTBmaA
I2ZRbZhBhbOta6Jsd102aqcr8ImZCb4MH82A1j+bv1Y9v6i9zXf+7FSWMA13VOfzvwbqE8Rf0xpW
A0KD1Dum0eYVzfcII+f/IRhyTAV8Z9VA4mNqtc5GFwwSKCpXuaZ6fqZ5zFQYeJNGmXI9s6IWmQ0Z
SAePx8+4K5Tlx9vM59mLaUUs5GEt5q8OcyOO2ApWbboGEKGjk8KGrxoqA6/9wYHf6Rd2Pzm5A36u
P+1CEIvnQdW+nTFOg4tu6gmAPld/vZmwNqEh7ywiTMEBAUVn+ckWMtaf5SnwZo+gy3riSvX5WELl
hJ+8B7EOSWdOgpO8QJQGQ4mD3vppWfICCQxNBX6ueinVdLO8/r9QAlmfMx0q3Hxo0r0XG3zrx5Ao
gi0I3iAYM/DtW44TosBf2uwNHiaFjRvNgVmoxwoPGgh/irMGKSOdLgptt03sPur7in/oumWsUun0
WUVCqW5D21cJXx/L3o3YGS3YeZp5eXNUKXHyc3L8OfEfa3zGV8EJ2t5772I1YlPlEAbNhLokqaES
+U+loWiFZaEbmXZklXqsYju+PToL4ETLuCMS76nFNMnCXweVD2tREgKuzwv02cTxzl1lXoR6HO+w
Tsb3w6bOmJvLOUJaQW9KM8docDj3Ciph8biLmruFRmbYARe88gR5DbAOvUHC/3XHB9lhINNiIyZC
HX0bjBlDNmLikPh+EVYUYuK7HTGNNbiPS35taDM3/uq8/uUusW9Ip8RA/7bCHYos2wF9Ujoc0xDB
cGUbkhfjVGUFUnowoo/kz0MISOTmRdFivT9f2KcYrMyX7uaM5/KD0+WmbEHn8n8gpNDnILUWnxkn
3bb6MjU9AgVmWl8i705/ZmxV4KuFztsSmjnebel99PrITbugurZWbwObBJPsaUC196KAVBO/7lo/
pGLp7X/CzlmRD6zryEXaW4FOc751zAxXoxPq7ybTWXxDsRt8XqtOcru+EY4T3/3WBZl+QM89ZAau
AuazrKG1M4Md7Bq8WPDrWdcmjxzC4t7NEFQQPm2thzYFHBkPzIfeVyq5+TOMLXcL6E6Pg5zgU72b
KGJuQB+KL/UrF9LG6Xn1lVpbSBnUjEYNZ0mBbuzZ5R5/kmZ+UvCRCShalgZTaMfDynY+y0J4a8kR
KrUBDZ5FUXOmLppjB72+ShvFseq5ivbDyzxvVTqr+AmMdH+RH1xrEcp+VXnzMhDcQIiyDyXuHrWP
GHuhSTrVmhSUGpGRUOX300/ShIVfnxYX50LjbWdEzvhAEYw+Q8S5mrGqcggo2gwRdPwS2Cw6e01T
IG9w9zqpY8bb+1pfeVdqb31dlZT4fsJCG4WEfMMIz/3Jr04s9vVc9wuYY64v2e2mBFR6JKxU4gAs
RpilWQSEzmh9fOewNVXD6PmXTRyRER0vQcq0nMfYkG+JjzPstMHfS1qBqnBH6aNett19fa1NePF1
hm0/p+dxvcQgkzWcrLvoSylFPKZmLTRGvQpXMAz1fvvEfC5Wz3VWompUTwmdWeZJxeRF+Jz1a646
R8iD0DMWca/l8qg4b6CLpRdBcKYOHGxpB/Rd7XFozHEGAZW5O4z3641HvcLMz+Q5vHAlhfq7JOnU
YF7Yu3b/Y5UKgpnXmu/dRnAWCDn4sz0iJdXKEBMHH24pcdiZ485KVoLM8gLUK8MAqI1KJAi2lFnH
U6a1aRpxCt1W0ROzjgQKZRyZqQnYmLC3aO/BCDCqppqtPChICQRwGgK59zEMSXV4+a2iRg2WeZgA
MIQ6H2mLdvf/FY43lmrMGRB7lgWOwrX48yab61WKSDKZj2ScYYhG8gdZD1+pifBe9hCSobSDyBUS
KSJknrp4qQH2kbedQjE269OC9Nn5KEdvtmlQHV8sMUSCQymAuyGrcUjC78+nTOIAUHOq/qTULzGR
OpVyWJDyKG5KhFrSzuv1ZZiHpPpWe2qCvo9f8cGXA0X/04mRX6odhgxmsHwj6MJYlkEjQKG2FaMv
2U26g/BXLRkVLZBWd53pCKe+ceOBffXtcCVASlGh8DTNFsZLK9/BxWHql9ZvuBaIY7bhIv0EKdlZ
IXHzj1A+AeG6g/ZBX6KnDbTW4KQVAc5RbaF597jS0Kgt90wBTst14dHIQzxDAWJ5GoYsRmWtWMcI
sNW/bhf5GBkvRgyGpzwc23cIOwsHlOqCCqDmpNr3PkCk/UaYiZENKlrBoMeqyGIvhT9H57BHFHs/
xM4wG1G+niq5pB2WHk9YyNYUYy+EmS4IVFYEhi7cJaewGGGFoiv9Rr2rZ/Ard/rk4OP8HqToDKJS
qcmIURpnOqTDNXXBEpn3MY4YuqHnnlV5i9KKoSI0JcfxB9UgnU5JRsngvHeZxhMSEpZ7jYUwJEt0
slU0T4gPtrArUE79w8RcHzhefuOE1YUvc1/HFhfnJxEuIRYLhXQMjR4EOxH/wjUVR3qkd+hWrkzk
Rp+UqcLskLy3hWYEP6wDduJFZq3FzbAGetiB09EhruKtZM0b64Xgnko2JJ427KK5p27h3KsSWcCW
zjP+22aYjcUymnH21Qq+oQsaoc154DE6W4ZxgQXQS4rqcMLVqsmuW6mklgXRuu8S9cW87W4fL3Bd
drSMxdvilbRjpJmC+4hJSkzhFn8TAz4n6TM6kkfqadBtbPEF5p8h4iazt/bkORDFinYFhp2DuQiV
QMvvMs718YGJry+60peQh+ZO4BxSLgDXSbzN0RYS+vGaI99gb/85gX8A3R8gjj15EIPzagZsxBfl
mn7rjAWn4jm0ZWptYli8yQCkXBtR+GcLoWtS0nU+RTIzi4NqYFgvIgrxPxrxv5TCAWRB8WIgVwRI
nTC8lYdpRLt3+5UgyYxErccL6bRbm5jeRIDuIiSDLfK8RtuK/BwR1oGdGg3dN8ZKWtLQlTj2goes
MeySAt6mPjuVm4c7kblwB/RzS9Si8jjknIyexDpzyP1NeOUtbhrAp7LPkmgxJXkI13Kjnxf1jgRg
NBkCVSSRfbzExlt+9P/DutNFdHbGXU0pI+T1A+v7M5kTfMxrhSe93sOB4/xBp3i+X2eIY07WncpX
o9J4faL6G3kxfwbU2FZIaTzyQoxfqhOueVEDst/60zJbNwnZV9mDfKBjT5VgAICC4TKyDoysOQT3
c1wEVFVsdewhF2duO4o+YyphfT3Lqkr7aXENv7rtCdgZUtsDAQIX+3ouixet9qzvsgTaLxhD/V+d
9+zym2igU2JdyOUFfabyyGEjMR8gesb+k/mrs0nHLDLoUWKe7hr++vIqzYWv/NjbiXGxoBZ5SGu4
jPfKDwVlsBZP6JUcf/B3Pa+Z99cNpu0TucyrNtEE+Ip99dMRS0NorQfAeYrKiNmS5zRok1umgywU
mAg++7GXqa57xJiTMq3qmgCWBTan5EFUiwDTLyM5mMKZuvAWPmT7bn+aA38FrRbGPb7gO5ofaEAk
XIbqbyLyXz3kmfVUp95I7wZkKmduOusxax1aQRHOc39UuGjZWtxOw6OoC7kfzThPJCBjl+ZOU7em
XXQrTMV0/lOJrddEcAyhtLpiDNuiw5P3oYo5193PuN4c1qn7dZIS4BdoLpq+HsAwZdvwpv5Rj0iz
SJVZg72QZGyV07x5UX+JSQLj6ckEKDHvG0T3WHLVky7yFVjsC1s13UP5j9qBCgH0+IOrVjgnvIMU
82sGLX41WnrBlPg2nBWkoX08GG0L1mMldmASVxUYNk+z54S3M87S1tQP562L9XEu+06n29yjcpBG
yHwNQZpNs5KXfgxjdryNqggKGFHi7GZ421KOcPTNSqbvNk/+hl9l4O3VznYUiCj/MrXMWGdKlgnG
LR9sjmu2u4DZw8k7ozd5Y4x+0UcSJ44oXeUs8Y2Ry71yGj7CaC7nBhgzt5TVbVBd6YMPQsblF6cg
mNv+uKMyUrZmB6PRG/awzWgD2t2ZeCgr9fwuwCoemaNGZN3gy1oMFjcHz6DRFwjVZXLive6YIdJQ
y0EsAjLc9XgTokwPZPVnPqJzoCtNksCnLp1GfQFnO9Yl4EauvG7SIXo4aAMVIUirIhcK0fLBlSb7
QrteVazrz3H25yijWO8mlXU6FDrEvIz5dC1ZQb550vMUqY6cG/pJDnsPQvHHm+G8zQjoQPl6wgGH
8LV/woBOcF02d4IQjh1UwSLKdTHQrJGqDp0GTKQquVMhNtLib7Tga1+lXQ2aH3ndC/qUkzvJvzpC
5mtFOpZ7al4DWcWqlolh8CvasZ/cCjm6Q9r3WBrzib5cytyPY0Hui5BcpDacJV46LI+kW7kODU14
x9YNdVdjFu9wIjBE6pqnECcI9dIw0WFVD/IL83RSXG95bdtp3AVIo+w0LoOjmakkpFxADrHxxcjv
Kp2GcKWR3Zp8fR6jeiWwgFYuxN2hTV4rxrUoJJFNQjDQ6omLWCQA/TEDckY2q38BUTnYkgvAOMMu
D7P/u7BdKGX0eg6B0L/wYlskvjkuh3dSQ+3DE+cqB4aeq9eg61X99O+JU/wdzGyHuIj/GnLxbUAk
UxH55DDbKVj9AmO93pAzhBxJuERkuhKjRD2u5LKopcg6q8utuBPszk+W/+M4jBV/8lYe/N9AeDYq
fDZGEwEsDr4OWunYvpCuSS957VtWG2ZJksI6AVWpborWlPiFGu0H/YO+lE5w4eVG1Lt/DxzI1TUX
HJ4zcWPkMGpExttMDK90i/hs38fTptgrlr6CUJYFp4tfQgFVFC65/GdAAOfYWATLYHhzkvtb8VlC
i5SIxs8XFWq5E57SmtYlUfrEmkqSdoDEZ09QtSszyOW7uMQ3Zk4xPSm99fob6dWYryUViLsXyB67
IfaXI7hHU0wudbhi80u/ayuIYt6lZVx84q7VPIN6IjC+SP66eUgaQXjCoZCCvSwIlrnerFP/cqCQ
fib06MOVPiWJyYdOY7Rm1VqdRi9Zjgci/el9eYLvK4u3J5OO0XYx8YclmxRNz5qIGPupB6FMtSvx
gJibmVVdUYMFsGPBkFs7ciBtO1GmLBbUjrR8JLKJDo3xwJjWGSTSqHA2wT+JJwMBpmM4pjeHhk0d
wKw2eaRIChA62vU18WIBKbTXlWpEtchoAaIQzVAOO0w74HKurfVLOdUAkFZwFT8Fo+K2uzScFMq6
GqDXomDWZd/MzEDrclw2L8iAxfZYo1yvKP2gaDnWfutuuKVO5lvv+DrNjGgj9XQlB5KOck4zcoZc
FTlFo/yVsDtI9HAAwz85d2frl1/1T/KnrggOb7rH8ZoXcxGzA6w2QZjrJOQgyXGsW3jX1NxaiLdw
3duLZzcG2a8bZeTjsoXtvL+ogGu507nxPNFcx2v8GnGLRvh0xIvnDwliPcxVsCUPutACJ9S4Wpkg
+lP3Yn+tw+aKbUx7gwD3Xh9qoiXAWRxTx4ofKEc6/o2FHVCbxGXDFmf3Ec2k8IFPvTlr7lQM1GzX
w46waqJqrVlUBeHtf85EyY1vtV24iLe/HgKbHVzJ7R6AW1Vo1RbQW3lIjCiKQ3hgd1EI5Rf9H98G
o14LytJ0q2m+nuCWbi+jvu/v4ZAPoUyOLH/COyBULi1K190n4xf4wadfFSxYxiEcAY5UYXdWKlW8
SAqFlqkwlIjsEuJh/ii+wj/OoyTOhXApw5dWVYFm0+6L0TIJFLg4PDxKS+oOas+4s9eZIc1ndlMW
xwhKGB6jI0NrHRhm1j8uAmbMyeRW9bnWUGguNQ2G9gOCiw24elb6Yx6wqwkLLhA+gaLfOmSMiSvd
Zlcmuv6KQiIp43eGMRsu65Pli5WqmRm0Sr/D+8lZMpYWLhfNDTIyQSMAdBHyXteHRK1071XECYEh
vRZj6k8JIwEfIJ5E3zlGKXVW7X8qvQKhMJ6tLbEMfvpGibDRTQjZuV0657T05NDTHSfeKT0Qwp4v
UjpJMsUbibtAymEjDlQIK5nKU5frIpJlgrvjQbDcqygRFgOYmvFpwVn7e8+WNkByIoEh/rcVSmSC
fafXm5HI+WL9676Ot7HFpcpNmWWcBjkSHjTx8I9AzGdNybPGj/yQsPrflNDjV+kGOLEMfHpbKW7i
itgCGg+2245gHcKkWZmxYV3kKlPgFmPliNsByveTZJu20i+5NBix9N5hhRRYHQlxWyX/FH1dEIDN
4GVM4IADq4w81Y08fXZS7lhsbM4mGtNAtUbD1XKARuXRcdXvffne77HP6dwd4iBBSAh1UGfaWcMv
XYf6Eu1QQQ8bTdj+dLl9/DaYcEX49JcMuXPs5G1+EoFH5qm//UaurDX7lZBszb5W+MpihxLSXa0L
0KtB/kSul6Q1Ln8FHl9MzUkZK6yEVzcYn9Kq8vztrNgCaZv6aHuBLEgNAutAtoiBlrwdkRiGssVh
oBw+0jrTtPw6cdHCYDPI35cw50EoEvASIUlPwhpi8Tp58+ws7MHuSJU2Zh051eNSduPMIUtx8w0r
miiI84e/J/H8maUb6FtlAsonepoW8xILmxOfXWHVLUCMj/DqZKWkpRoFp2xksH6CcmZJ+J/IA4n+
tNsEt6xLWvvd8QdauJ32yJ62mQunz0mNXDlB5RAJl/Z6s48kojWc91Mgy2SN5z+4kBH1OfsE4/xy
tDEbaOKXhwxvJWDd+wGprA8yUP39uXua+bi6kobDGzoWrrRRj/6HbwjuUG2NCO2TVsSY3cjspIc7
T0i/hnm1MLG7J3vA4bcTsc6lKVDH1HJuBwgQzHiBKdH4KUycYErR5g48bHKUOELi2YfFFIehWkmp
0MhMdep5nSpe8uHgFj3+x4GYuUpmBS212mT3Cb2d1Hh+mdxLfEUJtMWIS0Z1Rv2JvqhSFEp6rRmi
HBvZ1bOwA5m380f4D5pVDSTb7yS9iUfyZbhT/gDC5iOgCS9JGx9/3Qf+3wkBBgG8/pZvNWZ0uqkX
0mOFQsUno92sQNgeoNBu5QLRglYKJPJHiatCp+GculBcnHMFgHgZCT/dG0sufCuwymqwdj1K5nzU
YjDR1A6qneb06LPV4vGi1iGICYtcngFyFJeyOGiH8XDIh/kmu9EDwzkd6eclnDBd8X2YHA+1wV8p
ZK0LymgWedS3U8qkqlDbyFqIDXc4B42tWVYicEaEzVbKkDCL2bSPjzye+T3UJCrfhv9DG5385td4
prxyM9DpEKPIBg9u+A0914zOoDkzcdwt/b2BawDglySOtRU/49amK/Kbj8wH8eAP1wnh6uAmC9m9
2YFqH3gcGkoZJX+rm55RV8LWo1t6Uk53mw7joN/NjGgyB+YmI5U18AUfzUY+J3ye0ocGty5jiXLb
4CcL86NPv4yFpJ5u3IVL9j8gnQmsbZCNG+V3tq/VrRSA3xIsjXgxFZSvjf95wQLKTJPzwRVt/OH3
y4dv/oGC+wlYozOH4loA6hXNanSc9nkRR0LyaG+BAkGyTmEqlSdqYAMgpaqpR279Z6ztyxox0Ff7
BgINQz07BJMhxkJKg7ygbb7dA90QcCd/Z98jZkmxptcx0Yg/4uPxsMr2QxtZkJ5/Gb0eaNYCREYs
oPcYSdD5m44lNc2Spu8Ke9qhpeewnk8Fo5QOceD7QSmSAT0g6TDnR9VJHVQKgNsgMxc4LScPEs93
tlTX+9iC6J8sLeF1vnocRSFNVRWa8EApljG2CsaKFRo3HGRkyXCrdlrDkPSL1vVtIELZ9zIvV+3z
GfpkaN5Fr1cmHG5JeYBUu4+Hh8U9FRurRlrGnOawfZVJwed+PRZsDJ4m13uKgY89RgreWeZaLjYW
Mc2d3ObqqnoOB3+Vo21e3RKFEJmbCUNeZF9XcmR3VpTW8RwnzNyrUH53iE/eHNs9EISjuZyKin/r
O7cebUpsgWsORqYsDj2xfKSQQ/yVOTmh2QtmBlqrZaSvEdn4eKSMg8vg2bU6FnyoLh5K2ghChrPX
gUyF7Ce3EROnsgdY7NmwSraeyaxyPC/np6hGnpLkew+ECG6W04c15v8MkC3LoZ6LyX4e4naBCfqg
2fQ2uFwcjaehYG3VoGUotNB/QJUSSV/Il3cEaFbreWR1u1+PFbj5pNn3XDfl7vDjmb8FHV5ZcRKU
EIhx9Zl/Bs4fHLYbgu/SHLFztKuR/aLAzS0bV6VPHfbKK0l+bRZ+YU5iIIGVPobDTM6qE1zdbJWo
pKrTm8tMi8PuoQ+Wk94A/zc3M5RQKM9ZGIAsYoxJbIioFPSxRO/9ddtYqjwDQ+QdoJn8sK11DIGk
TFR6zP8f0L0zHiKCF06oR4jFXeNcpLuEmDKhS1a2fSuuKgu5p0m7h/jf3z1aYZItC1u99NzRp8Lq
td/wWqI2JdbNlRRd+oRBdOnSBh/7Cd9QtnKaGEEWWpCWtfnnEMJNtCOal93tmsdiS/dglE+Y1OKo
Di00ubnB5i79CArSSHrUSB52BU6j2IUNSLOSfOrpyjqUhyb2BWpqU0LMlJV/qmHIZv2IQcG9mj5B
t+9MhaVvx1uJsWgMwV5iSa4X5KdfcyuB3ySJsR+j8FlsQM3fWMYbxfLcVDyU1lNFACa1CuRMmhHe
Znr+tIFnLfwWrTSWdbAffgjjj6vQrsgud1hKYnFVLWSMrwTzeI7BINmLPasM68QdZY7SvsrCXwZJ
9Zt2PuVQolxKPUvenBQBcDAi6hxdnyk+oAVh9mpnqDZzapoprFA39cxlX1230qhFZRfhk+rJJQEA
OOKoC2joclDr+toWorGO7v8whuzCH/XthhSJOs/eQl1NAFaZXRrZBklR4gWBMKG5flac2QDyIAFc
+yMewEsZ5cjEyYDWmbJCdMh9cNSLm4Aa0cra5ucHLpvlzJT5c6w2T9I6rEjBg2iySt/eGcSD+VeF
o+gma4AsjCHp2UfEuVKoyIlbMLjOVFJhCTUR5FregCAx7doSMG2r9ksFM4Q+G7MbsNiTjCG1DFKn
R4Rynv6s7Hg5xvJlnb9/SEBbEycHCL2dHeSMeQ1WRrbGOWQ/M8PxQtAeljE1hpQ1aLmzHajJMdQY
nsO2fAy+50hzP0s8U5F9I7nppBR8i4+J6Tfaxw7otg/vc+wlBOfJdbSe5qjPIVJX3jsbeQ/eyQSq
w3i5V3EZAGxNLh4QHRjozzI2vKWIZjIgXLCDtuODAw7eWurRumEu1ciKLEsPrAOUXAsaHjb2S0AN
ICWbiEaMt+Dsg73wT/9WQp3tL2dsnp28TCBviRp7nhWM3YfYIIAqX4frnUIgyzn4mPLQlbxINIZF
9y7m/+DNDGyvSJS6hawfgVGBJuh3tPYW7hf/KPMlAFluCif00GlKwfnr7fIrtCd20iOc5kG4390g
MpL03+Gvmq62qfouIVSmWngbk4GdnbzDwkAW89Sfe8G9PLoDtHOLhxr4G9DKocTDpWWKHGm/1tbM
Daf7q03YbflbYmDL7+RFmkJ10DwK+MURZ1rBAa3StCE/AfytK/5xYhSVlDJGnfhyJqxzZelJ46Rp
4Efp8emiwm/XFej46bbMjNableXjQ0Wczcx7b/1qw4WkbOM2ptcgTozk95HSu3/QyEb3dTbDoeoP
uzftdTV0uxiMCMyGzq3VQIUwxkWkHRiyV0+u0yunwW7rtCOdh+cl4dBRt9IwgibIR0XKLfar+I9T
AMoFTe23ydksEiFEIbjpmVYCsIkn6qGZha4iSGvlW4WJFGzr6exlZcrvK/TU+/a6DfFFNs30Jr7C
xmrRPB8whbMri3v0KwZz8UthVfcMssnXVT1YKIhmMTeGe/1drgI7Q7dDpdQaUHXkGWrzlRFUbbaU
KJfq1sa8SRpf2zXgZd1FcjHAo1rNfjoJROmDHRpcpMevS8hqKztcB749h/PwyazM5J83NGgw+osv
XbUqNkxl7HcYUB92kz+7C5zpBUkcIVcMNEDoEF0HdM9+HpTpHsDurwCFQBWHS+uxMrkearwI6eNa
/9ZqFnFqfcL+DxAruKnLJj77CVXZDYIKEnL73qyBeoHm+i27sMZ4mqlZ5Y3Px8fEHr89kxRx2EPr
YOt68ZA/NEhJ/3emptinzbQ21zlAflnl/xs2r0tc2Q39qPYDWYWotDsGczH8A/ESE7EPShyV88mc
OAZ3bMXK0NlgZuSBUbSJgsOzxj0yvW6ins2E1d8CpALc65TPDO9YxyVwwOWcMBEAqyZ3lRHPFQvN
gmXm974niNLsoiklDRSH00F8ZOXcNtzDIEO0rFZWeAcZqGTU43DNi5Ie4PH11eoTUAc6X8cmWyv0
Avz1ck3LrwAGdueLTdXbw5dD3mIv5L618aA6JomLTejHjSUVQUU6lzVEjtdj40tuBwQ9TKvhfZpU
WVLbuA9VfFrYqzavpKrbjey1N5YbLM8506uTaSF/NZkAVKrcw9T8JK+s652xoYuvTOEkLGlbRA2x
8a2mbP9n1w9BZfaTCQFjCqQGofOpiTxpxDPgGjsvG0PqJOfKi4/steazCrTvVixK78Wyp8MjU5fO
4nHowIBWwm0US2kVR1S883guoSOmXB56/5G8zGswWmq8rNg/Kcj34cn1hc3vhFf6Qvn9fHUlBxLF
9OsYYB/q143DFIhMn+K9BcmdLF1XT3rzclJmyH0amjGZfJUuJ30ln2gTr+Zk/2NR0/F7hJzm8pLQ
jidrb8xHj0/Oh+MPdI767eyd0LkJ4zgQ7prJ77LmSdYOpwCanP8XVvut+fgQUzasyiqEeWedPrQK
oBjr1YZPfOqLrDfEJwBSBV+PvQD5DWh6MDdW5pcgAWXaTv8ciUJYl/RD4YgorpVOqltwCNfLYJ8b
RSZJhT4+7vnBrF6+poMmB5GSJ0/HkMAZ8a2fPhHmouzMUoiOGwkl0VbpFFVcqFroXN/TqiAPxfol
nB1HBnt9PWzvDFEKUBYFCGdBlx2INLOVn3i/fKtrUI9ZMbjcrQPvNcHauZCx8IjOitK3MZpJZLkI
2riYbAIE3VW9mlTMuXT621rvO5rrmqCICAMZTR4HiVGzCD7kLArssxIb2rk/erArVMxbolR6gjix
25DSNJc+jZgpPMqjydABuAqTUMjUyV44SSm9bMEG26FA6e1bBp+yVtuGPkLbdSRW0C2mybtvN19o
w+KRdugDuWrN67hydVyXwAsVPH44mPE8hqysmMytOlpzuih+RcANrHLrVRz/GzP3Jp/JRxERETrr
EIz26H7d/kSx104cyJBT4WHasLGChfIz/XnG9tvLvpkAMMr0bIsYrj5hUwJ3C+vcOM+45aJmqMCV
y7hEbuR4JgwMjOBVqlqvhgMjHWRnRk2IRNRJcVbjptTY5rgbMIxWz9P09ZtAFoHWEBPTnDzd8V/v
dQIS8gAypk6ySbwWvnwum3G0Ons67EEkYPCxBWpk0e8fcqhgHBMNn6vDpUV5CJ5pBDXzXwZsOuj8
i8KHKG1tL6U4SdfmcPDQozR26e9ebuXEjJby/qwvhn5ZP3oO2xQzGgcdDykh9Pl+MllGZlzWEueM
GWM7lXlRlFY7nG5QDkgMTEBjacMsSqZQ4NxA5ntpCU9pASeiJcdOWh7NfFzdjnT4Tj8iSQblFp14
qPY/GJOTmpcRa69P4KERyLVa88JvU9G6k3GLg1WuFDSxON0YOx9lomUUgxQtx4A1xYphY0JHCa2B
ElN9RzZg4dkDtM0LpkxhQfA1Tlr8D/s0AZnaFuFgo5qykYzW+WuBpVD+lXpWuDX/oOOOrMgm/mkZ
cbTnUeZPkqos4TqZVfI/qVUOYKpH5hNGzz9QL8p/OgnBYJ2QIRYv81nkmtzMAYzsI8qZKSFKLGqI
QN6fjB5RDOOvkefJRK4HX8+aa5SUFgbhPYLPZOyu9kFFsSCKbtoa6dHf2MJ4flqQk49XATZzrBKT
q5IrimL0FcArFxs1+kASsydq9uzqYv0cubNh5NJA/0ECkPqzh1HW0WjnnfP4H3oLNeK6MuGHROW6
VLT1IE4jKE4TJq4u1W2XvznsEAtjRGJauNwsRkuqwfWRIGOAYkDng2L0NrWHXHQd7nEJnojwjqfM
Bjc1Z1ZXjD1lCdH+1RoqFyFMt6HMEfP3KR8wa54vMhjoZ9o/XI328FryU/HaMgpW3ZXT82Sd17fL
KHjNMfPmEYpRR1Wck9/KUWEhAzH3tayd1Kc13OGZkx87XNd9xAR78k7vJdE3oy8FqWcUTkDCbAST
E/wyEJadUetig5XpLbo5lrwmtlxB/LNATajLmQPwmADh+knmHevNF7AFf41gxqKgBf+DuZWnu9Kw
teFeiPB8g0KL8+e6/3W8oRoy5PsgLN3czq4cjwCRf1G/UVb7GRvune4vC2aTy85OI4dKbJYNCfu4
qSedcZXhK24hgzZE3tMtF9Dt4uncwqsguIr4e65iAnjT5/Og5ga5ZCu6ITwlHMOWlcsjILQmSrpN
z8zoNd7SGDyvMQ12E+uj4aVyx0L4a5dOqigZvI8YBDFTp3h1vGFxnLGqwDJpldX1UMV8Bm7X36s0
S7Sr8aQXAo7ZlHk5S89gFZ5Zwb3RIdgO5kGEZcA+uTVt7yZCP8dLN47ojB0Sr4LFLp7kb1+XU8JG
GnkhiRSHJmq4fC+y8T9ctVNDpzvxO83ZIaTc/z7t+VtgIFFzJHgi8aL4HIm32INp4Cd4DPDT28IN
OUmlGIsHkH81CxfjkSG9qyCbSXN5Pv+4Ly4FKE3kUhqKLryQg6A2z8YfXyBk+a0HYJGhZPaEl1wB
Aj5Z97uEc0bWLvzYPb3bzpUbcAIEtd9FEoaA+jvjjMCpPmu2hqO1VOVhq8F8niaY5jT04TopVOMM
vs9h0VZ0Dc8DUs4q2NMnznM1HmagcbZHRMZSvY7gTx7p3LdILt8P5rShe488zf/fJBVd4ISXx+G7
1iErrXMVjkbJk/6RzhOdrtFqs0K3rvqM/+to+mH+8l2gayVZHi6ebu/WWSuyCvOSfroraq/9QcSf
OimiFRJK3ir8CIuCDRpboRRhP8+YaLn4xkbL8Zgi/mhn0idoBOd3V9YldPJOP+RRhjLZ34viGZI6
/o+TN3wufNo5MQueSHVMjDu366pVCYGQGbInetRXY8Pmuqj5uHdsuU7mhMWLFimk6yvH9w6u/xQh
0sI1qAMZdqhN40M6gat14GOpGJJ71Icx62CgNmXOlwH9KZVy0mvPcSj5TBgt2Znc3SDz/ynFNIP8
VygIQTAtUYAD8Tjd1MYbLAer/Fim4FutEq9zhZD0O+SE5b7D0GRKFTsVsVa4ImodqtVC43OIXRo9
GzVczQElo/TkusyEhMyh2m/0FuFwqLwRx6ZW1jTlpjWdUuBWeftFD21vWvqG0x2IWTStfXGpBlss
LHDhuSXiI9oCTxQIJOuFnXAnF72xE99yfDbUviPzrhR6s3tA0FAZUTmyPSfzIWsrp3O2YkG42+RU
ymipa4kBqyNCMMlL8utxADrMyVcWij9eMrvF5I53kVqBUJyeOeN47mIFOYd4XGmwcy1aYlXO/F9X
aoySG8/MGo26hXw1Fu0fWlgzbgaw4ZpGxog4MuMsq3Y0BP1rrJqA+dvy4Q9NTr+hlD4UrQ2jxKII
FtXlq7csPgXvhbMs2AJp6NbIyT9w3Ou/itOJDy2VI/jbQEiFIlv0swXOMA1GcCufXIqlGZLiGooO
rxeC2Cxqoxie9D6E7of2B4Risxj11Y8ZEDv+PvvJKnYyThgglMlj9kasL6QTPvHVw9hkNFUq64ki
pzyMZ9pa6woHOVL6lk6LA3BLwMOnrZ9vFUoWHA005Gv7Ssuo8Zb3FmAiRe8+sr0kdhA6IQKiwDW0
Ls1gTMhd8jVUAcDR9BSXB+0QUBFRVZMQ6+B77oCfa5ee9NazDmOmDDoj/5mNm+Y2QrFbhaUkl1wS
J4jR8uyW3ojZ1kAi41Kdl3ZVtW/HAzz5hz4gslp0cmx4HJlJqx5NEAHqqVJWHzoTpv/h+5oqqlrR
MgmYiKV+mYQqifxp9R3gCuS16JipWYuVx/nI9bVNtvwsmPu9ilF78hr/Dt7x+lBlEUX+KkhWw7g9
AkgDGfvfMCg63JDhSJo7YGN8nihwoWpBNT+82sn1TNzxQruuo2r4tfbjIQRz6K3llNtfDUftz+od
yhjcNZUC9UXm2p+vS3fX1k4QYzw9CA0yt7ZJ1h/Q5YfR8lYpp/8mCqGTt3o/i8xvW1KQmJrfcb7w
oMa7/JENqUiYPRDfzV/lXfoUKPfsMiwnra7HPH/fkVIzJVBr9e8hUw49Yp8pSeKE36kNoE09W7is
QQf1/qv51m01NhS1zQmIDdsQRllZvXjbVwOJVt2BfuhoMMITpwnuW7vhCUrUMNkaNYCjZHBlncdq
6SfP2gKd28SYy6s4mkjdPVSu82F1ZJ7kMrL/N/ucEwXacqHbNGF1Kr+Wn+ZnRsB1ebGXNZ6ftgkp
gEAnEmaJMJhvcpSHWls6WCmgJbflISJkkjqStj54VaevLXYsJsKPs7JGUDpc1pTvXfsXyrtSdzX9
BrPtV2/t/7DRgkmY2GjQp3pMJjOvDhj+LF3U+kvyxwhNewAPCs/X0LpO8hKyhhnfZuNM/ey/uIos
a8DXZ1+I8FlJUs+lLcBNHMlFEVzyQDRgE25QkKIH9kAQMSHPy9h2Cj/6XZcD0u2rg8Ml4lBSiaQ7
2Ps41MznCdyOYQwpNhofO0i4HfZ+t1ejFDaVRTmCLgq8ohIKomT5It9DzVqYTSmNjrNWgmBe/HIR
iztyWFsrVQwreP7/SGq3lykkWsjcS1ujEsv2+sVA4xl7fVdPuV4MEw2kvojXVo7pjaRY8GS874mM
CpQNRToyWv5XZRWOWNtNg1nlBeon7z7ia3HF0BUP0cMGBDy9+rN42v03ogWy/mkHMc5S6ETmCR/J
ueyGWm/mona25As5bhy9H3djziKBecEb1gNFEqxBLt36VSAXPXHLgwKdhqJ+Xu1iC6JpgTayL9eW
WjBKkBFK9CgiTTZyWb/9S8uLK1O8WIREpDMKd/JjHDByDjIUEZZeLjYP1PGYXWWsdbEJ6oxlQ2HU
dcT65eRABzb8AZaLbkwJRDr4uTo1I8WiRxoef2M8WLao1XTZ/wEw4H/S9ghuC3AmTZyZZbxE1dJE
aCSy7wVN5CqAndxY4E32sSAh7ZtQSBk3rwXDH74NAj5YiQeDmvagU6KU0UQoPnrC8ATkELTQyBsf
9whXrEF3KNli9+hH9nQ45Anpi5C8QzfcBiadalQvpkDuY3esZD8ijP2PI2uSEQE3FIWg/UnmUy/O
QOlRGzt8oNDDVj4LSLghxBILf2kcVveegGSuZJH+TVjax0ApHN5m6zRVSJTfR5XLyT3UAuvhI79g
5dMyky4YM3Yo6hyKxGqq9CcR6WdJnlNCJhN16imsBVlzcxAm/MING5tA6/aelZEFj1bO4dMOAVwU
PsbrpayhE2xMQThmClXnz/0nx6oYShQWYmiaG5If7MEWingucluZe+8j7eE7+tRept4NdMgrZCT3
io4CyOJuI+oLdJtARjUntJ3iPDkw9YHBl3Ernws1SLClKXfgG4c4T6gAA0cLvevfwZC+v1i9q58e
gU0fwjzUXcX9ze8Uk9/XbyT/Zp1f5CB3r/Kbk8ilZje6tewuZyPeOvu17CZppjbb9ksI2fNQzDAq
9mYhBuV7RQxSjWYVKmb54kBNlzCmMyaxoAxASWHff0PBWe19rqcTpPB8pu6g+d8/ra594zJwidoZ
cnP7vPcm6D0wuSvwexTbAN6UqXlGsMaAmQL3UK4Cg0ThpzXMV1iOM7c2VGsK53vFN9EitcVq/U80
lpB8IcR9w0EmmhAK9MpKuH7gHFS0VHkq8ruk3H7cArBP5j1rNhb166GeISlv3km/gahyIb7EZ9fQ
lmlsixy7MSBa978HIRXPkZCT62MIQUG6Ivik1vyAL3EoJ/52WaFk2gN/l3a/ieH7CyOQP41mTczi
pbcHKpptGvVyZ96UqBQ3cncn19dWAwuM2J0/IfdSyeKWPckeYc7sxmCzP8U9d/DbOSQCPW2hDQfA
SlnM8DpUJSVFGtLLQo3KOh75+uH1LGnD2bKTtMfZsZJfAVlMqezhg1PSckWxEnAiL1F/9ehso7Xt
UxHCS8994JXfbjKE3ypXgl8DIuZGYHUBFCSkoS+KPF4omKmDFcogZwDFtRHmXSjtoZRzSHVs63Y0
xywjniB74ULX6zVfxS1ocGwWWfRNoByqINPGi9TCG846VG3gHGjagjbC8h7inGv3ycoS3mxTIyhV
IbvpFIPETkEDeGagomTwwxyM1hRtMVinEUFrjdx2gJ3IjRQUw9sLsr6rsGzuYfCbEBceYrDYw59F
WjQuoqkQ70Ml9apvE0B7b0z3//GSZOwPg1yBu9SmdZtpi3stIXP7J2QO6d3yKYOyfXB7mhfPX6oT
wGwKmZKoSjLh75B09/perD2udpVIDkPJh0vzhRfafEhkTs2Ob1SVqIeksSjJBA81dN+1fQThc0ne
+u0pyiHWu8sjgf88uwwj8roy69xLxrhuMueDPU2clG0PbRj3BcO/yGQ2GjPnSQnEQ6NQPzcHdNIT
tShbtp1COLE5uhZjkCb4NPLvI2yjVWxmx4KtBTTWoafSG5nhFS+xNeQ1aFX1BneXNErdkWN4EMMH
OKPJpJY3LOAUc9wR1JFOLXmAxoWxSs0eaROmpOmQjii7q1UfwrOT6dipqB9EK0TlsargJNixUudq
sM+tYM6RnSVDOlhPRQWHPg5zUNd1GPdCrWhCFIkkhis+TympePMCYVX2iowev5LSMec3oCioN+Zb
2ZMmBbhz/QzkewSN6c+YLb1OnnsogXry01X8FCbCT4DZnTtlU1NE8aLhE1RpNUv1j9tyCxFfo+vD
eIHOOtatAAqgwn47O/PnchgxYpxG7oe4cAv+O5jmAoUpO4KlB4tKGmS9CEYQH8sBQ0oLLsoO7xv4
+TcaOxCJEtrln3UBnmjbOT2OkaH8FEpaTIA8BIgd4UhrJ6jIIPiuTF9QTHYkdKqVVmEnSrWxMMr6
WfySml+ZCI9JiI1xFsBlpJlqG49mQfAhdh6rLyi63SMm2+1d9/l9u/yXnafuUcSUj99wNYM7WTYY
ufipQna1s7qPP4cb1lmKzhQDmSG8KnU7fRH+DOtpyyTKhQAE7NizKtJsYwmcmM+zzqbEJDU00H5b
VJffizw3/h2VczrfXkA74aBxo702Ps5DG3yOBNxsJI2RqywdKS7YXF34zkl+tfHNlYYmSnTuvc+1
dPRfezvYNVOP6wD2XR8NQ2fiUeoB2pfyAg3hKTZRv4azmECksu9Oe1FW0QP10BN+4sZb9h7WkKNB
+XqORdo7/7J/HPJ6oqDa/vLVuqn57zJSwpr+S8llKmE2giAOSFdV++qoSP8QR49d/QWMB7uWWh2f
hJrfiRbJ7NStCLYsDVaLswARBgAYDerbYAP9QemI5lRQc3g7mvrEXk2x05+5bRa0YxEdAQEdt8cg
MpnnoruDzcHVWCs2DWsMvIIRHwGSqA+IJH1GOy6h7q5BEjHJ2hn5MVKLVSkMxFGvjpIwEH8/iI2l
bbmcy6NQF4R/pegSzt4nFyTd6xj2QxFisYgBe8iVoNdZ/CIhO6bKFZJJooq7z+9ckn0Go0ugBtkM
aVfY//ZqIvpxDzdVlA8sxG0P+66c08rHi1dA/nYXBWxEGjUCZ3rI9nKTd+MwvpWw7KEDB4c+JbXo
FN8W2ck6XVseFChsAbPdaXtGBIoJ1znSXYYtyg7v3xqxYzM2pstWUIyZnV02dnfDAdm2I+Rl2nKu
EuYTOHwCPMVv/qgRvWU5VUXB5BfIiqaBT+KhJnpCec1MHmZQqvjttsJuaxK+wZuoG+mH4aI2NjC5
SnatYZaVR+C8TvQEHr63082HqVqFSu1ablp8upAV25tVgu027wanrJ1T3IJ04guIYjAMIe07yUHP
kP6Rmx67Dt/+lM66yoytvqSfaA4qAVe7hixW70ilaerYivYf6wlWZ0BcEW0F0J+ge84MBdbtTygV
vwajvcbeywEB4UlT4oDzZe3CXULO2M4CQr8ZKS/vTf1qPFUbzEutn1FBGa85QSQ98v1XDpZEL1c8
7VPtuSjHbs25fqDlrbVktRTRqXTivuvls6RUCcVduiOlibR4odHx4W5yE9x0MuU+LXTPeufnVsSr
/rD/TuTNb5G6RFekBDc9Fmqrm0Y+skrH+emE0JhXfmXUkEUWl4SJ7RJolHhcI/HDAu8We/7pXaVZ
nqfVR8PJ4eJJJbEBoiydjFhgZV94rhRv9uJzczchDoLSqLUtqjHNfWlBJ88+0zUaeg76oZAjFYdV
vtGdiwXgdhyssBlzk/VbDelEUlkUz/+0V6sNTjDI3sJgOShfXWFPtsky8NTvw5dXfveEGXFDnJ4s
81gXp7XkTsTJUVlH32UAL5hWnBkkh9kBaxvag5t4Ymf9ixZvpsQVNP0QZTylFBF0rYfjZO2qdemo
w6ZDkJmX1nu5rCA/QC+6WeDZ4xDVGGEPzON0ZLIdMD+wJ5fSD7YFLMzj5VV3srla4zbg9Bg1z6aa
xbZnKSFDcoP7jsxlFJMcFQvDmxcAhvClvG3NlkO8OWqMQ57UsK3Z1RWC038mUnr2ZvcAZUvpQgAG
zFZQ9otBRCmEGY4suXRFpOz6iUZ4audw72D0ChLgs5RRMXOIj0CcyoKoicgnB7bGrMI51XRvEwD4
b0ttWcbdRRe0CXt5kK7LM8xJxenbkzGEAjAk/WOCUsqHfqRvnk8A4QA/CZh0mLU2kdqgZLWME1Xf
MReVNDpPJlKc96ojGoLNWHkU4mH0QujaNrMpRXOcj+NQWxFx28eQYvoFRLh0OSFjpbD9ousqXtxd
VAd2Ex286tr6SSG21D7cBYEmZkgQsT9GDdkuCQgrR8SN7wjcLmM5KK3AYuCIK2HGF/tnLxvMPddh
yLqrq7SA7FoysZ60xjvlOhm1fWmRFdNF1oersMkDmpipNB+3xfk2AZu85eiZli20n87RQm0ks1Fk
NkznJuLEGXYQQ3GjDj24WLYMznrZPx4rcwMd+fJjVXmUCCmIOa55mcaskeuT/kipNpaq0OuL9ruI
4FsmAVuLfrnhP2PycYEIxQnh2CVuJRAGiiKCYUuTU4fNSjdhtV3cB9Z8OPwmcDCePVgS46T39KSt
sGhzsDXplsY8bjtNkzIySSNvQVwVu7gFfyBoxKwPtk9Qx681pwvXK+f00fYmeBuPs12vrQikt455
jTo6bFNAiZX0NWZ1Yj5oXG5TWFxZ4fjD/U2WYOwl7/bY/GcBtlnMlDowhQgGDtKl3H1UbGkaVuCb
apwfUzAm10VjCZCXJfDJz0yPcL2LUfOL9FousM+SSavIjMhleiDMx6qN25DK5GhxdBZayaofJiJ8
syNZBys0Q3Hujy2pohYZ13TDq1yIFbbUiDzllFXuu8ej6R4Qz5wdZTvDHFRlLfc93rnt248cvtbR
0NBVk3RB1EHbeMqeq+qIw9OFVfb5ilLy5tELEz4UZbf/sRTaxiHPKC6K4WSzt5W0Sj7rRzoOwBYF
z5avyYOVcPPShBy8yaX95NaxeowBzC1wYc1f319/7VLObjuk6a60EfuZx2dbP4j5GhtnHhYmZypX
LRZt0e1v+ILOVoDleuiQsWEzx19ih8mP/COUSeZSTyGnH7b2StpY3R9a8cM8ijWCyULCf3eT7hqQ
u7XK1QABc8+itd90aQeQpJKi1ZMJJ10QlR7d6hOsVzQvmrepfQOHIFGs7MQE2ZaIdj8bfG6bw8SX
7nqJ/fCw7mydByeC/JpwVrw/nqe22Nu5ulFqOm8fw63qTe/0qpYFupwPQdaS6NCQVUUWD7noqA+t
eC3raq683wkyM3OapFKCI1TVo3AXeatCmJd+XwggmH/UakCQzKDJuvm/zOdlzhEx/+Bpkll4JDTc
APKvE5GeY1VuUxnGL7ogzVfLz8yu/KE/+lubwtQAWxjESQIvb8+cS9zUJMhghaY46DG89oDQpe8Q
Zz8dws9LI50AIfoyNnw2WbEh9A4ZoSvEsyErB14WiE/w9exzZ6tQqbW5LWzsNsrNpgta/4kfwqAM
BY1AFeC0aEX945SvxfLVtVbnynhwwQ8a7zwkhcwCHlF1qmQdwbV0OTe8z4d1nGn+6p916woSPmJL
5SCauRDBx7SWfjk1cZ2KEFCK1L/bEBaxM3uOS34WV5zmnE+0BB6IUBBmBaVzyZhY556A9tfv230a
54oG/DmukVsycZ7jR9G9jdwgfTLtgDtJPgby9nNS+PDHeBlJeTHKqG2jfE8BrLh+R+/9adKvnKrI
3VgUzx2rBi+bbOGkKS/VQB+NCWqbNn30u/w8ZVKJLcceNPJi2eMu14+i+wtC59rUJdrhkIL5TQhA
lqdKKjoiQxomIgt14IwweCPOFrUR2fM+CGK+WQgP3imv3UrU4GEXoia7HsheU4EV5szdbvKCtMQF
dtDRiRTyk7ox6MVlo34CN9G9szCqymZjxGB3897yKSPQUBuFQmg/w9ff1e7s486cCBRS7lA3lSN8
j1ju3D9lQAn1KVdKKTDli6eZssaVHrFuRKA658lHJL1dQ0efmC59uq9LAWBr1wgmuQebYxNqp+Ym
iYEjpnyzsjXZJBBm0mjuJIkhNLr44TT16/3Pm1kX6x9JR+GH4nfoUHK43T93W+9L7ofcZr1DXCUq
OhtNG9naog160HoJB+IZ9YvmyCyShHwQ4AtbH7nSmZYOzTPtOAiwGVmco+iKmWMm56+z1Z8mYuIJ
Ka1hiPuqRG3QHYxAvqU1m4dgx6AOC0uLwS35tblj7jJ8WuUByoDqmiF6xPwzKzyWQ5DBvZyUwVrG
O0waXpvqmwkJ91pZyoO985FZAY5D6NPsTwJxh6XfNa2qG15vAm8qIn6YVqG/lzKAMY3j2UD0YiI3
kKaj+4WrXj1SZnTtYprlqEmZwZ8XnFeryXQ/pLLCAQ6wGju2V521jSUIDC2C7eFhMFxpAoE3p6ER
QmPqtetNYqvR5LYM777/QSHTS+Go3RACb8Z3Lp9Ov4Xm+u4ltU6rDdRY9xFfQOOZxDxhOx5Jyngx
kybQ1K0VagDPseH36K1WP8vKD6STg0ZuyZHVGdKnBwULmTvo2CtT+UBRw3pnrNuL5R38sMHlyPJ4
P7NHxjYZoKdBvkwp5ylxkkHKaF7nGHW06hfamVynyuiSP7/PyFfBzZ/T2Nz0fcqJjMM7rBum7OUP
ic47QYY2LnJlJG08LBKnqboEkVmaCG6NQ7rr6txIq77Nj11nFeDjaA88JLc1+eMbDkTkROO8EULe
MTZcmDxwnGVzLrrk7/2W4vYN64Mhj9NR3TQwLUBzJcMx9TobFPliFXQZyULhb3z1u0PX0ZLxkYgx
hemf9YnC8bgax+Oos6yqgAwkenNiL+XmONt65sojHGtPfUyBfqNBJX3hkEnwPtdgT/yLBa4Y5TnH
YcLW1QkCPwMJubE3ZGBLqGDhiXYoN4QkG5RV8FNTVB/M/3YDi2kgdCP/bzCwO86jiPRY7tbyMvlV
BGYo3nG4u5hY8Xj9bz0iv/6Dyt8Xpb9eMxAX/B6gNXkv5HKjAKlVEvccDCW8LBhHGL0W6Z4i7hxW
R2HCFEN+lRBWy33yEYmiYMJKUV0Yq7ExzTZgvejRu8yedH2EZRD8hiwJkUqAZovtBx2zkqIftMe0
qBAwQ5FV/42ph27fr8NYwUyvNDuMIGuzhaIto3uEn0MEbJMfD0R/O60eT0NzmQmdd0SEKDIVSCEY
oiyHENgQ+DeNZNv4Y7tPEVSBFyL3iD8P3PCwXa+JLUjtTmCRd3fBFMPmIc5DpDHrNmGnJsKkFWei
ae5Vt2adxxyqnPLECKX38vLpzv52U4nbM5IeibqGer6t0nuHp+MoUaj09oy7cIR1CvWWnUo+8bx/
Np+oXVW6PB+JUX7kiDra6puLlHp/XGxYfJ/WIWFGq3SWCAI/r0nKNaSLgI9qtQpKqSPb2+SFUvwm
+b77/l71lHUxrd1OCRHsjmkb8lMSLO5H8bomFA3+D9Ugq/S5t9bc6I7vZL6f60iFECuckZPHm+Z+
69evg5yHVwbhJf34bi8Z6ywzTDILEq+E0/bLTjDFpoXifZQfn+wBXD2e0JZJCZsxRWIqT96K2m5l
yMcePQ0aIyGaBAj/6AWUnfpt963mkoGqCJ9tzZr/Ypu0qDPRObYg6AxLplF/O9WSk4WzUNFwkf36
iOIHx76sF7AXSutRqfKDhFtRtz7Vq/H+kBejWJI00g+dbVj/6q/HVMNPuShxYMeTTHdFJ/o5mCzS
ojHDJXAFYLPePhpWKZTzs3MBIvxU2JLRZMOnukYq7BmPVoRrmyScHluLONkV0zTz5nZTgWNjS3Lh
YxfI+uBbMSBXMpw+fOpHN+D+ulKkRadaiH1DCORC711m0GLpXdWo6t2Jvsnz4aVKkoSjtGDZ1o+g
BzpCTKjrm1hmmECMiJf0D30htEAcmcovSa9IupATpupKsy+TIxvEAXl9dn5gdUiSP2R83EFNwOKw
aoiJgxz7e65NOPl4FJIVLjtBjlSFMtT3MU9a7KXC10Riav5peJJd8e0XoJsRDJL9K1vEZOiMGnwT
miyPFJpT2FGgcz+TzJO2+XQw2aGGvjgm6P+7AUgjDO11i2UFTSZx1OxvXvXLzKArJJjElUvidgxA
U0z97juJ9LsBKsLuCgHmMGwx9gviPVTqGq53x45zTzqBSGGPTwg03N9OBbwy0KU55+cvMrTXY5lU
tkAKFpAcLmOR91eZJNiNmn7CMSKujxUfykRfHrollNGIj3KkcoHDmT2+pTUTv8KdTX3keWpvftrp
5LlrF4BEn3gA08F7HNn8yZf/e/XEGqUN3HYe3QSdkAPZ6S2EFMM/qib/h/aDu0RFb5M13dEFiaYJ
hMytpFbZPROBeQAAPiThS3EQTaWYveMX1rWQ5C5yWtKKZ7lPLU2i19fhaE18zUAXeY3H0I9Q6Dly
p/npyczOXy7apIBSZCWyLcBHH5QaCdMnMIRBKjV5PBm3hN1oO9y5SghmtUzchn3T7xIs9eQqxSRt
XbwQTypxcsKCB9O9/ORDub62skSbmI3FmmD2ndWWCb2bm6cWUtDpQJYPIdHnO4kLI4oOaFt3qVPo
UrvwFZ1BR695sGEs8w+4VmqesoEjmYqwsi9U5TF+LYNhcqpcTxZv7un37n1SZRI4nmFdo5TxiHZP
RgpVAkLxXdYoLNU8C9TGCGKnbxePRTrK6SlhxBwc9edIhhdB9x3IivoFbpg9anPBq5l12o2DatMq
GtHMdRMuQbRAUi/7V4Br8INNKWT+YMzPneNTs7n8xkk+cwEmjwy4+eVkPzzx1Fgu+VCpj2S/+zps
qYTGx5rNoZBdpo3E5nO+6SuQlr0hbCiVe/vlFkZrbgFPfkMzuLRXkqByaCLBQuGxoGOzWvwXUL3j
htylLmcjW3ndOX4ZNuwehhfQkO7RcCuSrduWKfpJQKB0VYjEvlyajPTXI1rGk2gNpog8A1AF94Ec
H+UNjUHMLoR54Go8Ba+vdCVAnHKrAiBsUdu4IKkzMUNYIVgRVmTKElIvWP2C9qUDbB9MXc4ET5ig
Fvu3ye+aa+tXS+gpp3YQ3p326SMmxkIyIpDmhMHZ+pytBhOfn+9vMKKKF6jdETNyQyXfV1hWlURV
6z2LjOnodPGA/L+uVUKUIAONBvaYPPuC9GheDB6CMzdgwJ1EVjuTOz0pTJbZvV2ZBsiOdVdbXTvS
/K6n/+NAkPkNMcSCKD792wiVhIfMmaVc666TxRV/vdqzJlzpSQTrEC4MwfwLa8Y62ZAwIwBn50xs
bU0kPzAM4+C+Y5HT1McYsTI6RlyNC4WiPo2jSrhZ0kcYMUZbr0zWHPmSLovIJJVPyQEPtuO0VsU8
wVfFuDGLJkiq8TsuqPLAafwLLLQMxryuyWGcamulUoD81I7CUz2J/FrIGoe0TeRxT5+9WxMqp2Lp
BuCi6buYQwiJ5NuyWGA8Pl72GzRo26Ge4mTlFuihFkQvbtk+qWxYEIIwHWtEmAwd/i+HleRNpyFj
S1vXoXZSbb3KFZ+eUyj13uODkF3F0yBK/k5lFXyQAmo3dWYQTAC7EfdFGH1xwlbtzX6wMJOaX7uF
0ZumGFXWND330q4r4/BMhTZGXAxcWd/RxSCPejaCdA7Ss7vMYODTYYLF+wwmWRDjQvZpo77YdBt5
8VxzMiahqeYNhOlaHxvRUnsfwLCUsT30UNaGo6qdUse/yhEuRyYOevcpfcN7TzAlRSC3tGufgOvd
9BOOQqd5agMMgsI7Nmym93A0QxdEad81JOGM7IyoKIobYJDeOldDqa/4z8Jy9Kl6PGbAfyiGpXHE
i7lPT7Xfo+k4go4SxlDz70Sl+uz0XBGaK+DICyDY7FoWbfNW+Ht0kHebDSjqqoxoBzFhuk+IyioM
wXV3EwBC6t6bHUiol0ZpZSbknWvOszRQze4BGovJESsPN+31/Cq5yNvqR8pHQdMuue2QjEpdR5jZ
1ROy47lgUVis9LPvcrPTEhfAanbuA4fyGLPJkKG3UhwwRJ5CK92RE5PPQ3BoE6rnGEmh+HpaFhsA
jv568Iz4DSIfYp03KmL3LH7Q3O8QCxcyz+HuvUpDvbvqseijXQuRTkDSlP7zClmWHFYUZ4qq49iI
GxGqmQ/6lJQylUsOqzls0wIbdkoasjhdNC3lbFJ+r99QS6KTACReELbEbZYrATzBe3qmTOZMt6fK
Au2LwMiIS4bWG/koHAhVM/t3whtzSWiGBxT1weVPxUYeqwfO85Nq1f7IqoNn1PWhkPkYiVaGy/eb
afwDAnB48DFMCBPL80DQkJCHn96zqkNEUbTWNxiEwQlZQl4deiAjtwxS3+b4fn3VKxSJU3HUGKB/
oRCpjjefQghjX7LER+gbzGgA0ksKCrsDxUUYLJs9heC07mR+VKlh7pOSAHqjMJVV5iQNgJ3P7saC
rKtB+cb/+44GO+vGtDB3qs0Xc3PDJXMYnzZc169OttQTxhWlmTXHpP2NnYMd8v18WkjNJ0BgPeef
Prp3IZ++lm2SwCl0+pBykzdrip6cS5NGoc00Xf1rYcAvrnS+HhuanlAbWD38caeyV5hJaVi8RUGX
9TY9wJTGwBmJ1wDXFqE650ZYGhe7j0nytksCagP4oAs2uGXwURpxv3pHazxl9TIiq7tQPVWjyYXe
KcBv5ipJi8CkAP6iiQOxpxNrTMKOOko8rkvbOOlXXZzBV9V42G3HCRSn3DNVqEQYJSMxnqbiwNcy
yZI+Ot9ELUqUPx3Fn0ZwQFFUjwMEi8lWBzU7vguucSMQ3AsrHYSAp4nThcm6sqc07rlLHUgbv6ZE
jV8m1fSUcmq3OsUqrRFCihcs9R4bidNoDkEYwaareY5SZnwMKmMajYX8hwAgePxQQr/9GVotoI1d
ZAeAcYlvGdUi1CFa19/+LcFF0Ui9Cybqmio+J38nwicLbCiZHe6a1fdFYQpSPiZ/mlzpx+9YlwF6
RX6KJ5UMfs/24eoPxMUT1nErAPFVT5+E3ans1n4zUpULg+suJ5U6SOWesOYI5FpIJcdKHCIzvES5
ZcCgZuuYcDmjZM2PcYtROduhFzcn/sydLIwG9Iw/csje9nqLTRCN6ekESSHF7JbMkLtx5Q4sWblD
3SjzmmgSypnpr+oApNIFFA8wEWLzIVN5/DbxXAbiapn9ca3mh9UHjICYsQUc8KgtS7bQiPnym2bf
CsJ7MX0lPz9IP9ZFp1m/SuZkbYah2kofWfyf2YZVQ8ua+QI97uawpPCaCrjP6/I2ckwnE3IC+pTb
IyLt2/bH2FcmNYKitVMOcxcvYLYQE8rbdBI6eS9vjkZ/oOQN3DuNAUf8bOYMepYxQNldp4KDES+t
Rj373FAzDZZGzeeqDAr0uSBcWrsyGsxWmPKnrGXTCSCgl1+YxwRXc/Hd4514UJMNAceV3iffIHLj
TfUSEEqCf6ewMaM4zSwbpbjEKPs1ecQxCEbGIF2aIq7MoH7Xtzs3znIADWWhgw7w5FFKRhD7YOOU
Xx+pYP4yv1aUYwH9gGcMEL/djlQA3WpFzh9ESoSNUuIhQ1Iy01OEr9hheiNC+7vgrvOdNFAfADDc
x49auSFXTxKJXdBWtklLbt8kBXwbGHgBwcDilYoMPGD1Mey67QCubsu+G9o9TzmaJe7Hdr7/aM6W
g7bhi97X6WMI03ozIFso9tPAcr6ElVYZQU3rM6Dn4j8v4/jEYPGzECDv/G8JySdh4XAaVa5FMd2B
ETT1vmCHWKXD3crQfDPARLbA4vXWo/AOd627J5oCxEW8kIYgSSD4gicPwQAW97PYtUNtYflPwks9
ii4ueWx72MlA4NOdZvwopDuKICQJPeshhVvoa87lO+YvHgc3p6/tJgKC6590xODsNi/eWrbbh8hw
Hxl0qSWuRQ5GfhlpaWk9uenDalYQGzt+VXuybNMBIGt0mosLe3Hd+Q08mZQ19E5OMyw32zGQxleN
zdHyqQldS8S4mmiZzTZyNug+vAFQLBpuAtrIYasujz8WmXrObagPGbGjXNRPc6eQXjfENVOWhMS6
g/5rkQ4yxfpou7OBGy+zG24iVLNUZSixMepdnI+oheCbL9dEezW6uNd9rxe9zVc1uAybgIB+jJGQ
S+jvIOkzCnWbLYwQEWL5vaY3ijHMqnFRDFJ4OPbERtMHnMqkkxFZwmKvy622uCJZ79DntK4Vz2DE
jxMFMggZDMhD0xvEkQo8j0gxr5v8xvEmw1h3cZ8Vevm8AEo2AsFwEZwlcULzA3jyldD9cgVZSJdX
iaznWTGiV3LdzAG2PgVTXMg0DT0g446bQnK72KATSt5VxRkrUPzhEKCEl0wW8dEz//R4kOjiC3Xu
bAkLxqvfTx7CP9C9taC86j4jN97zRHUqph2Twx9C74RwFVyjj7n4y6nY11ej4CyP3+CEMkrJV/hm
higBYfH/88p/JDLCTPaJuLwW7fnXOM810WZHA9gDJDCkAnKsum6mdruYmFG+s1/ZMslfIczOx/iN
1ohgG4rJ5HSh5d4zaLagqZoVaKqhk0SItX15qKzVsrnVq7QbOor1YpZXJPhP++PLPVV9KFrx8g9A
lNpbazmGayzBD1mdC8hyDFn1lQqiic7NKKMoOIwegczo5HA/fiMHrnts4t4UjfV7yIQ3A+mg0abP
BfrEFgQIIeHmQ5qYFNk3nVnkxtLJoAO3E270UOvrV172rh0AaJNkLw5PmeGCsJBT+lyoGELINMYO
SVwIXjjHuwL9gOYg8WdCu/lgSk6LTg30XL90TMfpjhdgZNAZsNoci0ASTK++jZMP13gnSfvb1eZr
HTIgb/xjJWDj4WpoxHA6JPbE4gA4OwsQeH3avgybz/Y1avNgQ337jQpc78BuJwZnGpKfW/ne76Mp
c6ZH4TNsHpkLWfHlmNj7//hZEbsA1/6dnt5w6eL0u31oXWg+GTyR62RFSP3mx2UKnNq6tQTA+bT8
SmhLBeqtAKzUC8+YRuFnjl2q5pSMagjg2eAzrEjbbkfOLSNmEzzvkVwV9w2ac2uLhF9vYFFIBhhd
6jaMjsIWQFBNKPEVwdOoUfjRX9CnpuZbWTc28XdiWPl5foWs+43pFE7BHqYa68/hfBEzApOBBtsZ
SpdGsYFwHjbHdPCnIYaWeVECroHJNh8b/iqTCHvu/zuVZ6XBAwMr0mFs6z1t27YaBjOd0Qx2HMG8
/ysn66FR/7LPwUx5zBTHuOIe2Bkqw/LKnFGkf+fhnCrZI91321vOo2QWrVGz7y41NiSvB2NpBbGp
WFVW0XbuMamURSSVUTIWwrnWZ1C7hDG1aeyhCnuxlpjDG4yCaJlJkDdKsXPnngEgCOyGJFmaaF+Q
e2gEQA3dH/99N75Y18+bOiHxuZ7VTG6NUx75Lf/CoJe5dw/zDliUyczxqnXm2iqXDbe/Ia7sW22E
KwQSYB93rORO5h2NfIWihAAjh4oSuzLfCxr8RReT3owOc4O2+DAhDM2Z1qJ8fKWgSJQdoAar8xbE
eP9h+vyv9gvuHGxBmUVP5G1Y6d2RGf/RBQheYgaCtc2F0uoluBcyX6BXkS2oELs+rh4+LGhIcwFT
wZAhjhGSrxtgYzr8cFMA/h+tTjqBFjNJPE3hpUkram8P1O4QVLLsdwE1O1+ONbphkJftvH6+kRHn
04TjUfF4Kk99oS112m8RSnIR2qM3996KLGPpIIS5iKyw15uxusPhTTLwk0QHqIjP4Dskm/pHmL4Q
J0VPEJwGoQfhFOIdQPw3p8PqsQqXeqHNAJ9D/Ts+kAcQ94rDSuohqfRzX7nSSGZQQwf1ovS96mDq
mpxKQrFyLErKztP+Ui/okxpRSzxTN6syuKzAl+l6XrLAXf1p4u0jaPbcMFlHqlva27ekQhdo1Q/3
0dE4DCvvRzQao+2pHdZ/+xPlDmcOn4zLCtOA4W6xGgI1DtDVETA5Db8Lv+9fFgF/EeLV09+3n7k1
QufHGqV87q74uwiOIPgp8WfyzRc+Sdzx2oCOJoeWBqIetIjuRL9ROYy8k9podiwyCdWYrtb+uiLG
MqXLYTuSu4eFuiWMrKwg2bhvMJUpb9MYsDefxjSsKEnkbiGO7JCghydYP0iNjFhhMRugup/LUwSN
stL7o7UNd12jzNJnZdLlzaU1rbHLNqJW+cBY84HlVNWACpeJhjOKeo/ZO2fIErc5L8+m/ElcYE2P
7IY5NHKH0A740OQZyX4dlwuMb5FFaU/YtJdYvmsgAq8ugPxfEhDHFmWCgjQEG9y+ncLQHtDuEV5p
k1l4BveDTQrY8917wqJw2B7zZYCii7ZGPXt3C5WZrog0f+9846uDPVR1IUSsbTtRb1sArYNCasq9
UpoJ9yr4+lHYBaQGRVKlN5UU8ejHJCSugYxzS6X5PxAWnqys92vaIMTKnCN4q/bz5mrYfOCYBmf5
nttCiJwLpIAnhDLRAYBzlzYO+jxlghW28YWsaXbI+vrh7BPHfu2n3bS+XCA4mWL5a4+mRqX1Hc7z
oey8f3GguDJ4PWoCxtXfq021NCxWVl/4UVLM0eUDngFc3zuMnOvMQbJLBSrGLJu9sjZv7tkLz7Ri
+UT3nM7qq8uTbEDxpxT5lCMyDd488Ix1PQ4+i9sFGQuul85xQTpyJu5UfsO894lTrYQGPyliYOhC
S47o2afAvcj6roVSnn1vUguHUvMlAJaV6ThWzYa4jIXqLPQ2WnX+UyGv9wpi7lA8GbZy6fUM04vP
FRahTsY2ENcaI7gbXmZO9siTXdKOvIn6I4OD2lnXRjGE0RHKmO2RgpzfiNTKcxXuG9ZcnPqFUln7
dz995GGf9ioK480I2aEw22Vx8yVEyp7PVn4QkREFIjzkRHMjUrblsi6PZWe4xVF6iyGLoyedvbOB
wqlRdZsZIQCK9vr1DER0+y9Zr8PGAJTZpNxiJ5cwqUHlj1WupuMTNYphSaDxIeSNk5vQwmtjHI0y
Zt6B4/2b0zh6XGJoJ3C4DLJF9RGZzXLpNOapOkMGGx5YwoIxkIG74EWdpG1q0ZuX36VhDXznC/EM
RWEGQvaDcLvD8/KVKmouGkB4JMlNq1nWOW9bKXhFUldpqzPySHTnoW08f71RFYNdDaAFsm2UjnNK
dtSRnHtdl9HvKuI2qZ96D5g15BAbIx1cN8zxugK5NE7cuCKCOH/lHNCgW86kEu6o3GWM05b+XNov
j4mRo9Dx2H1l2A2iMNjfWuGFYLwZCpViFKai5m+U9pDgHO9Jx2LT+EdOe60gco9KXDMmxs3GNa6j
qOKaKMWLDC6jzZn5kaXBC/dHKueyRuHtl8H2RrUHLxDtLdDmhWZNjwnollE69Dy7N06+stOFgqKC
xE8xykA4EEIye1/DqRfL05KusAgpcunFEFKpJrag/rVpnNEYxP70GwvuqZsIZFVdTWvmFa7XdWkI
FR6+KH3KwQLnN/KNtzhnEjTJFUlr2pkt2PnMXaNqvlbVDkZx6ScXkw/do72C9Zs2rBfn5gN0LYN6
9QtkXX4zDpVq/wZM1daRc+o1aPNFSdv+762dq+gd+QNK4gQQupPfLcOM46YE/2H3IqbHj8PEs5bd
Q0z8wNXgo5u4AE639gyEC57w7GTbgEKEG8psN1OazAaHNA+GhyodhkW/aehyyKu4s87wezCIAOet
VyrKAVuYAnhV2oXS8tKPtl/zMPq0Sw77BbpWu3/51jqWYggrju/xgv1pSZwqPsDSYoE5SR56+fvs
/aUdlKBLcKV/NobpqD/hMG05Cu3852AjdFzR9Uq+29rC/4SVUFEM3+sIF53FT6TV/D2vfBPijG4y
6bFoPFmV+J5f0qidqxF63Iob2g56FyN9jqAPGwJNByPB0XR3s0FbttTvdkJ5ILHoWV4AvFhCqj5Q
s12uztAyVzEnJ75SJwZudynM+/8xtZDV+yk8iaKw4/1ymkBGivFO+xwe4xJ9dh2h5JuhHWGRlgUI
z7AHkHCVouqwRkc+/e4O8dELbX9D3ct+kIXJAWCiz56zJawBmO6txYMi6/FPGjsziXTSeRrFIA7Q
2s6dk0tx6hkIpdJmcdpapWyl5MhK/9QWk4SpXiUluP2zx2kq7HKaS7Tu/qLcqGXes8vibgwg7Jy8
8qwv6Xwkk7GSQMSIhzZ+TXDCw3vBzs3YizzYqgbluCmGdhkjSOHofZyNE4Z7wLGMTmC5+sl9ZCiu
l7K/rev1ft4yDBHHvGEjZx1va/fxtPqTxrsJESqHWtPs15Scl8ioQOZdRz0DMIW4NHU6A6C072Ls
Z+W83HEufSCAK1OfYbG8p+su8Dt9raZlMaVqOlyvH9lMybLExPPGjId+74A7n7QDlmPPLBJjamyN
XZoVBbf4UPqF0GMxgpIrC8t7f7PrqIjxs7Ly/T6lfdQFjq6yFnuj1QSApqb123BH/vyjZvV3tlLd
S9GCrjfXVrtyxPiXJ23updtJOm8vbxKEyzIHvUG9+/yVwAznWmrpVLdyY4v1+MzfnFiOVFedv/qA
gqv1uHMYlR69+1Hw5cHUvfBtVDekNrb4h75oeDon2DDxVHdiCxhFig8XwQoCtpPyDUStwsd8Jqmn
wpfYF0DY5GgrcWs7meAxEPru4QT6h8zhcfPK6z4k6RrzJUyS8UvCUOzq/LzlmWj8XyozBntNTrHE
XC8MvMrSoEcujS1eXP9oLOMeTVSyKVz2bsgBmx5ebfdUj3kobqW3wbmm7baW4oheTNwhHBSV6qG3
t7Ycd3rlZ2uV9r3irEvOYcOUnUurfJX2wxvS8fWBHEnQyMgEHzmP/wLhRWWOvIJbn4ffXNo+cFQD
UL2zmHdxI/VxFAcNbQtL7SJXbyZib4vdvur0ZhwVAzAIkpLynAeKhjwMn5wiRXoDulMQK8NFCeib
5FPaH4excZvN5FABpvGV3oIjNeS4qljpukmVrHrtP1SWL8F5tiPpggnLJ5S5zSIErluK0UeufeAK
Zfmda28/17IpNoB+xReFflI7n+vA/Y3CU3InInSSjizW+EN53caUV2GrxwQKSd92IRyxHjwoWjuE
3fr3V27IYaxygowsQDDd2vKjqlVKbGahifcvs3Dr9I5XcLK/NcWlij1eUehELo9BajQq5FKrFRrs
NjxiLzuqtVoo9lcxVqPEhF/q0x67ijzMZPdahdPTbWv+0kGDGaFEtS32Bamyf3CZNnKWNghFom9l
nFz/rVHLvX1cxX/dhzDXWhLfHmcMpU4JvmvIz6UnGupizyUoRNcKAyWtZOvuJtx89KpZDelwPwbB
FzbNRdIOA1IRci08Xe1AlSwryLzboBg1uBl2ssXw8dZYLHokfTfGJO1fUNLEdUfpcCYfoh9ue2Nm
HRonIFsYOw4P9wo/Ouxhi98qmVtDhd05H3S+RiusDQhzmT8Y7yISnh8uVwXgWhSpXsv8YYuGNaBu
gbEJTWxgULBXinaS8UePiR91ATgOUTWtfLHUj0e8kHjTtVt40u1Aoo0NtTMSuycAhwN/NbkgR5Na
cQMLnnolnjKjKXlbGwwkf7AIJImm3MdlD09ekQ4FADRuJdc4CR8vdayXueMFZskQuXd1/H7nTH1A
SWa4uNQoSYdhjqh8tcw4KPBMwN9KK8BPHXODCWJEoIcL+fCbhfw/uvF+0YKDrZ4g2hGAh3g10TRf
Oi3YYaA1Fto91KiTIncbttw3U+5EPlNoyuvKcoKgtX+CpZ0NsL+OX5t4FWV7d4QPCJcDG6gc0Vsx
HNRTzbwkqZ5qjx7aUFfKWmpM1DKW09psANiXdNDXMQBof20S2YhKTRpFLrB7Uvufv+N/OENnD5kk
4RjGp2QLM5KMs/ApWpoviC+dxGcCoirla3jsL1WjiJIh1uBsSyzGpoqsBGXg1Wakag440AKhisvN
B+84I2SbjuR7IxKRHTuIdIGj1HhO49Tymt2Ip1MKuhV7TKmGT+aUeD7uX51K7UP0LOx0i90ViBBT
Dptqtu0mxJn4Mi9ZdWS2kU9fYOX663DgVs4YjU9Ah3zJb6146+i53JhCI5S2LE3GMu17nbDOa9nm
BKY6L47pqatbR/qMiVCDwcV9anm7dmu2PbBs2nT7MoM4UWNMmPneli0cKumnRpPVKe9pdqIQo6zV
vxM23+LD4w20eb5A8/SlV3BI+sQ7Ib8chUA0GEBGYKNMv9xb3KQv5c8XMSbjJNFKmIk2gwTo3UVF
7yZI4+iG91Z+zW+ei4DDf8JVu6cHy3+57V3wRSm7Z9GsSL+vqicKbyHGuAcAIy+78JuuIp/nHjBU
jVH5g3bbzZPBBYKcgMopXgdz9VHGzfnhplr+O6Dy3emMq5FC3Pl/Z+oi6OACWSgTcBPmRxSdhfvk
CnMyRBiQ8sjAdeWLYGmpIyikWLfcam2tFxdzJFukiZigj8FhvlULqbDO65hlSOsvaFXApq10VX4Q
S2UT7TtI1igmpxTNJpb921dgkvF6YnoX7NJq4wKR19NCzIc11N7956/mitD5GHBS+8k1lZU5fLLW
PMUDQX3sMNOQwja8MY2CdYIjYIj14rKOfQiCwlW8jQU0EiM5qtrqDC8gL1jCrV7mZ/g25bJZNjf/
thHeBW2DERqAG07W2TnqV0fxVjE/WWrMipsRDNburMitj35vYWveuQLNvmKc+MDutEJ25cgQLarK
aYjMXoFRQ9Zvf8603XPcOfeGXiyIVdkH9iPlFnxB46KUylWyPXP4RW8IXj3z0a/j5Zn/y+A032ha
5h+iFBH2QgJ4hGjOq//xd6hcBfPXouPWAwcy49cYF+OUjYi0JJ4h0Vcm3w1freoDpJRmFhhis9Qw
BrjOzhPYaoAXw1La3mkEYG9qU25DP7p+G2fYa3/dKTAqQMTY43icPmFMvd7l2RftWjB//mOvxALc
sHlZ7yURLstVGsJnO+N+/IQ8G5mw3TkpY9TcDLdPF+HYyLB/AF05ka1iJIt3z421JvBw1pbGqrDl
4dv5sSO4ZFVQ4h8mRQaf+sqZKB7o5rsZ0xBOBR3UwAX2zPqwUTxb8q7Z8LJncJvef2CAusd5pCcN
6fWRrRKBeCR3B4lvGxHv8TaH268/aNjdyqEDVfptZgvuv7VYx6AVGnsBpGv7ZJi9Je0i16BjXO/0
zFaoE0TCGokANw0cp5DJTCoPEw9GQp2lRAj0Vc+xFTlQDO94YzS1q2mzvQT8mNM7GJxgjKGD9Zl7
oQxik+M+HYHop0GSEOpGFWlAzDpG154SeWNj0crcWzm3FjVIl0G9nsc7voeHNdkhh3VmM33P6Bjx
KuhkFbwA9rzXejAtRB2oj1wlO38IR56xtyw9F5XlhGLZFZwhgz8f5m/Kdq3xUv+OlhvRmkyu3JAV
mDnSMATVwksjN38Tm9R0lIjZzlB7s0jpjw65n+ykFc8pssiqWs5PoMU7PO7RvIJNjKdwpkW8rPIj
n9B1X66GA/UF/MPv9YrsvjNR8lOX7Y7pCMgwvkNUn1O/x+1WPwEGAl5+vBnpfhiOa8pwL9TS4hNs
UUjmVo1/aUWMUMFOIn9Q5xbjVhz9qlJ4WKOMnkXyfspHiwaMcTnbcAxKOYayQ2ZrEDKTC08oqS2r
qzGzvRceFO1pihYUfTCpKaz2hys6mGNtkfU/BGy8MYKlN/ruPHKkJdVorxA4qOsWcXHKjkfCSLou
E1A65aw2RR5hg9y2owsKnuCpsUiNeq+FQgkEozMb3k5jMCqrGttx8R9ucyIQ+b2a856/bSpBjq3r
8HoKg0InuU6B513KNB1a1+tBhTzA0I2p+9vDW3HJBE9PFk1ypqg4wIVU3MQLruV/JeZhjB/MllvU
vbDRA81WiY9NY6YbCuOlUIqfrYVSlS/lAvHILsy8xn7Qnw7Te7YnH1HY68kUtbirwQEi5JUu1jqv
wlD9BZugTwH9wKJki2AOyRBYKidhNwVZUPzVlctss5togh8K1chNZhcnyLxlYiLgqZKmgwxwrgrQ
2emuVAY3EA+IQ0cOMuLeKk0+yp/XL/WiXChvkHxPyS9ol97rQqc9nD0PQif3a9DNVk2XtIZs0iCo
6fzwpuyZq19vcSGFfWM7sfcNxs4nb04o5wv4D6HbM/4hX5mZZQNoNikD1tySNUJBJwAxcXlD5bij
QuBuQ4zO/3NG3Fhd+2IZIp+YFvsZkW8+UH+TmwfFN/SIZXrFtJzydBUnYtwuKnnvB4h4+Be3vyu+
z8Mc81lCWvrewaIDTalNkxW6xQqqKNQHlikkgQGm37pC6c1ZvsvIe90MDDSA9GQqwxAL0pE0OArL
+muWprBkSb/noaR4B4Hb84AGGxN4UtGbY9OvANHQIowYjdqoBV7IsZ5KmZOJNqgywBtCNbam8cQt
koyna9sC54gnJv6wrILvdbxN8brDlivfIMq1JUU3wXEBq1trc4UTJCduQYzpcHNyIishfRY5OOIH
mrL/IkuZxo6r2aF3p37xtNkGjlcD0WubG/+bxep6yuwFwEfK8v5eCv3773IiiNIC9voZrefNkCQE
0Cg2Z7jL5uuTctkBGSRg4Yi0aSa5YQydAq21PkOVZ4kI4oKrTzvF+c8KUBYNqHag5voRPq2bkyWy
XBKCZBFGj6H9Kk+qx2WxuJDfESu4BV0c6IPkcLaoKlbWhIoCFL2l4BpwdJAVV+v8sq+y9cc402Cp
29Mln+7wLV5ARn0oIwWiaPxDoMGjof8YiccwuHy+lL98Fq2D4XUsDFRdrXJ7wwRNq1SBtOWenTXu
xR3z8Q23fJjR/9yDb2Gu5+vhCIZIHTRU5jcVhNNQcLtqePqbTSJ2ya79t3iBGIIkm6FqYPXdULj0
SmdP+adKWPyUHp0Echm1vBTIPx/CDaXr7PYsvt+JAoWumDQdiINeyHopWSmSNYViKrf3z38F2qo2
dzfQ9wRyQTaFJbYNJYpaniQDFD8IEpYuNp8FvuGpXJ39hKECs+2CtgzcuLkE4NM/8l7aW2yi+oe5
+FNLpitECQmOMgURnHbtjCJCE1EN61CmZfLlVdGIu8X+bSu24UVcYekFUzsTMn6Nk6/SaT4vnJQu
tEcdwyqUnVm32mwg25Nx80lHyoBHlWZqXx4OEhcjCF2aCP7Klz9ApFbSRIHwHuYMVetrga5w9ZbD
w+6qffVAXqt/FdEY+3dXZ8FS9QhpUc5AGLLEu8F2l+DeNbqsD7jBT0dTKHBcZVd5DCru87iU+4zZ
SZf4/TXOrV/gwNRVjIkZbA+SNKOnEoQViXWl/4/bG7PhK1ZT0IYY8hemgj5vErt8IZq8Bly6y+Fs
5L5XH1qItTz4m2gzmY5Nnh9gJXVn+qXgWune14zFpEeD/0p9L2sPmiRqDDazJbaCD6MqYtiPEv6k
+DyGXN+QdYkzvm77wDAryN0dh0IJQ67O1Ed43Jw0gdoDdmbHhZKjRs1VOHbM/7jEBMrGxVeKOb4z
mWR8dtseSINT6leo2FIlzYbnz6uz9I8W56kKQeOxNoDOjZdkqftMH9mpxIx5BqKsJbavr1aziIE6
w+CEOBAdh42J3DyjdwtXrqtliPVGYoMrqzEVpi2BWTdfv2CcR8PE6DtxZ71h8Xrp/0H5yD3zSqQd
lst1mojEP71kd3Or9O/a4SD/bJDnmosEFPDcwybON3T5T7Uxq6VOnZUTY9di3CEz5mtI0XFOq1/h
D0PXt2+0Cnuf6qLTa5FoGjXujI2K1pKE7q/0inXWPWqxBb7qGBnGvXvG9l9pAsKhDMcKx72ZJBkL
x0jwxBBkyqVH/ittgXH9PC62qp5IImctRCARbQ+kfCXX4QYq5fa+k9RQkeqUhIBxVTEHdmBy5TbH
COEVUvzW2bDmY3rZ6yr6JdGaVCgd06Xhg8PuSWK10165O0e57PMJKFioClDKADO7qPopscQYFlK8
A4fR/rObu67001WGtHx9z7NNJMelDWX+mt4cbQcg277IOupH6lxMq/jvwdXKHqXlj20P6yp50Hel
E73aQe2vWkIt/4aKjU85J9GfsbQnLEMJsTd4dOoJd0aerri8nZsMjNi5XDFRxG/eCM/NL3yJuU8J
N2e3kqtCubrKaVbIbUW+1/paUGCO+U62oO8kmnjd25781W1K0gdleoWwDURKNAeR2Jf8nuQC+vOr
C9zBIv/qVBfS0JCdo/uV8vRsquq8gdYpvd7N6Hf6TAJpOP8IboFKPxbW7iQfDv7cDsRkFDuOAGQW
3g3kYerDQQBfo6Q9nhPau5LHS6eAEb8ZcK5+al5u+ddZEbZI6NkPBQ5EqyT3jaqTp5MCT3eTk6iL
Bw4AWfLb1oMqQcYydBJtpLGDrGtNUn48nGPdJz2uv8LbQNQtUkqs6tI6/Uyja9XNpsDskd+AUs7N
cWPYTVy7sF0PyGkie1+V5fqD5gA0qHMLnWdq4YHYzcCreAee3Eg6gEY/jS6C6FhukZcbSfHXMNNt
MWyiblpm82Te8F/8llsao+Vn14a2NTkXMC58zG2MEsfn9hSIzy3lKbZFqU2tNIO0WVxXocCeI1SH
1tQyK47PwrtWoPG+6xI9fMRUjHYBShiAeJsEMR4jGcu6HxTZI2xQeQuzm+dkFtm3diBpkch9Skpk
6ebKNamlj7uDdjuJw1fva8Rts9KSzPmxPRnWfayeQey/Qp9/X/swBJXdSaFtbCitAIItP1dvOeNT
EH0mxK9lln7n9BeWHYUPqHs+zjiYz/WftT+T55lshpR6IZUueEhpSnOA7CZzbYN9J4R49V/MIvvj
W6QVCQ2JKRIvou2Vusl8ZaswN1QSzglksITC9YloTNSQsPTAwfhDn9n9VOSkACtgTJD/3/weioKo
zVaB1ElPCB5JSyLBRAhe+3jXcLq+MeywTpCj2kcKOSRciQjs8cFzIutVDdNa/MRROZh4bF5yLa6M
YfSSw4bdj+4A+/YfMLCg8s8qgSV/4U/FaADQHWo8nRmp9snZ6jfjU7q2/t5x/khI880+FafdCvgz
uEXTCMvSqlcdLJxTnUQHOPJ/SPejadqNdK6tx9LeV+yjRPo0//wqdCZBC9b9xfww53E5xfckstnW
DNaZavSMXtw8J6Hltrxh8xQaet1QX7fQc+MR4pMDaDtYl07Nkm7ck/wgHJJ9M3SrWf1O1dY4KYiL
riVLSCneHCGo85voSjhxP8ZBQACrmYT5ct6yCXhr1pCmGXRKptilRdhm4ep1DzU3ggUGFmg55RY7
q4TOL13IHcfzqu8gRhBGyLX/xEsHPFyhUbdr+OWTIoLy0+ykcRJADeBMZ8xV4iXDHXkXLFKq1SeR
TuVh2ZxgW35UOPQJIWE7oRKXaDGLMRDCDdpzziEx5C9lxet2zm2tqm4wOAj99DiP21tOl7iI3dET
DZAst5lXCezy9ePsY3J7I4+0iaqeIA6YsHUJPWt+HGVo7g342VI4ka++x1HYJ54G6xnoggcBVLQF
9SkvNKuCGVgxP3Gv6g53MdeF/LMIJ4Vm4V34cdpfDzvUxxqRZsjLt/BnQ9rpcHR9GeyXQWi0Q3Z9
/h9nXjeivKDb/RCirXI12qkdl+Rj4mlAAXvvV0GP3rqWjVQPCCNrAarH7aBvifDkPN5end7Ff60J
ejNESxzc4EAuh/vmFMH1Dpe+hALQb2IWD6vcBftVvilgzy165+c+LaG6UtsyfjhfoDShwQ+1YIyQ
QZ8noDdebfjY+Zr1mqCzkVmELjr6zEcyeBscC9N7Ap4aObuMryPtL2AnE/FdYpH51VhmmZhChoLA
t61Sd/Aar7yvcqVI29Qm23CePLzgmkRCK4uEaOJnkyQXePFBbB6upecFvNLZaXlijJ1hz+F1ZHAr
2QpbzsSKmJIFByHn3fQBJ+7PieohRcGYIpYIfAcia9hJKcS14mdN7Eg2GGv6imgm5DUH409y/uVx
c/BuJ3mzVBjrhX87QwabJ4/eMiLhyOCjS52ZRYZYZ38ZhQtmCGi4f6rHcOI+/t20d+d4p0LyHwp0
lqbCGED+fTtbcHUUJhGbZifwGBXl1+9CsWvY0Tswv31GHcNs0DvcDvGFJoirjcL8QFqo2xemfyml
5twnw3rrCh3AhJjHZAxZvxmEsKb8zfC/T+o1448P5hUCks5LR5bWzttK4ijbpPxmbF1eODrRpIgE
zuHadRKNLEUJUIwi5KlHIr9SPHwKStZQDQn5lXfGFORJFNO90PRIZBmWgUiCwQOGUKdu5wOZOHYe
PhWM+GNOxVPEnQ+NSjKReE0YdUozGBn9a5SeIDYx2DrCEI6F48AkOzhNxffClzfmHUMBn0iJI9EE
492L6Wjzs6ULrC3q3Me4Bv7kBr29ZWmHcU1dUrlRksVTDkD96or9ZGuJBIECv5ubtxtUoaftGMM8
Vp6i89+5jFRQwwjbIrC2yH/ZYmq4eFVG72yUR+7QL96yXkX5+4HwNTud/6P3EMd1ZRV4JDI0G680
0AmHHxdgsIxCbq9mtOycGGEXmlAyVr7y+GWyjJmx8CqUty8YM9/sKEVKvtybSqCCcyIAN67C1S/y
N0Iy7aEM/RKp+pfLLpkl4iM+881zuOz84SCJG9BfEZzQBwWi03vzO4N0NDLRDi65LKkck3/HIUcj
5zN15pDlEFMxXJ/XnlOYHjd1kOyzRXXhCEpU1cvZn+zHRli1Je54Y/3/QOqpGfrPGyJ4gv146ydz
8469Qiqu52LCSDkfsy3HZvijbgLoX7YbMKzC/BZngjAwd2N0I72ePxcddRtABNG6CRM0zAzNG9/W
Q9tY6TSgyAoo3aAkU4cyI5+dfG5dr9z2A6SVCWYQknzhVopSEbtTDg4S0cKmLdE82aFVRNbO2LbQ
Emv/y4a18luiNY+VwdNM9ysnBmVVImFxPIRcmCFibYNWDEbBxWmSOSKSZBDD4ZDv03mkYWGRR30Z
a0OjTDYSWFUvHx8c8WmMvIgRdOLQ6btxwTfDnY+6xeC0WFIZQhP9oonoAa3s6aqYTW2aSdyIBo2a
2qdMp3Cyo/ee+JuM/QbKIF4sF16z7vhBum/iYgOfMz9MQ3PuVEAwVBuwpW1SkWjGNIARAR2YMmOZ
B00JPg8T+Jdd5Yjvca/MT8SYxIX1dKGsbt9Uwa03oBQ6Ix5PtRPI0vbP3dSgBAWmrm+Viulm+bnK
t0y0kxch/yQAFLHKuXcGTbsrkUtRFjTFlHAkNGMsO3GAHHhB0CMcE1zUCGvunCHcMl2uIYO4E9lG
xNDQqI8Oe1eLZBR5XitL3IAQkdDKwj0H7RM1pERAR3PgfMz/HfbHC37eAjNmhfVPgyoO59ddFM1U
ZsSzTVwF9RT02atgpyQg4jm5hEt5GG9Y5zMX3whWBWCWAGpHKIBikOXd9UlPWqGib9dnEhVKk8Y3
1uzJ0QcIZrC3nUE8YxvbRIaBHlaD+rMz5DyBYmV0PUWCb+krj79r/aF6NpngULdncHORhGfFEmh+
w59t/VIXs1OopzrO9d1KFxvaMXmOIb2Jke1cFs2PbByin30twIfH+/UzyqWaHNZP0GIojeD6WbVJ
KDiyFanX9m7uVlRFjoL4xCFnTJydCbwau+bNBALMZFGKCOHJRSXySwK/2IyicJM7YepHFb3b2B1U
E5/7D3ERqKdUAFPH2RfqkZrExIDJk2HoRE+IfGv7IeNgRJG/6npcrIcxKUQV3t9EQiEh2JytystI
pFukDC/JZa5BYwSJHy9CWhq52x/PZFfOa7NeTp2yZRMIV5uxQoCitQYwOtfjI78fkE9NDoyvpXFY
sw1jmhm/70oJnnao7Qz1Ol/SqhM2cco16qoyLq3qx0Fj6T8gWZEzCXeOAcsC4it9I1KNbb1OP0ny
IZFNIT34ylJFqujiPADgzTURgUNfVtgu1pSGxhLDrkF5gUndT8jqHC1GHjhgOZsmGer7d7RomqK+
wba0NPoTDJLdaMlZrLbDF1F968DqoTkDsWwq5OMbFLi76gjJ6NGQ2FGBBGUpZx7OD/JlKbPXb22f
mRulc4Rw1mFZFqV9VeT3go5l2cM3YlAlA4PX//9Sbz6ZFhDX+GkwcxyGJJLQkq+HuFcsTHLtXYnz
1G1RGHP0xe93B1f2BksUtn66N8EKHqzcXK/2u0Y7HxENMryzLlCt0i5aUoirT59K80K8kZLe6UL0
Svr2klS1kERK6PqZkLkqXASIQ3/KMEuwumNCezrj1n4Z28UpCQqM1+tX1c7C13ejBkNJzg+ILS/i
RHELFWr6FX6PIeZGhDg42C63B5YrmSuCaX0i8Ty38Fli8qLMmn6x2xcQXcQakSmzBJ3mCDyyH9OR
EU5Af2eojK8woLPLnYReot1EdQA1ydy7tE2Uzr96CvCC953TRG4Kg4bXAYBznBfA+neS6Duhdn/u
5bh1MmxM2yyeKeuGJr2dEbjcGMJL1Z79f8d5olZbe5+++yyyMSGv1c+9iAjEKdxcA2TqKxdmOsle
qmXfd0ZaTDb915UFNzNonFM9n85W/oDH8VUTr4wNKR4eWsIlP0tLjUoApRDPQ6W9vFXsCho6335f
+QdyHlDgpJWA64lEPSg79JqEDkV+S1sMWYaxPiVrf/49V02jvTJ9N7jGrl9rpxunWxt9+nMlyHQ2
ugKAjvt0DmAh8rw/n3wu8407QGo5t/Rtw+5T8EW+ZHRgqUq2371YW7lhbjpwtKK6UsE5npw0I8O8
dfwgeh8AFzBHGflDbkiRcxylza89qcp9XbmEikwVC5Fjj0wK4/FoGsxvodWIBqkjMXS21+X62so4
fmlzHqj1TZ1mS/uFiQR97Grv/Afd8pu2gYkJQQ/mB2bYoNvs1yWKxM2g7NUi4DMQEHsx/TfjQZ4V
hl8XBk0fPJoSnUsqRnByln4SsyGfMeqAzt76xghFJry1Tq5rC9RWSRjoVzq1gNZBuNURttJIPY8H
6XJHWuLoIlNvqVKnmSEI1y8mLHQ4qmdp6wgUtMOznclD3yRBWBnFbNadHBMk8BdvzmvGJNVJo8nG
dIMhqlT+Q43FmupPgO1aga5PoIS9YG2eqbqbUZ1587y3YuI5aZGBZZknjt4rzOQCq2QcchXubi78
hIpHApMzygBd5zFmAM0hRzCpJqiyZe4J6IRL5C7OGg5vw1xFBYMIVWmWxQ2vbj/vmAYUioMP6Kty
BP4NuiksrgZv6JuG3MkqJZxWLu3bFgUKGznSNop9N2RSJ+S6vr9kknUHocZcpUwMz9xlK5bfIvOb
a4GvO9j1C7lrUUGkaZ+bxdSZx3vDygY/E0UMq2inhByj0Oxl/gcXLEdIxK3Sau55+AjYKjxpRPLQ
p8kL/X069dnLC7yFUh/UYkdq2yEmhYGgdc9KUyUlq5Aeoe+4wgpyNzVATFlQXDh24iUZfx2JIbDL
MpJCyzr886bT5SiFvS/qW1JiF6FG7SL+6tJ2qTDqe/Tsxd66NSTnbLFlJrJWqqFvJIZSFZrpuiTv
piaNZmN3IHX7fyjnYG4nOJ2ezfTfHvb6EFc+kpQD4/e0wU4/+VsIk6IUT5/y5u38CzBHbVjzdmNu
KCeJniUDYM3gPS4gBOrEVxxAH7JGyX4G1CWCAd7WXFYZc5QYHs5esEL4zEPp5VY679gGow0pl+k7
ghj7X/KZIsDi8PmhqtpnRvjaU9S/ih7wsY3St9yYohzb6sjoqhErNjyRHBmUP1CoA+zqKuRtDLnO
JrbYvwb4ENDdfRkHMi9CCn6Ia23lTfk62BeVgYX0R0E4gvOzjN39sxsa0UhdG8QZ+dnyR5x4PslR
/Z+UVksa4W/wTIXEUAlHouQZ+JVDUKvsVg15PyHXzS8Yyfj0aW7uWIstp9+adi/0IVKiGAf77eMN
zjMKeiK39/AwK2wPRYHFBKKSpl+t854j70IRMjnXlRMg8xx7ZCTw2Xd/rVHbVPPyixcZSYiumzpB
J/Gsn6L4358GImN9kAopEWgLEp4jiRAQrAUMiMiSD6JkEA2UYv3C99wFNPpDoBJVD0vsv9facNhE
IEZa8a3ia0OqQhhmD3LHBZR48dl+EJ0mSKLi7S4A2xqaIxFUzVjmgbI3HSLXfUmdS1jm/LiL4lH9
3WHugkt4wj8ddmXMOV5IBL5/eoU3PKAtRA1tetzwt3ck5S1mnQAo4IzsVXoGZoVsVAHXYHHF6TEO
xLd8LCWDYG42pxH5Jq+QNvxLLow+AJSKr8OFqn0e2WyKh5CX44+B0vIYGJioE0N2DcyduabAn/a0
BLe20GbiX2AQKgBg7h+SVRaYaGvPK9pPX59oI61Ks0F0OH8dX9mXaQAeMFj0uQMCBpGXZotibdop
Uk/IqN3WzkKojqjWVAJECjIHAkkyh+G/TF1TBtUrSaHpojOG7z84+LVXiK4G+pcVRulatiARO8J+
J3Y5ibN0CTADyMVjBOt22gQBclIeQf9cybtdIsNBKAeA3kT0NlZuLv7itVIGRPdpHPC0FVPPgZM5
kzmZU38z4G4sVad43eakZZlKeVNka1z1Mq7RsaNFVa9VctwPeZS2RIxWV6b/tvEvBhc6bKzRoEOD
wO2xdtPgy2bcgFslc5he6xuWvYTLSy4voR72daaIDcLzPCept2ArxGTissx7/yrNd4dzBmtTy5BC
vqB+jFGcD11G8i2m1/HVqBBpfalrJBLIcbUEp11Y5/++HBcFTiqf40APlAQypoIUtgmf5zCEliUn
wXQeqxolKkRh5v+yWH52h6jH1IjmtRU/zlFcBd7aS7/iqJSIBwU4Z6zrn2WCPxLO/HJaae/HnPvp
4T68+yswFJPJ6HiRvEvDNWql2SgTDe+ETJRSBA7FKTng7l0uMYQWGcoGj/IT3ep8ASB+BfrKAiEk
FyfjLQpqCH5yDUOw5utOQxaMH9xr5cGkFEBmt5erWbMHBi1w7V4N+HIH9kZ5aBKs/xBSponr+v+P
jSKU+NpjCPwzezIeTRahO3h7rFskbjPLsJP7kVGBj9hLvWShD6kNU3qChCFciQSHAdyv72vOtR8q
p/aJivnbDst4oXmpZ/7hCY6RDD6CPcOMq3LeCvv3cPohhvpQg5pTy4f5Wx2q93hsn32+Xa9rFSgY
qo083s3pDpGnoyxIgbcMxGEfIBMgZjuo89AbeiK6jIBx1hRTYWS/f+mPcKqU7QPcUAloS0rD/nAe
NotSUogs8yWIQIV+E2OZnK6BHPGDy9PKsJzJ/j2qBQFuyF0JwprpH0MjP0+lE8eoHSgiUM4Dl3f+
GYI5WCjsZLls095bED+SLbkvujRhqxpE17XGsndCPdvYy1wuwr2mShsMabcM/WbOcXvzwrAx4uYG
jCs1LuHW/SoPeWpU/GkWRtp5o5oNZYTkKeAlaC8ecbNBSQQ5F5M2C6+UJpTKRFrBvE60rJAlsbXZ
W+mV5P4dKeoLDkkBXvfvwGRXPnLK1iwn5BYbwjYwI0IPQOZ08phb6WhkXKDb4k/Rrw1mR1hc4t2C
MMmKd6dSzb6Hpuc9uEYff7tmvVU0tf3C9Z9NQnMz21/+P/w8LtyzUajPOb7FMKd9uPZjlPlLCa8J
1KPeLhhEmkfZNjdnCLA+Z+nlnoqX2PvE1BbXEaCnhd9vdb6FMn80FWzDJvqI0jaoZuWAdO0EFYge
qkGw1jQ9A2Gm8KjWt4YngVyLJh1VK84U6lPXIUL7tKo/xeXbs/txQGQ4uxrR5Hp40f6gb5DYx0X7
+20ZDZayQORepu22BoyZYVOqWeAazYOjFrpQszF5ykWXy31WxN6SuHVUs4Ky7F43Ij8bnwaRg9LL
z5sk+Dk/DpKnVdfZcKixAvu0WiO7I6sDzd9U7171lIBxz9kbPS8yDnT7izmzyGyMUbSCLq/Jhpc0
E2WZmnuUdAlkluSmlMYaxh82mYTnB4MP8rKO3vxJNGw44vtbscCK0rLvle9560Thxq7qHbaW/tS3
toSV0kL8cumV/+AWOX4GnuiyWr0+8vLMSQ2SdDq7hcuF6fZ0REy6KFANUQ+XlqNO3vyu/k905+wz
722K2ztxdEmb4GK8aam/TYbiJGBKFY2udTjba+aekMHAEre3p7sK6vNCcJ+fhDhFtjdyjBLLb40I
8Kv0pkm/iyCb9VyFUJfAuNgzNhyl0j429pufc+Tbozcf8AfAhatyGaYz8WX+0yVyG5l2r13mpnOh
JmOQLIGULB+lhJLxlGXVcs+Op6o5RTQocjKaOx52EUIcTGMb6+wKkInNAm7yv3C/BCJGHiyWRJHX
kX61CWGjF7YqG7Y7aAsUqc1kF85tyR4Qiqa1BV4OqV2T5EmTYwbZF7iFApjExXb+wlHGRIGwOobG
peofxilvxy5FlggsnoR1SWInbbTe8AUzcQWd0M7xlZZQnCi+tWu+tREl5BmQHwCT0YM3BDlJRVU2
awxugK+BE1gRdA2y9sllTZ7fOCIslusMJ3WJRyk2k1Rowvf/aC8OYnREPdiFGKl5MZHsN8T2s0Kw
t0HNidFo6aJJxwA4ZVxaI1nsz5G8luXnYxR6aeexOTlw6hjs20Ck3NTqnYBKs3bGYolxEmxH7Kgn
lX1DN1ACc5Fdc45fG9nfE9C5bfb2l8BY2GPNj1LwX3pscKu59RmeyPqkBfbhFy/5QDRNpp+NbumP
tJhPhTjf46WiP1aAogDD4yO10YrQZIQZ3cQuHhSK4oWAdQMGNR5DbztzCQ79gCETzbEJpEaZfAF8
HiVK4tgBLJ+DFwDXWPfegrF9sHA2rumYEiWnET+OhV4dyfwbPRV4ZFvlYDHv5SyJOkEZoT/q7HxT
WDiVo1es/GQG2tTbqHtAvVaPPn7Dqbsoyda5gJe132OhKtLUkRnYVrGwxm3UnklqNK783nRcfd75
3ZieNrSs43n/nRpXuz+b3iiR82Y32cTl4hIDJ4pYhpz+Ts8r3cLKJLFuPP0lKKPOyymW7kFYTt1N
uzaJ7RXamohCReEQ/Qv1vn59CZWBbNtUdZfQuUpfxFhJSfAhJ8S1VSL6sNIaOmGgYb6eGfH+aCbC
IzcabI6zcMi70Mv5sbDXQTRMkXezSAO+EDGu9MgE8UObVE6nasTP7gjsjHsh6/gEzt9QoAHTSQlV
OTGz2hh6G3cENThvJUuKWvgfjUvi+2w0lYuA0uv8kE4d7SQGlTewb0RPJm3sw/AjzNHsjLkqVxDH
+5WU315kM+yhgRTrkPsxo2XVwX2Cr/WnZsC5B/M+mryfUylAo7l506zEUHVqTo7n7lMX67CSardW
lxyXo9ecrBTpm4sxVhO0bzvk6COYxzbtVybVtE5ZaQ/8LabKnRvrq1Jg+Y/KPW9QhInTMKP+t+ma
0YuXf33TeSieH/43NojC1ye9PUtnD9BbzcCdjzFVcQv0YMb1YxS1C3COhA5vtoXvpH5uNeAWdiKN
vVwbXcYPcbgeq8frPQW3bpPuL+zLi+3VZtVdhPu/R2AhlqVdBMvheOEKVBiLPHVMaPcKtbvE9CZu
uwIyOFKHrd0LX772sWOlLwUCx1kFM3csG4C5Qg91ijbCgFbVq6hSvzM+Qjrp70Tq7a0GUmfaudY9
O9UmPte+/3JYlSiihesCtVWMtDO2YYGCnHABw4Lv8j6LfVIhYWnBE5HUE1tEp6CZx4866Mycq+FH
2hs3jF1ScYBDctUjLR5nfh6902q/1amiq3VmJv6jLCKiSf397svRx5IaZ04wXExCUoOs6mX/E6EK
VsKKlM2onuMeuOWbbrhbXaC9jUqNhTqE4u1szDvqMtsdWx2HSvLZ4KLixlf4mQ/NRprPL8UUFsKt
UHRljHofcSy+F38thvDKkopAXoN0RSdv11Hv74fy3JNtSZiK5nbcW8ORsvkTrrdsEbcyjjq9wkvW
JBId9rI7b6PLtDNQNjraPVJ8H6uDu5qBwXSf1Rbob+UobefNhJLDeA/fcs9YOlIs/T3SIU14+RBj
kfsWI2PFuAll6Z5zRKvMmwYoD2RlDssmaAZq8vC7wAHT0/9dpbjzSRtu66Bmg+EDjy3LlVHAi1mw
qIyFsCpj3IhJ6BNPilDWKdvtG8AinODYQCqgzVd0zIdf1RvLKikaLUBfkNYfYZxXjdf+ucwXMKCo
bp3371pKzteAQde5LhrzVDy9/cUVW75VvEQWHuzhNtNUOgNmnM0bU7tdOXGLJnUHyrpkER3/bApH
5x9abIk0ukBSQX20FLNamQw8lIpLbqEt4D6zYm01arkTP8/cdnUfRKufqzrPzcacIHWfz0TgsI41
CLyZtbG73h/JGkAxvxi6PFb7lUF1+2Eci2QJBySGuaemIjhBu9kUQQFcrBg6DVtdTYk/0km3MoZU
XCf0LlXeWL05Y77R/GJzGqTabci/IsF0GZ7Lklzg5n4hZ26HQUCwYxqOxM61TdxoQRIp6hT0Eiyv
q7eAwBhS7fVYbzZuGYyswjHrsR3tmGvE1eXGAGRwNBD6oQ8RZkHKSoY4hg9/qxHAU/Vt1c+Hmq/i
M3aclVk1r3v/odsDC1a3pxj+V7SS/XYWT0abVsqIBMMBDf4AsQAr5Ts81E4htkG+AjZauNI3lK49
sjyen/3SxlRnKzHxrqRTKMgFg1Adh8zCaN678BZVJrl0ABtf6x62M28Y5mAsfXwzCq1i1kb0qWqq
arOY9y0qPhCY3M0gkEIXuvm84gU3zmawWCJYPmoxpe48zLBL/U7JDQviaBvYUUa4R9tu0/kSp2yg
HmXEkytj8bGuGNu0FhUQhAQZlCjGWOxbNL5tvqnwpYckmuSOujyFmXTGlsBIbawTz9uCkQuuNe+l
DhVjq56Y7zE5TDPT5JmczbeiAMWPf/YjXrdEyF5niAOkVzGFpKnc/UCFvVGNaEjQokQb41ahcKSN
oZ95hXtbcZkA4bpnQ8F7I3OCDiUbXMPKXtQ0WPNkwaAX8Q90oUjGy3o0sad+XaOE/QEJ9z1rtoQY
LV0fxVbwv6UFTI4+ObPYQzp9zwB3uSdAyfdg3l7DBigYsmSIu3ZoAaWwYrjUEH6KRc1fRCbzw6ed
U6YZ5EDk8F7Um9rCl4fvCBJG3LQ3+m5CvLBxzk0ZrvKqK92sO8BChQmvWvxvN2cvKKM48xBDZ2LT
v2naUhGLGG5aTCxGcGU8Tn8GWDz04hhfxdyFTo5fzGIu2Qg9rVR4LLkHFH8bOOF1nGXTgEmadA0w
6R6aQRdNIib0pB3K2wOaVj09SMLiZIygrlqjWSb5sIMU9L2S7oFgdyD4ZuzvdmbdzieXJ0tDcOP2
trCyiB8/T4YV+Y6mc1pVCBW7OxeU7CbClW+qSiuxW9mtKVJWEnfpD3eDFIzlEBwicaAgHpIk0nNQ
6QSqitUpk+Kw9Vji7a6KH+8y/muSZH4TivlpDKbRJoFLFgytMI0eDq3ek4Yx5r6wruysOcOA1ETJ
zrAnp22qvv93Z4TDR0cTc/qiXAhlsUm8l3TqTDLP03M3mJIZXIX9JL1cfu8WyAitvbnZPtAdLjKG
KAfRzKhs13RJCcgl2vPv+nHHj0vdED080pJs3MeWaQMMHQKh2PkwH3QvKxKqs/ABeAVmsW28SliZ
Sx4dZ8nI1R8KdnpcF3KYTj94Jljv+Y3bUs0HmwLboGXocpX9FHLtC2t87UOBaNty2ub4IWwAmCEO
SC//Xdkh4r/CTZr+pbz33eaQWQDd8ZCajeqz2xJVerkEOl89aa2oTLvffqeTmjMmE2UzQJsIpb3Z
RML6DBx3XlhUd7X5pqLHgMGwFf4fiwCiQekdkQBrpVujQs5aHfWACV8IskrRzgPL/1GipqJopuBE
yugHrB94X4KdKKdGpdQeB7InAJAFmph1vT/BqtZYLzEPlVs5b9vAG72aSrGlcH5wi8rzhk3c3H4f
KS8hXk7MQAaXr2gDrU3XOk7M1JigvExXzhv7dGeP5GVoOMRCPaBsCuusH1E2oLdgVBItRIIzgdpa
vPODMJrm116458/ZTm/e5yz4sCiHW6SG3C9C1aYqIYGVxuzhU/7cXFvXwKf55OcGNkMwJ120fN4X
Vai+skMsdKkUkKR0zWYBcHgVnzrpVjY4Bab+iz5NreO1WqKXc9/MaEN3U8EwFTTbUubTfBHIDklH
oKbOp4by8J0nH7hANVhBqGOTtfUtp/ca4iSAQQdkR3h8fWk9QIFJBcPSBNvI26LYnzf9udeFJYkY
6Rk1c/mYZPsn8xo+MVKsnJEdqRfMNRaV8kSfCZng8IIcjHjSaq/MGsllL0JVpY1mKbUsfJmSLw7Y
RgYMQpg3w3jKLwi9om9XF+7VBuwdXfQMv8TAZZVg5k8P13O/P/9a+OHaUypWPHzRg73EkcUO57Sx
JBHtRMvn42k5BroxQu5/jRFjG66xsbMDoYHZqVaJP4PfosP7MPKKEZB1JRV7xii0QIz2VltcGSLn
q+hidl0F/Em/obSXRF980SP4tcdLDO5M9EyAGEcjr0wS0uRBIZMR3NtiqYtu2XrsnJFrB/u5d2O9
Gh7BULddBfn/EURKz4OL8nBm4F2TdSXZBowN8z/Vx16NF+uHrOxO7AUqLjOrEEgWOxV1b8kyoXnU
4zGsnCYTl78Ilr8EkO4fgh0CM3MYo1jjg774RxPTX8UPpCmaMJ/fyE4JQmYGtpJnaHLr1iaV9BB8
GKb4H/utYkahWjBgWeFU8DStl9A1D9Tj0o8aRqL3fP3/YP/ThHyeEG19xsUw0CXHRvt13GTHluBu
23HGBY+FYMwIDp/ziePU2Vr1MbVZukO/VE9+xqR//O0Ls9K8HYdhFjuaAHO3Zc8e5UGMePIZLGJs
NJPCd8R4yW7wE8duTToeaNA7GtVzDhIJWaUa6h/hgs12+gTDgvJ5tu7i+n2gZVc+a/53B0mx7p7K
BjFxnN3DNomMPz7/bZUCMSzRZHKtryg6a483UMkNNCczSVnCp1EsdHcc+R2oGwgGasoKuA8pzwgG
48W2jOJ8ZOXM4umtmukc6rWStijitZkt8oNk8eWnD/gMP6t8vgi6jx5NLrTLFde1UdE1x+4C/lsK
yQPAN/80vHvKii4IOc9CigvrWD4hLoHAI5B3bvBskvXOiOHj+h/FVZRrQ+Qu9i0rr4gGC2xXvRGK
Sq9uXgbK+zRUM7nsDRJObvVr71GMOVF0mgAOYx3kYyZe5est4NFhNbrj2UEMj+e1fq9k5yryoRVZ
hc1CPnsowkx93DzVmZwnMu/+qA8GKZCaa07yxE53t+IVNZbEax4IRQ7t5VWsjLsK7CI1ujWiCZQv
P5eBPYigQhjsy0tEGZZtkirNH6wpLAqAvFCD74dtC6L3Imz52Z0gFjmUeCIvIEGL++tEsk6jNesV
8tedrKOW2tNPWRmqBqEM/7JtDbnA8sgYL9jiefCLtUwOMb2hSqy7jdP7vlSi35mqaEErnFBCXHyy
BvaFOE8S0baVb/AqG8veRkd52yqpiRIRADhC4t3Wtoh6g7F18ylQZ+qj6Qh4DJc5A5IDjk+reU35
8jdWfxZ2L03Fj6EyRmV/VSbGYzhaJjEmq7kZjQOyKt06qQu/udcbFX5Qyv31SZ2Zq1EfiRnlXQND
asPK8wRs05L+rGbxit5kOksR7ELE/q4UyjUYsdUnqy0Udd235E+i1G8iNCfYgoGLO+Cmf55bOLFM
xH57bAXJXrYX7ifrzDtSJg1cSAo89JgsGcJmAyZW2+9sGlRIAcBo7NoQjxz6m2M4jbbrARD56H42
RxM2yTT0QKtxyKaDPHPBsZN74mOn0EpXiDHQfAqxgvzeImbj6JXcXVVzC7wPfoHXOfaWfBesANg0
1XFInoEc7VktzjB146ZDFl8zB9vlWzPrI2dVmPWfcSvwhqTF7nLmePbOejVbx+75TfpbouVwaVXQ
yzo6ympo8pCK9DxB7tuWlbF2xj6SsTqbTstXBKj9pOMkuJYbMsI54kmc9LQd3EWCu8WCelcfTlQO
jyZW0Z1wuJWnKcOuS6vh5rNNUuLFVegQsT5/2+1oJ3Od2AylF8BXZwm0QcQBOUw5iETFj4dMIE7V
AT7ie6mtJ9LUFPPQIDaSfibx2gSLiGrr/VL5H6AJhrFNfSlCtXn365rAJwaKe7/CQCQX63dLjsT0
dNeQeagKqw+ToQh6NOqHQoOUAkwA3RzTca2pIi0yFR2IOdPhiCkMDS4KNX7gfgtR+BvTkwgfwCRX
/Q8NrJartkuRsLJBHUhc5Z/uKy3l/I2j6Ed548dlw0VGcDA8D+1i8gm+geEg9xbRezEeco2CqVlB
JQQacIyRBb/7I+RXlEQr5PL0skgyGH9MblmS6B8ME499oPi9p/15dUU5oYFNCJoj4Va8Ixx/aYmg
fUfRhqmrTwi+LcFsB+TBxQxFZbabr6mTDMHc/dI3szFThrrQfHmnT+xntGOAnWwVMu6Mzz6ztKhG
BwxbHVLX8imD0wTEtQ9zzJ+KvCa2uT99UMzHNHFmbt6SWDUpFv+xgOOk2hu5UCkl/EHRB91mdKJU
SNezNCu3OeKCwzox9pb5pEPFytBXxU/Dy5bGBBa999DxKFgf7nFUGOCHt/oyCkqZrk3C5tM4ZrC6
2tEe8pVRrYEH5zLMhefruSq0V6lDU6WvdraR4GWzxMYG1pDaGew8lOMu87QMJcimIQYuX7p/MybC
8d5aX0W7+MD+d6njJvr+409oK9uQKgOA1FTXz+gfCf41KBvgKfPVeCugZnH6Nc5mzoUyuEXtzFpl
qa6FEWa+CWS9NmIJM6H3ak6Be74JWF1KUs1dWcnLNB5+C5YD+u41onUyGidBDkjPxQZizRjk5YO+
ZuNtVs2UnSJBWZT+lrOC4kC6/gxH5iuL+gQ3koZ3B6fv/SUlewRk0q812KxdHYHkxMVTLzXRQ/st
DrKHsFd45Y7XFhyfSlKRtT6K8TeCSAVzYKimExr4glTCe1NN6jyszanpsppxv1CJIO61DP+fdadI
kgg7yQlwXCW0SdqtrbyEMkmV2NeSfM9ZijwY6jLloCWiIipJWn3SuFRo8Z8i84gEXpgG1idbl1Ec
v85YAYVobLVWZwREo5HB2lJa0dMDKV82/lWTeuzTftQA5m7svi6RJ/fH+J8TlBGGS7Js08Z5tWKS
PXU6xjMixQtaps9FD2kPAhuLD1CtK6A2JhW2TSwZSft5sf7pCjsicL6phAl6wSbhzYm3HZnO3Q+H
/M9sB2VraW1u20hM9EyuZe3wjmaWHs2PoylgGWQzeElPHkIYJvmh3A7bpp/I/ed/oem+cgc42C4h
+izoAXCpmbzN4aTmLofZN6WkDJL4DU3dMeWVymAYwqKLf28jy01DjwbPzKdbDSVzgGDjQVBbGjzT
y/G4IjzjNBuO3EftEPmf+nWmCMsHzv//F7yo2PF/BKyuDNA2KAhKPyNkRw1329sTNX6jAvuMJnsr
LRbfTccHJ7kt4dSB+SEui9Il2bAPpC/tDiIzsun7Tg8pnaRAXmdlqZLqBWjH/hGc0GZK8N2h6QSf
vGvWfViOZ2Mu8gOQ4kfiaEVo1O7xFzHrr9BB8J+DWrb8+so6KOCyMWEXx3VzrX5WQatY9YxNyDCF
EK1E1lwDYHlBp7RV4PcvfjBdhlBOLZRlTXJcS8XI9UXJbQHxazmDNywOJ14kPTUQTe+A4nibmxAL
2AoAmkfVStIeTsYeKNa8r1mkVMA5/l4v+2pK/zgtgmnlme8jZbKeUjg5BHqpFL3vAAyiE5UXfwH3
Iyt9AJXkjWUni/B7HOqq82JdkbKkKx0y4VbrYXFFdNpb2zHuQ3BaXA94zMSCdLcGeM7Mcx9/2qi7
r6GIbmcSDJzt1kcLHN1EzBeGpplQOCb2LhzRi5umYD36Z7ZVjZW7jisT3EiNpMTaH/5v/FGx3v8e
RzubS+XWm4aLHMIKITY5FXDH+30zY09AOwS5VEVg41nJMbgkKqXF/xiQejAR8+zf17t0UjAeaPzg
ULniQwB2bo4FfnXKl8jTwuBvF/F7tKFo0jPcMXqU2Vg1DhHyxo9QLsJK/hj6KmHufR+7OOn2Gvlm
lTKlJt8/KMlLHMQLQwbnZ6AqXGpZl7GwZ5bsOPAPcz9rIV2qfWG4JD2RgHyadC7VHHV1HDC8qkkN
p97Vo74gscnkfsYKkC+K8oysTysfU4gx5JOXHE7pgiRPsbhNNpU4rIxWDFnHe8gv0+0skKiUSMed
hSP867XnncqoMrekxvJrayWi7w/0yVbkIuGmHOLIgLS9R0Pt8cx48N09lqbmRTjcMOFeBjKcrGyQ
+E42Z18ko9hKYQ/SrPWExWwxqjV5H6QHyKnqCrZwRQs4s5FsMEOk02PEwfBkpiQdaE1z7/19+aTM
uzN/nDLkI0Td3sX+H4iDgRCCJq8cIh75iSFGLdE/Wmph9jONqH1ZMECpwb4milxMkIGyZ7Xr2oav
Vb347rFOrgCQWQnKk5kbN+Fu2g+KLB1ncUCW1ucrluuPrRozwTsyl2eQBqSQSgUZHuXbwJkrh6/T
Vf/DakFAxp5QYmmtAWE/8Nm5kpc9RUG/x2b6uq8YD4MHTAQKIU4ELKASq+JXwV10OtWc6a0U0N4g
NbRRxCyCA1radvDuXuQ3IuIfFnJwrVpk9XdkIAXsY56xj/qED1grL4KE/ekOXc1FUUIvCOMqStGb
CesdHjY/5vQk9NaVjOv8hn3f/d3oA5reDn3iLbsbGK66HJTnlbY44LPSQ3Sblo3sfRC52QVLcWk/
82OgCtJglemu9kkFItZ4v22qu7V1B5j76NSlRJ68vrrVo3tY9l2QBa6WHv2o2SCmnkYbMgeguNVP
d9dZ3fzo2cvcqI3AShQJkg77j9RtTLXeUqtPHU+sfjMPUyjxrIqJurVCX6kEYDKOTzDimv1LZMTf
09E51rqWsfUPAZai6avFk1hYOJLWHfhtAFvXN1i6uQKtDac+IWHuB26NTXV+W6N8v3Rd/cGEen2s
zbFj82kvV8HPleFDpOeBw6AufQYW5GafOBeSd6nZ2GUBuPE7LXRv6SzzYf2VyOmWOEFfUvjk6l2N
VCJuA9JBG3H9eO0p7NEhd6ut5eeObaQ8RouWw7ntoRAYNCnm43g+VN6tmgnfFPC2q0NLnMl9tLPq
n1SZhx8hYmbkikqX0wI8Ja+aiaY5C4OoCb15/rhZmvojd4DEeOTHNj8bta4NKL868yNCU74KB/hE
sSwskXwom4vZ80Tekvl3u/eQEtr2b5BV/WT4jeZIq5GlsJLY/d7Pqifb0j+P45YKL8OCvrNhvZpr
Ep56iCuDw1emaWJR0iEcuCUP5J9h1jlOd8u5vc4GLGaFa9qJWYcy4ae2E96/eyskKpUScjg1T9ya
URCRv9y9kSjGKdCFshuhM9RchVKqCU0bgmd3J9LW0AAjAcNZtGd8aawU9wwxkpxpgNHXUHKCJxxs
IBsvam+TdyzH3m6rRzWr7+JQ3BAfRBNAFEnJhFuumsrwViCfdo7u5VCgP0HrpOw+LSgtRE9NGN48
VJw30rrhdSRL5oJ3XYcsdwT1jlanfU4YGl9jQX9HY+WftIyj17AouQFh7ITnamGB2e6K05r+INym
Na2iv5fOqa1SdMpuXWizkJ7pmWu3RcmcQ0pyAR930wNDGZpzuTn7DVPauLfoyzzejgBOgDXSBaNF
Qvgsp1fuEDBn9ld3BqFTXc2e/YjC949yePWZpHd2lXnX73kGdT03e6wdC8f/IT+tuffsdmKnpIE5
BIxUP1veUWQalURajaYfjT1zxugKJxeKRKn1ELCbtuk6tB6w7meEtT5AjFIEQiXbFijLu5OmkmsJ
EUBqpbAHRBTM7mhBEnLDXUAeW8/DUDXyXA35bMaPf4LXDI1d4myPk+e1ZPJ6Tnv6fIfo5+nW5/AJ
KpDxoqXDLIj8F/iMJSltvVAilWASylCmddiu3r2+Bz8LUqcBJPA9YZ7NKrMrrmpXOySemNEIckjE
4a5fAwjeNRGKz9loOoCVKqWrrD+G+5otI53+lh6f2ArZdaIrRec7nUqndW4xYvccicBQkPnW3zEU
P8zDQz3q0Qyopzs0rSbVPrkhhcopoz5bzRLZB8imoszsPEyR3B2UU6yTfhlJN4X81tKCUCw81AQF
xNc0f3dqoXTx3uHR3Y9K11VHLTxVtEza2RKje9s4HSSnP4VNZaCT2Rv4R7PD9xwtdgR/lzL0gFWa
MKFBH/0fS7zbFaWfxi6ULkbeIZCVRhhTH7P5fDJPdtZhTfvET8IGHnnIXGNMt3CIztgCSVDp+3yu
pjzLZT00H4hD3WpMFkdl+N4O+dWlPWVhUTNk5G+w9cbgPkCFd7LXXdTNqvWRbxvaWkmom5CG05sP
pq8PDs1esvkxUnPFN42igbM5NUexZRp0NxIlELKMwG9pREHyFuU68Rl7zm2rLHaSRSpC2sfsEYv9
mIJZ/XaKW7TZeUeUiXXAseV8B13kIRyEQN/RswzKI+BB3GK//CpyC7XLQf5bzu9fFzSDZIMf0mVL
MutebvKh4WUgYEbRUKIrHFPtSky+Z058z5Rc9xyfh5Qp1SWwFlJKZnYvyigtW06EfkyWGvxas98u
IJj3EKctop342gonnr/e0SnwRWlaAgJE+xRQR7U7qxY16PrQJ+gWmZRD4mP01IG2wYZWaojJjaWu
HhiLRtXhZmU/C1YIDQFYM6dsj7JhOh4UxvcHQ8PrtWXMiMvC9BNVaJeQelLEyZFchWbMP/hPV+pv
XCLKqMOuIN6GpIk0fL4WsUjSi4/00e6wnGwKsUm5MHY/7eH6eySbTch1mP5XY2HFoUFNK3VDYlUa
TrilddAHTSb2B4ch+Iad7UZ4W0t6CW6OBHqj7OC2kPGPVcOB3vvheauH7hghaOWznMAO1NfmBU1k
kxlL05kFb7QqdXbPR2vWxAAt9YY1zqKXD4iLfynhHu4UoMJ0c3/Sge7JgC6pqpj+KMCLv3Z5xMMP
OVDO9loQmTvVhdka+trlpW3Tmos4VwQbGArpoh7tk4QCik0YLWKTUgEpDUY6+q4+TKlhiPRm/zV1
C1Ve2MMXALFPmDCuIvVVhHoMkBBwMtFVvMyINnhm3U+oZmHnuaINxmuh+2nUkhox6t3HlRwnElXr
EnlnXjnz83fvdzD2kS/0VPl0wic1XE+m/ZgWQDJYFwXupuR6i6ZOdzj0/prG+7TkeIy9iPw0udR8
cDvxVRkYCvfDlIJh5E4DZLKXrdNVZub7esGQBibggdvWvtIIhLEhBWApEvf0U06e1alT30uDnH7Z
s+HGIOwQjYg72tZhexJS/4bDbcRMnDK7sl3jYSA+q3aF2CPc3WJmQbMIciUeEHNNARq5gSvFpmS5
0My72tr9wpCddd7fD0hxK/49N9ZWJFYDWnsImZk0eHS6N169JJD78KlhNZO3ECUtWdFfjkYv42rT
964aVC9t/SgogotBxXL6v+4pl6Civr7l5G6SGCXf/v+zVHbe43qu/9/ryToMrceSgNR0+f4Keja2
mHb+bRQbnIiIkGMXmf1i9z0mP8sr9nQNGT7NL/nHyz43or4FYBvsDbXYKvyA/efsi9Kkd2TPzccs
jgfKQvPMNy2+gFob+3owhPU1Gh73HN0NZqhr1ZronZqhIV6Ql/luum/3d68ErJv2WALxZJmX7TgI
yt7w/EVAIgx6a87E+4ewR733+9OQD/egoJJGr6Qb5sfv0dDGsYcu2ZdTDHUIWnwfH75JK4wY1yHC
NOkn3/3IMrCPdLb0j/HKZ6BJmKsz/GcYCVUzwK6PEt196wSJi+bf+f05CVYvW2drnWvV3OBDlCfP
j3sZDErg4x9xnsPVFMqiCxft1bWmwnzv2mQ8LkhyhzjECx6Vl0rS3QRWMMuvBaDSQBIviQh9sHsf
ykomragQFzJI4uidYG/weiomZaIz3ak/ZMe4eCrvpVI3G5TQwOxQA4VdX/lvzMM/ZS5y7/aNWqGK
S2TXz9+ngpXdfd6H0MJxoKj1MRNNoT6GRCVloJbbXs3OFTmzKXSbikivlNpJl7hghAC8J0hj2QKy
Cd1k1JpL/SL+iCOUHavFMq1quUVxAWEgC8j/geCKUgBCmpt9bjJqHALrKFNdWlfTohH+hO8vUstS
G55V34/NdZYPKYoL5FLjawxTepP//9GAm8uC6DjTWCV/lhfFrpniNVo/LrF5fGdvtzxf5/4xePeG
ZpXrMoRLaFLyI3oC4XmbYMsHDaQVPqkxS9uzAkqYzp+dmGCXIKMeL6HFp/IR7UEmxTEQAu23Ms+Z
ed2cN74C7ctcaa0S+4nO2nKntgnOxVKABk/k1rO1/oFT2ZoKRzpsE+/g8V4+dXIl+kK+Cdy7ZPRz
wxRGbTXJc/y9p12OPq0xOpXPjOe8HZgaJR0CaSzKF88ms7BnBLeHjY0/vLpyXkk6kRYqSzE0mgSa
ah+dkYj1A5FRG5p+7oMJmVNlI1mpTsWuJuqASM/pTFu9R3JFfwu3iaxjnAXXtMym24Fd7GnxVp0y
XUK8Dz3kcLvUCKDgjGzO4HUcmfy0tdJeE16x/vhP4SI54ZMEfUdOoSV/cUeqeVrk2gWrthlkquQ+
XQHV/b2ozpzQrD3Bu2wwbSgxc/wHdh1HdJX1kY2zuXyEj9++mbjLQYYGNSxE7NID+cinDxSJXH6A
1D91b8YGkOWzJP2HlBpdTxS//c1OMUba+NHPFQbABhZa4ZMw8SbjqFl1t3loZRd3zkmWDaoJ0Uea
9T2benTt4lFn5AHaaedhYEnaeCF0/PiTCUBzLpTfkt58vL0NsqnzPy3Eh9FffCMbeycNWt1wI0Om
CYqDWjjj3YepsSRmFgQdicgcI2CR1DTW4ywsqRt0PLBQEKPXYyzTZWcOFm/lg+JHwkGvxFvnT1xR
E9KcX6/ChZMNm9rzHvQGA8nQoU0ifdYlwaPrjqdlgfIN9z2vBP3UVTZPUgv8LI8fhleE60QVTtMy
hSo6koJ7+ZCSv6AAANvUFE9tH2RYIWIKvgakJ6fWc61Gviibe513h6JeMrE9AWLiXm+dEe+Ei4is
lUtad49yKj7x0SZt/VIRZ6eb4N1LF99XQw/8ckHpjDjPst6eujcHwhTeNoQbGFwbaPyQ0Mpqu7qb
FZqr4i3BAhrfShYVwT0OL+l0fLZpTm7Umt6q1iX0JTnpDaBLR+bjx2rxFQ1W8iRkSYGjzPycOhjU
VWj/jUhcm1ntFJGD7bIBr86BZeqPAiKet2R5aaZ+tbrcDknAEGZmnSV9qaDzZrWC55q0UGalNQwP
xosgdQpcCF4pEdNEuqfJN9QoAf9smoxu1hEG1QDmTGitfgg3HoJcnKv9WM/403c5+McIRE4aq/eu
GWvEGyhu0ppfQYjVH2R3Yh6UBFKTWVo0JvyZr2TaoYFcdhoil4B67duNpAGwcgCgqDcinV/pWw4g
F9DJRhxv7crTQ0ziYFi5mFhqkUtm1och73tGg98R9C3RjEA384QGIxrgJut+gwJ/oefxlSYbQBZo
triEGZ5e0m+U81uGnYjaHJaIqQr3MQOU+4hSj8+EmvovRnYDkyfyzrS86D8QVccSjg/gkP711uAk
SsnoxdnzmWqsXjqyh9KM9tqv34onqdKQ+8UFNZ/Uq+b+oleGkwDLSFs5M43chjmc7nSCZsFYtfVH
wXh9fVQc9+f5X7VLWU6iJkGfRkEe0Oo9QTHQGP1iOVAuoc1+Qp1Geo+Xi5cQo+0Eg0Zmknxwo8sJ
ZJHgElmLYmKqHH2zHuTDQiS2fNHHeVO/v9pI4t8pxyrogecj/zHrvy+Y1k//HBsGPJ0KDD7C9pky
7LegMVITduaL9deBHozVxeMyig9TKI7ArmRu6Kd9l9Ibnw0A0HuYXn7W7mP2nuYrQCtWYARc81Q2
FNajuH1AgULdmKq60Bf/WQ2WKkHyqOuzvcN+qN/m8kj0fT4HABOBVHoXfvhxw+iVFO0o2vLolHn+
CMbot6FaF6gQeEUQgXDmEyNODJXzUGMQNo+hXWHfrGsz02B/c/MX1hwsEenZXSdSlA+Ld7yyYPOw
hc06SB544rHjibtpbnRwKh0Pzo4DreXvo6FGMTbd3a+bjVsKPQ6MBAGDkEEZrPNz1DRFm+3ADKdc
0yDe4PNsSkPbI3a6J6aO3zEJgiNs5d7W6JiLjy5haHVShmdheH/EzHgdOGJh6KMCXnr6RC5DQQer
l0+ByaaWiZRABmOWV9fWNMBFX2TqKv7GeWHjuRbdDnouff/00028kOQusRBIOJ6Ta+CHXUb0ZaUi
IgK7vcv2GKPs5OppYX2IAPQ2+UK8J4lIn1LKE5NLsMfvS3YmSjT9gi13qbfqJOSHr88L4Dq3n/2x
t+0yafRkAVGMPBzLyA2PSZKtgVJbPaNNfg7Dpu1Q6RoiTUPyUWje7YTozMteRVtb2oNzCsoTN1HD
fY6elLEebkbtCgv9mcubyBtq80Y+ZodQ0XCswmwojzwfq139CG5lbFAWT9m08lQALEH1zKZ4kYSE
w+vm7MJaF/L7v3SqWHHRqdqrwFaGr6o4ojzteiwFBm+ilpTLZlePEQuiZu8al2mqzRWPHpyCziqr
IlCTwfwuCkncQVnWgtrj+tCPSLxhMAZX8Z+UMloS/AhJMuojap274EI5I+fuf08dZLbJ2ne4x5Cx
4obqQr19u98uq8zI65N3qur357uRU6rkrWFrKZz/x/VEAds90b3mEo0a8bDIP70r0iJhAmObysCh
zlAR6n4MW+EjSPVDY4MQx9htA/6/DOgJDFFOLJw9PrSJLPdK+4ccbzyGYrOrI/I/K+F/eIb+FoK9
lyYJpm9Aa2iYphUwlmTBR6RpD/YQMwO3L07XsgDnF7sWsRJXPeU7XSSL8Acr7zdVEzaMpjocYYea
peE8HYNKw0TBCiN1ONNwHwAwg5fBU3PwRsXYTvs1jqbR0Twn0YP/IcR0sLEjmL+Q6SaeDiaRlKYH
V5kf0hlu7idTVE9bxX7LyKWHYAUvCkJcTd2yDrjfXuTzCXftg9OMaB4HQaYuh9xjmTmlWeLeBobC
xbnyUL9M8XWaxVvK2r9vrGEvDdhIX0SdMdp1ul5ZwzOmbrCsQpbXRxlxFpuaaDg87p5oKkKkwwDf
oW2EVPV0LQbWT7kNXmWD6bhx3AxFlKesj334wdFM79xcpM7aOmJLqED9nUo0EoZR1+frq5EHWYH0
CnNd6zfrpHdpLH9Duv8kAkm6HnJUF7bKT6tHwPD68q3+ZQ7QSKc1kyeqtgYlj9d2fsK1vDKhxN8D
w/5MINWIqub5LPguZUxT73q21eQfBn0tK9L7LSTk0SR70oVr08hKwih/rHv35CxrKlEKrW23qGJv
YNAbeKp3gpGj9eOdYAciNxDXAMZAOuTUeLioUk7mFTXi8Rpxw+VgUtrNPJzf2guXAP8XSY4SRuPK
zuNo/PceTA3qtDawQRqDhLEh2GUAiK0G31PP7N+xiE/lAvxy4WRWIRrKar15JsaHW8eAIgOJiiA1
Rkf6G5QGCY0oOiAAJo8oQ7Uj5+DQFXRXmaMHCQ2W16UXQuunZUAYV8emHiPq1xvVTktXHy6z35J6
Jvs65H9s49Wekb3f2h43qChUbpOgfNAivsp97+nE05NA+Z2XWczHd7LPv32blZz1SULF35YSp+gP
wFkgEUYRAz856H19LQN7gN1CNaDVWBzdcdmH76R4uCSkPQ5Z8ykXnDkEn1LvsWZMbIBUAkxSo9bK
T7RfInt6hqVFUJw+WtTC0IYBbYjPZM/HAyOOyu2f3AMZTrcJYShcAwKRRzTV0J+zDwb4NYZkMd0f
DoWznYNGrdUFhmJtWKy5uKNlXFazp2s5rmM7tAERhV792HW6ekfJa5A7LA4/FIfJmmR+ev3nVUJz
P+gfu/oBddLRcJHBVplQHTJ/2iADVdp/1TYsAFvPOqCK+PeX5onZZNWxX4og9RCJcn0coU40FTzX
d6JFH7BlJRGtCdUio3GryrDAq6Fdg9deecv79pbTqMlTq9GUk0ntjrSZJH1Roq1FmQc2tbuXgblw
83W9/jJLL8zHYM0bf7uff9vVjWN7PJA9VMMkGF9c8Ir9/3844t68/UQaBMslRXoEfCkEbQBt0UzJ
YYXhZhRZqkXtsIeTMxJ7VzLMxzYIV8dDMEqUFfdivZ0QH1VkI8zi6oE1wv0gyduqnFSJHW1R2l2t
xBGc/FJBjFImaFiWMad3j72SYcyaqO23qke+/EGMFbNlS+qNWwPFfUU+XnvpBqqSkoXnPzEBpibC
a1ZvnF0wxMtchFpQSevqSQtt3V6MBruDu88HU20i723zmjH7PpOAWsGzulY8iMIsfjtWo12zT19G
rxFOdpIHLisQbymsDJu20C8wloz6yadPMOV7aiWk+sFsMqD5QDpUbolSSB/zGGvp/t10WelbNf2c
y1CFzZCvjw0/jC55bF8GIs5WlM06vMZ/3AGtHiuaTBL8Xo9HguOboOeulhIvZK/rP/SgRg8jtNGi
DWH0lbFhKt46BZ0EYbIxzTdre6dwG1+3Go/Qrd2+Qpz/APbrz8C4i7a3ANHKVFUTIA0j/zq/lg2u
MuRDRw/WESCzWTOaORXw1RFIsSWUQtSp0V2l00ttHAcYPbd7OgFUH6TLJPQS2hIRYKMO8ZaCiP36
8Tb9lRHU0ynfSk3S91CQE/woAtyToS2oZWDGaLxWPdomOzpXPO9ZhGRvlVcRXFBdxlyQkWwSRYWU
mH6SJ1IYVpEH2o4kCyytiBrUC2tD54gI0DY7YEkTn7Lj3SDHadyfvXHVjOOI9H06g4FxybQOMhgo
hDLbIfLvQX3hD06rLjOSoN5e6kOVUWb/kPcQEsg45Q49hsaY1RCu1R1+uwRx26k00W94dcXIQxJR
JNvVPK4vJWLLy68Grsq9cL5hfTmWBSyjpYfhXpy73JTGezDiRwo2bx1szqjXBLBF8d7kcv/PSAXR
+rui/hFqS/vGllGJz7tk0a5uZUQlu/0sGDG4UwSYFxCsqk76J6BpxE08aBQxt/Ux0spImRLQadYp
+axf+1gmemMqsOn7W7076CpTU9hqclU9PWav1jsAnQYfGsDUEGH+ke6lr5+UtgPd507vSyRL2a8o
xBWOrqDs1drLgP7e8gktVoP7GAqw7Vdawj+0RGnSECcLTjjB3eYZFpPwiwNJuwkTv10fX+vLydVX
MLEFvNwi0MnRlVPJ6+3DImUccptSLpaWjo4GF18rkE4bs5HUa6pkBx5e07PrSB+IuZtMKMoWuah4
sIv+0UWvMJ3YJJKslEnVyR+4nBwiKnH+lTD07htXl0TmMz6kCdO2lBOgd6zr0Y2vNJWLS9sIaoUr
QIM5AM+X5US23vubVULWpxeM7j2YGtYE8EXBxo+dLdKoHD5VIibaJIdplwVgADF+Mv77nvLAQlvt
2Az7fu4LlG4CpWGdC9BjYvm1yFNEgo6EP6oF5TmWph+Ib9nMQF9CFCx/KDM4mLAC8wK9uhFMvh8P
lHiqUmWbJ1KNYvfjgP7tWxQBBTtBAwM/p0/0YQJ6iZ5c1WXBgm3JGXYcB4uUpHmPewEXSh82FPU+
+PEC9NLXYttdRkjkq+CD7ALmP6DwfmwlwzuJ9Mv72KPPw7dR/J4VOOd9GRb7B4toXKmgu/NPhzZa
Svtlpqe6QrQUnG6+1LUL6e0eQZ8qdypGM6oRWRYrnBrjttsLI8T/jjR6wbwtLe/LY1061IDXEG+6
9fIab+OvWqhCOwNKfQe+K+a5hjAA7umZ971toKAHBrKnsQa3vTFxQFLPGFBuM/6FBezAQbB+tTLn
BbXQ2LKJxKWo7/TfZsdp0wJJlHokp9xFoZBpa4LmOmttJ30hhG+jfuUTcZUARxj+IesH8z6Lfrl7
0k0ME11mJusLRUBy2UvRUZL9d/gdxfGMrGo5b8zhnEYwm//dTQZ48ZaF4C3+suc4Re9y7Vk3qhAj
JpjAcZzd0j4MBMa7IfPCFUGxJ1oUmTG4InxvqA2ndjvGdnq3VLwiwmU8SMeUxd+vZg0YqnU0W733
mdKHeWONypZFRRIntwXZAcUHu1eZQ3ngBY3deeUppDAZ/Rj64Sd/EL1gDso+iyYpORMUK53OQrEt
VzS5c2QhxJb7HB7/lFNSWO4rfz5oh+AS3q/xjW4MhvAv9WCoS8vqqe8OZw5q7YEYiaqyz1S230oX
tfUlK86mZ3MqiOzT24f5pJb/+sHYe4A7u4Ur91WsCL0XvWSWOdUOieZHiF4KwxUmfyp4d9mFQapn
86aODatS10LJXug68Eu5BiqtBeQHj4xnQsTbOTds5eC1oDIzuO5bTLhzuMrFy8fEcNtJdkGIDt1K
O9qoqVU4PK9l18lrgrPmv1WbwtQm8B18hRaW+cbARmoSJgyhng54TJ3ePEff2oNY2JgfMM+FioTn
RKfsPhXyvXE994h0/ucwrdNCIrR5Zh9mLNNyHF0U0IRmhCRD0J3NYEld/F8YPs5YteSGW47yZmNW
S773gZ1DlBHxprYOhhWIyx/NiitG5nw0QM55+9u6HAXcR8XOe4AUtu8EID4TBju7PgPUkzc+Ntvj
hJy6iTQDFc6DI7khW5VjNH2CCcCpk/sqcw5imzVP41W6NEWiQwJWbI2FMLqBi8YRrw9G9kZFisFK
sa0VgKN/BvP+6oTxfHnCfMHe8tZvUn9LrrnUe7P/lDnE7WapDFRR1YRHt2bpvWszr5IW+dLT2RmG
zzJfxHUAJXcEpA+uRH2fCeJFkClagzHREXBlrF3uD9aasKGkrFKjTHDivAVLPGHlIhHPusU/qt3o
fbmkGLlh9xv8LTgJXhAzLzYXBOIzYuffD2CRX3sZXYgx/s0vY4ZmWThvmG7vSW0T/GKIrnIkhx2e
/t4oFQagOBsIjukDvcspKCYC4mEu0Ea0K0n8BOrB3TGzpu0oyXrNXDaqNVG0OUoFE+oZ5Bh/5KED
vFCNIdAjUu2w21/5Qsw4JDpaoOFWP0K0gyMDO+9X1xoqVOJVDRy41M4o2UX2TOXyJ+fpt25w0gZ0
p+GYe2p5mn7MIORqQ1NnrOen5A20tQ/Ki4MOu3URrjR+3VZOQXYXVGwJHNed+RQe6f8pFV37f+Q9
X11QhVqbLB03vve+0tp0kWlJtjpuuVm0HEjY+nYhGLTzwTyvgDpG48Em6gw1TWPNhCRa3CvXQu8M
ARN6xKaMD99y3NadW9KOUcdYIYKkDrgmlcNxGEz/l6lyaUhhHrox3nJt9pkdXMP+C9LNsfNKDX5P
5zDOCAOIXNn6+UtAauHUyk3Enku734sG66irA+zZAMAP073C8381A5nweCTTXOOX+0NzKby6ALiR
9+Or8Y4yJV+53VLx1Ki6/XxjyqN05BgFNDZHy+HrK06P4TvZPBN15QiJfOO3csBpzfdsVYN3+E6g
Dz6sggwuW2idN7QadK7uk/q1akjr4srgtXSYzl4chDc2VpPpOErCDoF7UbCC/l6TtPvUipXWCKhM
R3/fkwXZ0jmuEjj5+8Zspbd+50H+UHL46kX+DIYJC0ZKG5sXQSnXcXBRfdjhQDxLfdcy4calWwm/
2sgI3b6eEJ2KgSCJUmzTbagOaJx3tSicaa1ilI60V0rzgU1MwsUWpz1M6PamS/Iw91e9t5wjZLpD
sCK81Ff3TABlrRf7RZrb9YVFWYm9SrqTBqpnDWf5TpnoDsXyCdNlMvHZTl0ygh9IHVqY/zFXNBnb
UeChrCeQXppukMJSHjztelw0Mp42KcXZMR4jKycCb+xZLNu97CBOv6jQg7RdNj1vn0guxDmgggT3
0+fnycqQC5Z8TN++mRHeRfm0hwN8Lr/xl9TFxEpozaXZSppWWG2ldyPL9GabjPO1SVEIbjn9IvxO
Z0oaPAjpIIzjLP0TjqHGBRdF/2AUjwo7rgoYg2pKkspzgM53r5OYVf8muZOL/pmKauFNx8ldhwVP
dXBfY6c2WdGLmZJlou3FR+pgoAJNGYHFcUMCguKhm9k2ZtaM429EdZYVvG0JQ4f5VkY2eUTEPofL
E+o4nITLJdU7Yk+vq8unE+TTgkPawChT5Fhk3bzLX3NPMFYLR7bd/EwhVDvEr+4vmoWCdq5lOaH/
71yhrlvO+TgqiHp/h5SyqjFwnRoqXvvUnUoDfAGdraoBScJ5VIOfLasbnJtFo8H6p+SdFQQhVPOh
Y834dJT/Lw0UZ+qShlyQYJfLPdvhOyjIxmQNMFCUilZjXEvUBQUzPG5FsfYTJwnHoFGsXLeMqXq0
+8KBfdI39wDk4fKN4Z6K9GezKxAvQ7F1Dn2RE2FEuS16vmlZsr3W3O5RBmzq133kDmANRHRqwGRN
OCxrvk6zyNFxHVj/S0gXiv3BydtAbO0QUir9vgQzwIHBU/WFG4ZhAC2mKznxQeirm4GNvkZU25IR
JLAbl4Rc9RZEssMVgkcleNrfTy7U7uYl3l0zTY8BRvKiftVpGzgX5k/g/WnLm1b0eyFPGdLLt1RE
EkRZ3lGTGY51nCqNFqIMxhRdPGE0LUwuTS+OJeDSc0sR0tUfbB/RLoFkDaHJccqpm5s3xayPhvHP
6+THxPYuZx2F6Lukvv9sczZ7M4/mMIeU3KCe3WSellU0UGCHqqvzXWv/jmydCcgKtfmMeEEt30lM
nSQWamj+Wa2fSpIE6YStz+Tj2zLkb6FTTbvLbDOoAAMlsX3Mc8sl3a/Tph6m2T4RDT4OS9KL3BU/
c0GWYV5Z9uHZazDMcJsc60l4YSnAkx+VWjxXo69OpSo7wFOOK66Er5yYDFpjKDdNmLg+pKc/GxdW
CNqEzmyE/KjrP8ULjaK0c94VtVxMY7TlktJsTmEhjaYaKJpm3+xDzCcxNkf94dM56WDlmCXGOFIf
GA+Ru8IWy6DcMRQ3T6cpmEw7KI2itcV1jlQL+3wej/5mTyCjDOh6FPRO0KXpjHxD2+KPBp1333fL
BFUrweYFoOCRXKkatzXMg0z/RKkau9qiPQOAdXThWNYD00a49CTx0cSHtGAWxQa3OpA8g2U2XLvG
ycQ8gsCkrNPE5RiyeuwmfQfjPhxGHewMoTvjKthAcXTqAYA+nc0OYTUo88rY1Hh/25oVWzhdhMlB
NhNn9IJa8y3YdONNkn8PlGzPDGrbjpUYg/DDjym7ZSGoZM8crEFx5O+qeOVLGXjW6cp4LQOW3hSb
r1AkyTY/MVHTxYIy/LdmOewVpnKVFofK5m9A+fhB3lTZGUtQxU4tKhAhQPPoioUb22w62dZaQDgS
A3IM3Za9PD1W2syn28GyN7fq1IYZ4E3WlHtXdc0HKlkcrzck1qOlGP1RZ3oI84mw9ExtCUAd7b93
YBy6hEWQ1RgWqL4HFgMdYWLgrsCB9gpIAKr7sk7DiHRc6zgaYZQ4zYBEQCwxgrNOGPMfVpLcTtls
BXSU/8EDzP+LsEvfNSvyaWMcLUL55BydfwDAGhDLWtnlu9rB35+dL2FFOr1FxzECcpgIFZPY25m9
nLAOk9AzEM4D3xH5JFOKe3+OgjbwBYDeRaODYkaGPYjEIGRAVpvpfi/RBDeGXVIDhHXxSnUYGN6h
+qCZXQWJix+U408WVUNwC+IZGFzDFXMek0mcktkPOkaSYy+kzzDRhiiacz1RQ499Z5YjQuHW9z5Z
YZpoZzMgggb+63bMuWlKvqOJ77ZSfXNCQHLoAV4LGlBvlu+9fcGUzZfAA1Jd9axFJVhF9likUgos
r//O+jxP69jdilnw2yibSgN3cTTddExVqy9jlDEEWKfVP/KhVBHxDTSIH5MOGoq19VKvb+abUBeu
lfG6+08u90sUVXkprOar5kAOgLSLQ/dT3JM2LTcH+T5DGYjkifeIWCYrSpVkZYoQSZ212Ty4MtzL
eB8CicvmdclnTncKhla1Cl7sapZ5si7THZk5FALg7Vdl0Hifq+49CdVSWwHIPzcXEDNptOrPWcZe
8XVj8Fr9PsM+cjmwSc10M61grYW8rKCzp+OaZCiwzApKeHL6HaS2mG0MOuOLUBsdiB6uncq9TngC
1tMYZ89IZ6zBEksrJYQ4V3aBnuG9GT/1ag0Famu27CkOZY0paU+ta6N1BvGFvGmMOVTAH6r1dPGr
Wc+fpcwqE3Z/WlXlSsGB9zh3Z83CqLnJtSrFYbe1iNy7oGdpo1+uw7lA4qawGWTUztyNhYgio9sa
oXSpPzPvKmCFSEsfYpjF6bYWep2rPTGSMk2ynGKgDN44BqrGdLxLiPhgEOTcmUcE1fUU+wvdC9oQ
uC27Nhp1RDvQetwmFtxu3+jiZIn+ykDrB7ATg0MKMtrvxdhnCPE/NLi045hfYyiFTSdWuKWz2N0M
3bfvcMCDK6WPnRrYGzSsPbJqBU4PaOIb69aTdSIU43l5BZt8rA2YIF9erouXfpPRNkTYKLNWqrRz
FTWiaDS+iSvrwBTXo8PZpadGTUK8Pyr1cRBd9AdSLm4eOZmwVL49LoKMaiIhwbgzAg8O9zsQEuIJ
Jclopud2IZgFwZgcvUgvtZ4Lsj1o4A+LxaA51XsWQOd0t0aLPCsrBSibFdxGCiA2VmeQY2Hz/mPm
uEWClAASsQ9Fk+8k5FGjXSjFXTFKcnru8XqPGgWM+cBkPfNlzK3ReCJ2/f6wsGGlPTyzpj7/bJod
2WDlM23Uj5t/+FmSP3jfgV0XB8cBzLvDHMb+0hTT6onGaou8cOr/iQi6767Mis+2bmIeL+8b5kZo
Npm7snss92mNoBmPiJL21rIwmjp3PrMhzd4Pu7k9t5MfAZpPhsB4rUr++GJnekw5qry00X+vuLbd
Rq3lt6O1PQEZXAslX/lYUZivWRIjZeYaXGg7hCbuNmeuyMXZjUnh+9qlI6CtJaWkUSr/Vrz7ZWz4
DD2BQVJs/Ko9jlI8L8Vj/fwJix9HT2YgRvyuYOtT4SEHOawbLixM9SaD0BHqWfNBaOSOsKCi1aVG
7MdO9BJbCWEtYhBgAWFDKRVbCyFlF9g+4Hao8a6twefHTFsFatfWtCsYiDAhlwzuCaOoTc7vTxPU
+q+j8zgcKXYlKHrDMtrP/7BTIBGOWrAf4fL3hBCtZm7Oc6dqcBZylmpW/t0fDLydG8CwATAL6ays
MD3oGhN8qZ+ZNSLS5jMrbiSdnl3i2oPkuQUxx01bVxPsoyUuObFtmAhER2rkWhzPn+nBDjV3333N
crFLoghU/GUAnyTj9LEDaufZ3O4IxRP/UIaBrk1AL+PhwaVulUdiG9me6Qz5MbExOQxRAcK7smLL
di1RjIrP/iowPRMBfFx1/q9R4n5vQzo8y+exx3+F0etW/aw5hjvY+J1Cyseqpcp+LHxrPRLl5huM
snFN6+SLmiUzu1XAB1Abbf8iyg/Rpvj98oAvmU5iMD4yLCKuv9sw8ZjPhir0Dvm8vfqAvTcxAY8q
V3DK8jipji7cPfxPC9+etgMLCSgqp0ReErcFhkKeQTFn5gRUUOFXK4b9g9b3E69dSg49E/UMg+66
Z8nTml4UJzMVm1AjvM6eYREbAEd5vi6GO2Kql1epYXW2j492flXoFFoiZj0VqqxMcZqXPEi6lHWW
pB8WLfSDoVf30qRYtyQXNE23tKWm0FeaJfbrz52bdMEKFT1gxQ3/mpyBQY26ngsJ5E8OYlbT1r1z
l6ZgrSmU/OWRD/stTivpskRziy3zA1b67D2OCUvpw7lUhzoqPKhOqUUfViPKTusUUtd5dwnmaxe7
j0siS6iLefneKjgIjQ7KMcaADfyhnZFLFqRTYH9DmHR26pl2ivyK/IKKR25Oy4umSXsneSlhRTkQ
8eev+r2QU1m3yKGShyCdBXXtpRd+X8apIWsqtNycbPezYJ70Jokn2+2IFFTgMZdRplNJ0GZi1mvj
hQg8AqPMwFwhjJc5DYN2Kxs3v8bB/R9zaN4ciQXj1UDDXMabaei/9vEp/TyqU/Lbqtx8T2Rf2OBS
B8rUBBFVP3FAmpqUH+vXOjfg6aHOJ3LQk/7Vz6G7GX310sKILXk88PHBoEHHhRFJXielIv1yJ/hU
wumaaYl+Zo9fUWVMOeGOrrSekEQ3NVldJSiwNspHpHM/uFwFty4mLXcookZymB2Tzc9uXKL3BrKx
ReDZ8XUx3DxR4PFXK9hx8bciJa8aLYi9i//aBewEtkwzB66TqQ3mn/3RIDYCzjqjdc7EMZH4e9s/
9z88JKlFyiv4bP3f9limQcomCLoPm2mtmhM3PbN45mLiwfAavrzBhRJbspOUtAMSoxBQLmNyZ7Ze
9jkAjBfZ5OpiglO+FsKsKyc3WyI2VRb58/0MOM0YfOCnWyY678k6CqYwcHKWr4rOVVHmuviihrvg
bne8xJmY9y58i/l6DqcT/kIPkxq93kv7U2dTUAyn00Kvt4RDRQdtMEgwkicxxBafAvH/nYIhhp+2
brUhp22u5nLc5kmS3kIYRKDa52xbU04FhYQWvutU0f9xi8dUhpQ/7anlN+V20iG4mo/bu4FQrkWr
tEVTUAryn4NDNW0BsUVqbtp6yM0DVbljAo/5AFBxhqrEp7ByKHdAKnvAGTBRww+VDlyGZLcuveRj
Dq23uhC1mYYKVd1KFtYpGS6eqY00oSt65DzkoYKZR0yVI5qEFfx6sszIuu83a59jM91JokY1q45k
k4z+o3UZ0B5L82L67fDec8P2ZHK7+DPQxgTP6p8s8CvRhp7hZFO5zWIILBL1d5wEkFvBS26rO7gy
A3iYCt1O4HOFq4yLWUtxpSPBszCb6FeHPrl+I0nPG1R+gPIfFsaLAkvUEpQtRF1RFC6JzY4bobmT
W06myjACtb9FGAcICgW2stcEacJySuTslNIpUDC9dPh1RV/YVDcii8B7/kDvJVZL625iuzMsXbRR
0X9ea1MKhMxeeNtAwPiHnkbzhEyHHKBgQmytKeAku7KfKTz9CSPKdy3zvGbDW41udG2gw74tzSFG
S99jk1Dl88ej9vWv9VbSs0uA24wSIM/lTnq2RmlP99GMXJn2oR3qksIo3XH9YhFKfRf/Eriu0q8m
IAazq2bBDRZAkdasmB0haX8uQhRKp8bW1nGOC86QpYvxJZ69za6/tXOSl5IxjxzBqYvefCLTnyk/
EmNYKoJoJkONssqkc3zsedZlyscgnXUEXFNBFfgnw6NiAeHTDKQfkAqHFKdCoQpSHUvhjoCARNoE
Y4sgksO0u3mgJQP/LLpC9t56jOKZAkuCiKhsD/GxA7TKkeMRzwaViy3XiTyoteDRzLxAU+zM9QLY
X8h3Imc4SmzKMMObxQbj/qTN2QxdsEFdwNRKdJj7Q6yzd0LxxK0tg5LnJDDkqWpCTeuR6zgetCun
lO3jOSvXOXLZcWoA2NPOnyfM1T4vsQssTBYROS9bwEnSwT+A/QOBnHPRX8uV/d9zUsNaxcfSTBAq
ErPCGxuOOo9FFa40b5fYVo+/UIrJmSnw6XtHGNHZySbHfH+n2q0Whzd8LX2CYPUOsQ6uS6vENVOz
7ko1dCm7sUTWXvYFhf1x0QtyFg3jq6NESHjVAPNsWxi8AtiY1YyXh2yo9CdvMuQ7pBp9hY6zZyT6
G0EIG5kslBd+mxSNIbqo8HE/yqikjeWIIyTzqUeTTRC57ZYvIgLf1BVPNqEJufN5H8cXxA3LXpC1
nLUt+Q/W+7eY/J/735HSG3mtLsB80u61SCl5XOiyPuxqgJvSizxRKLW5UACe0bO1QWhJVYbkPKik
GbsxFGFYqRuyU8DbrGF+ENjDrEK4HOzEi8i2d4XV0liB2ZZyorXJQMedJqXnDpwW2D5QH7gsKerL
8MoS/6A6jidmlejCIdWPMckQvt6l4STiiDRZRmyGaNjp+TxSQ/Xam6ejE09Hw+pcK930CABgNvQQ
5bpksnA4h9OArOjPQmRLSuJdPb8pysbY+AC8BSgHVb7X/d+bWvbFf4Zo8fx+43hIsBEK38L1mSpk
B9hlSpmpj21SUodHCFFiuUdGddXlDD4sHrmi436WHLKZQPkWv3IX2cPKLBf9wUDrnQoyCaSXv3wm
73CEyAhlU9GFdt22obRWtlb/HnvwCDF7Z67YKfIg4WD0hPwBhsJyfC31yMGaPX7wyDoeReITXnQy
Ft8eG9USrNbVJAET3GVWKKTccjt8bfDrx9YG/hymMq8E4fmYRHNp3ZZ00tBicIZoiz9TbRfhgeC6
sGd9jszrKugxUdQJLjpYCGq4RhNcVpmce3rGM44PK6D5flguKzu7s4jEPrh95fH/YNo0/PDBe90w
ro5wjhsxduuioB5ye4CUNHI8y4cE4UlgjfgkPcMbd6ScfhL+u2hJRqpZpsxLPu5Eme56RqBd2QlQ
widAZzpeWlGIF0LmxV1Irpjfg1BJROeKl4M3asnhPqRWptcnA7DW/ww9ZKikE0lEFmr1IJAmqDBi
5wXJ4EBerS7cgv2093J3XrjuNp4tyTdSg+hFO2gBLSsmmOjn4laWdVaZWYBVPFX2EBO1JIBauQ6+
7+zKUfVzf/bP4MM0pnFZewX2Bx0/mYJlfwGw19owBdAUVQtcjOU/02wWn2N4DBPgcl+x7Uu3NS5B
87Yk9kGe++pennmu2SldAaVjz840+ierlvrRneJNFEhlEXSrUIuhLArnv9xsZcycEEZcOFoqlNjJ
fNWO0XO/UxYZYtny01B31SxKdszEqCT6h8g4jW+LZuS5M7rdSdS6Pb+r/C0DexZ1NgX9EREzQNyb
FKDl1dU9SlxJP/1Uc2p5CTtMa8XYXajmkKEu+7zZYn+UG5WgVEHfA56O0ykXxi1qw1MlX0Cx3zEc
+Xpvd+53dKz6myz+SL4D6/aEaQWOsXHcYCQz1OCM89wXmNPvZXz+0ZghHk3SK0Xr0goOgfbl1LpN
N2yXU3P2trbjLxqBc1MfAkmGp5uQBG7OEyoXRTM+kxNp5L8Jvq6e/Tr48CYSMQDG6K16Gphq0PRC
WcN7MoLCJznA78T5CE50tO1d/pgf+0wQiXgBT6cwMdoqQ+6uL3Jf2XwP7bUHNBRcJmcMKbUcXtv2
geLgFPdQNjbPMhMnAg8p3VsPh10rItVVS4FuK6EeyJ2QAj9+jm/n+UKxb55NPAF5j5LA68UenDv7
9Bx05xI6PHim+CLYhqoDd75AJpm5BmiFE5f+xDeGShh6sMmrL5CQhqWXed1JjWwitNUt1ukKHGCn
3cR+1ImL0fSXOabSOjY5Lxby35hlGrgO2wQzJni8qzFM1VdyLPSH85Iuu8fDXxQWssAEVElecS4T
pARfUc4gsi+FGlVZP9hyFpvQb/7qmqJO318b/xD2yOdw/jUsmJsE54n2aVCfPKxU14+d1vgm3RnI
AASyAMdu41miMB/KX0mgw/ZN60GsG3NkVC3xKJwAm41ndMScVIrA6hDVUElapZSEPDgZtFYjKSvN
vgXu4Tqb+RiQ7H1TnmTpN1gRsgykt8ITBv+rSlROmMY7kKfBmDRrzciw5ra7w7RqOjGwE4CkG17h
iqI1ZOm9/uT/6CiAlGFQb6AHI9sQ7Gord02swtKWOi6YUf7nUOyf0X/fepH5ovE/k2otcrONqF3m
pMOe15dmWWgNF+cC6owrXH1XkVou+PsE/XfmqBEmKjNZaapORk2n1bYNSqq/5wrUFOdkIyIu2Xhf
gzNIobxb7eS2hWEJ+Re63CS3YX2UdHpwiOPW5BvYnglseF65OtBsQXPHvUS3h8hZbEGFkdpVrVn3
uoUQhsnQXPEaVVAEgzTVOXQa+cFGNiMkQsNcV0LCdhBbtuGT6Jf4lXq1sQG49OaS55xJva/LyJhp
HgzG2U6RYIpRCZkYiVYecccrSvkXRP2zwvDPlPU++43UsB5/fbpsuMq+Dsm1R3hkAgfgYEBvz1lS
fnoPsCDVcwchOc3pjNzb73iyMvrtzGTBwLYF/MKHUfO31LRnhmIfN9wkjSKs77SeRVBdLEU9Rsa/
K+F/1HqTQE5X6IbF8Zj3oxYVYImDF+nDrI81wjEiSZAEYDKb/aWGuXD8VuzlQK8e6OP0LP2vmTn2
GmvueaDjRz1dSZd3sklyDTf7YaEptvHhm1kaU+wK3pbacgJduLKioq46kKu+05yAMnqIBoAzhMw/
uMyU6zNOgNd1B8uOyog2b7kzz0QkDO02PL46ter753Z89aNoE7iQsD45gahDH52kM+91LUIIyvJ2
WyEEoB+V+Kr7obnb2kj9VfP6WQam4z2jLGOL1V4bbALLKuTWkBifiOtyJFP/GHy2YS/QmW4lUzdB
Xqby5ll4uGDQmeJnF3Q23LLyqnKcESftT+voAGa7ILAjbegIaja47OaIHGkQXgtToCcIDYCm4z1r
sowns1bFGZ9Uqg0bHEYeRr5EtaRFjX8DXHH1/fuaxT0lUjpQ/YmHEZTum5l/9GHHrhm7meaReePn
8ECEWdFeLQp0y77KAT6zAh4HNi2/myNnr6+bBoBtKazarsg++F8e1TcTN80CZOiATWPJOeedRIAh
aSomxzBkOzfTqyMZ/WoKCqSucfBVAiCwNX4bL+Mw7mcJ1WLXQdRzrboycR0yng8YF/7FnEaAGCpl
BZUO2+S0qcYQc/2kkebAlVbedq5JawL6FshtyT6l50osaxdms/OJkRTQljuURYM2RQI82E9rSD4Q
humxt75eGT7S9YZep+B0rKcXsGE7K+iMNkgRmaK3/ZnsHxBjPuDWjHaQ1huMg8IgxbSDtzg2dHKJ
RYST/ACBFWMJoI82DxAgpWNYtPnbcRzXW0AhmPhmBfEB25rhAkZoBgItkMJ+iz3Ebf3j5uajM9iv
SNWBQk4UCrTTUWIXk8RZDzHp0dlddvqxEsqU22ifxtrAJixY7qg2xRxlZG/6COsoXwOeijrMft2X
xCasm3eOoKccANQxVC93nuOnhH4ws0cV9y6Rbcplfy7BuT0fllKkfPO8wQw5yRoKbQIt7/yuOv52
NstyjKVcdyPkJDAiFzvGFvJEzsIq+8+KQ5/H8dR962UPQxr6ZJVQ0O06qURVWGV8hst1N6UQtsC2
DxIskAlLzqmL7iN4FeP46b73JFkoTZCX3LF/kvMaHTtk14NAL1WoMhuT8WRjukK6eF8G9z/YnTta
rTVBfpBHdD1Qu6AWM3wpF2JV+EfRs9rDAH3oSWquORwFg1rbvkN61sYjPrGFUVtgnf42sDavU+G2
hp07PvXhS7plR0cLt8crX4ICHyxEeQ39B77e1oK8ZNaLnaOrD7y36dRr9I7iqNZ9qJfJIr36KU3h
xVdYQcxiHFPgqOebw7bT8YUDopQvqUi9nFl4MQjrK8RyWYACFLBIIXy3MUohlZfHmGI/lh5a93lw
dSSC84Jgo0diXrfNXwX8Eda/fQUZgAqMpK1WZm/6mM9dA0VLGGwbzvuPxaN9r/jXqyfJCK3r+Xev
8EtDPyiSf/T3/zmpd24hIUXmfDS30gmMXteKB/UbXBztnf0MD/NIdNmb/5EyfAED2YH7d4a7BHaB
mGF60CZ80FsiDigjmnFl4IDmwjh1h6xOSp+pG0aZNdgktxkNGwSqpPI/sCUtkryqZwQ5vlSKo4K6
nztiKC3tBOm/HIn8bb/PGQzCPl+B/jp4B4mF4+P3/km4W0aTJFk2EKU1rP0jbrgG49VI/RrIiBgy
fvsuxRj10F+VwStLktp4v/YMiE/oeHWW634AwPM56TzjfW6qGtNUa73v4MDNZfeEPdqTjPlkBQ0y
aRMaAr8xXbe+LKwasdI1L3fjfe7NmgX0sNjjdzzWOf/eFs0ABTr9m7/F6wtDbo9I4dainBN3+jGc
AclHj+AcfAtA4hh8h+GQj9iK2BOPrkjLMeboywoaGXDnyYx4uJGIgsMqJIiYfY7ugj+YZTNwyFXo
zLDOsB6WOLsfpij2jhlV4jxZHriU974Tf4zKBfDPi+2E8qTL01byUYuhBV9AzXD1KJXu15aC/DWP
nSolOH3a3TsnwWI+bUnHy8ZRkjaxffzprb5d2ruAvRuJgTQPl+vYcQV6XCwYNiKsSk+QVv3jsW4a
PEaFqLNqGMFbl74xf5OppUbFS4ZFUfA+6h1HyAgUdE+PTbvMCOQ6pDDae7n8oE8RkMO4Bg1JnwtP
xXk66KcsltqgjgMQ0+uprzTcNkmW6cZBz0sLZeudG2jP51JvTwBXIywF0ie6v/7OXC7uLq53YADH
tJs19O8pgQI4hkb63pXv0PolXXDbx1SsrBcw4cfuVwSDRb+8h1lpv/Exjlc6ujCC/78cInRdG1C+
jPhtuwoNGhGJSZTRi/+tdBH7Pu5sraqNesrpx+AfP0a0Md5cGDyFx/xXoQSd31NsSAHmlEkSuk7Q
gkbFbSFUx8oN9Bwt66GRJ0U5vjUesi0BjsrXd65yraNOkfbvOLED05idku38wPjayI4/Im0DxwZf
Wde/sZelpuMmIm6aVPePLjrHvclEji2VLy1OPlatKM1uhsfWztKuMdBRvxevIfZo5kQK5UQ9vUZJ
/4RXpnVZNLS9bm3cB1CbkBMpG5MLwnu8WLHXqo435l9rwqgZv19KDUfBco1BedApmHq2KWl0Bfu3
hACaZO6jEnT/8+fPLmLwMhWmVOI+7fo662E6775kEmg+Ml3DSa/ymB64KWVEKKBq7FP8h1qBAGzr
IoN5O0BYZQkvBHaD086ct+9cs13RDUTkiNAH3gXgYpqz8JBctS+WEXgN9TRjUAJT7EscR0o6UYt2
kZEkYvsXMuklaF8qRSO6thZIfVh4rlwJAbWmQV6gpFoV2KZVbvZokm16bU2CLHX03rFmCV+HvPYh
6+NbkC0J22dOTJborKqLdU8GF8l/yrNmgSaw/qjGu0rJuF0vymgqkzowBlM9/EHBAm9KZGQl2VX+
ApQUV3wpGvCSAfM0k3eADCOf5jeHvKgs8KGuGPPoBJJboLcysryax/SAm3DkkUdK/83el7FWfbVI
p67xaYfMXfa096YNSnFfl+++f7NDfu2UrEqMAZN767bsKwtN61DMGCjvyhRRLlZ3PLWxBiEl9Mj5
qPDsDTxT4GK6JP+re8zVyMNVlRz6u4pFKRq1G+l8J5L35Lvj9xc+7/OCBoYKb0FScQWbNyPbtFxy
25Bz3fnjrrLdG+eylH+YV8Vl1zSZpjATQb2SBdUjGcqRi8YKzh++qjmY0tQEo2Y962o9yjfn0K5U
UYb11SiFS1Hxm39URKx4YstsZ/IIo27wUy9hAoM5uhEznw4T0AQzEwRsMgbgdqbx+lEwSFYQLpqf
kyF2WmDBWsqqM7S886RC1+BTxT4meiMOObQqMSnp6t+dih3HibdIGEuak32U188iErBiOzCIk5Ha
xlh7qJ8DyAtaDs7Igo9yFRh7w1W9r2ptXSU86iS/UXpeY9R2KEnjc0R5w3Z9bwDPHIEBarPMZaBl
hMAH+B9Gdk4SI5DtoF4hIabYYCtcDQt0jXbEJPeYFM6KS+H3f6mlKhoDp+Rzf0qSy/I9+H5AZX4L
ehSJiPkIVfxgOTeAijOl+EA4g3fdwDN+rur/4hmyQBkgVAb66R8C51Rb4J98hL0wiL54qAbkBRuL
c5KxwkPUTSjTCoxWQgib+TJedNUSqttmGcEq/vEikdjOubWyfWUBUZNBTAH53IEQuNU1xCAXdbZp
LRqRbh2RnMfFEMGbejqCpzeA1B4Lkian01sOMFvC0pc+D5G7ACMHIMqjo9cItH6u2UOj5Qsbx65W
hOe1llQaK1X8/9BIMzIi3SzuK0NuWue3rmN3tw7QeeSTZq3dE2A4obDmDea20458CpZs1TJHbSpx
ksn43+wHHpJqSo8AWy8e6WPzdfZZORCknCU/RHpCVFWsMrTop251oTp1vP9djJ+h6ZxeZva+rj9L
7Jvzv0Lzi4ZMIEUN7JqUHKPiay8Z90Qg1n2upJOzOadxPyipQ4/mO+JAEL5mm515cf85GsOLEmSM
OCGEIMqP0luEEf/jSn4iTTIAscAYB0CvbKswn4JtzzdY0JTCU+Aj2VR2Ag3QfTeE2ZMO/DdFZ1k2
961xGUzCC0ekzCddkqPYnZj4LO1cqSKQBp9Qlu6m7EmEioOPQdChFJksQi8rUBPscNBb28Qo9lPo
8333keBtotCJHgHXK/qsL81ecFgVjVZFF2HOY9+8+T+LOPNSxxlZ5/E1OV5z7wJC+FNOEQcf6ZT5
PohurcUGq3X65l++6kqxvsU13fd5M1VcuiIoPBIDayra0mrC7Fcz5vINNs5d2GYt5/lG48NKTJMv
w6rwGH2jPSxmv0usy/TKb9Vj2VL9fuTmrsruGoTRAfN9ykY4hQDqgnBTbNLg5TAU6KUM7DTOncQv
yLnfWjSNHuPxRugNG3UuPhBV7BPwrk8ZjokU19XMWIXoRSLbmBRg9W+NqsMh6+BmL7Q9DEu75rGh
/1YcNTwPeNsWSibaZlZOPFtoiYY6CgD83BxJf3piJOr6kryEV9AAheZ4Ab6B0x/qiKsvxg9MPda9
hhHNywwUA3bb9u4XmRIJmipjJV+Cc59qhYAw6b8loC2yaCv8jbqaPKDDELHJHyIpEdSRBYOIUTQR
0hzdpB/Hox6LiAvsP+su4t23xBmP0BXnm3TAytc/BtGesl9yaYN+mQdYOydqHZM8xciPeuXALhbA
HDfWah0PrzyTi/F5NmP028bVt2d6UfyQqBuM74YTQrBZ3WE27IH05Tm2ndQ6q2v8xIP24e6rkXMc
hy9L7YVHHWaCD190h84qYpHjLecAzw5MMJNjGsEOOEy7KZ35V6z4YFhdT53XRVwrYbdj1ej6iuoS
pAI8GjBHBhZh4uZdR32E/QYlneD+kCqCmGf1FZrn8pyhtdcfN+J9iTMP3YXT8s44eXuHh61rs2Ke
wzL0O7cV+MUKdI1KZLAens5XUcmV6NlmQEDrjMNqF21PLokSdv6IaeKiFLEsx6ooGxRsVu1wMfdw
gyTNrnSEWG7PZGEbhS/BtMqVqjOR2jlNUpnzzl7TwN+t87dSitUmPOY6Q2T4cGSH5Q9rRcCRC/Jy
uiAMy5gdWK5gfCnSyPYE6EAEJkFTRwR0AVARXoD64Qrtecg3mVoBhg23Rm1d+wQolC7hicfAJj28
Jr5jkv+rUHxLoJKTFnx5wyhRau4xhZ9OpEyWDtnuv5/WRy73RoO0LawGOatiP+bkrIeL6Ut8bntH
j3mZSXeVwgBrlicBXHM4jLPieqMtPIptvgg8SzalmhSLhPDkHRCfMI0Tm+bMVegOQUnYtfwOv5M+
GVQkpQ4PRAohuheHxpUVO9RWuS+jadJbCJk2xhiRMcmyCqT1o+/ivrd36SBw+8TrQ3HYi2Uw+Zjn
yrDdCMT+1asJQjh+EpYyr1ftYL7zHsuEEsAXtoy34zt/az594Ew6t/2a6eF+t1MFWtDsnn6WwQMK
lZ5OSB6nrDqYFUAN+nyc+1fFj5NQXrJ0Ip5iEcx1mQvCBxZ4yrwInaplYFSvtdo/nxiJqOVaHZFO
T0S4QxW+8N/5rmnECt0nurcA3Pc3wq7rsjRcuJpIBKg2qkyF7wXIXORAHin4L1mErZ13psLxP6+d
j5VeBFuo0lLZ2n/JY6LKyyk7PbadRajczhqwqxEKXUq1vYm5QxbDkzTSeIjv6QIKIktzYHXBQcIs
kinlEId4rPVuN8hjUi83d9EpsTaegChlenrDrmF/PoA9blOazKOb5YSirVXI97XczoxQFl1/4R2h
QZvhg6cBg9eb3cdGM/59jOi0VlcTYdjYwUnKhFRk1lrDaHR534lHBg0Wx8P4om3Ej41i8CnL8woA
9E3ZJjtjdfR+yAS+0vX8R6Bq2iD5uH2O+CXfbCiX6o5VwT0hvcnN5QyN4Fze+XS+Rw4pWyG0laX6
qK/sMuiTX8bW+sCfopY/B4B4cLmH/quCxz4UWSFmNFRj9T/94RJdXz5o6iYjCFg32mT7HFBctKFc
6pKh+PzbqciDElFxJqXSHaubwclCJpmeT7oMjksCdOTobpc7Mf7g07b+x6KCDtsbaJCrmown0SCL
YDqn/HQuvKKXgQH0wBCuvt2P7WkjG7omg3zBB5sefsnwCv10XMxuoFX4BXR30No90KSux1LPaFH7
U0PpR5lOn6XMCrmyTxKfPSxg6NDfwuRZ+MrpQBvPnU3JJJdl/woAaFLI8yo26bX4RWx40IJB6uWR
nc9XHwvDvalWX0hdMPPbKfj1M/4tXir7dLX+QkpGIZQqnHqmwvyyk47WjZu/YTOCDvj2OizKbmHv
wRDyhQje4cN5cUokmNLuhzAdpOmt5kTX+NC+nSNSmC6hQSWYEEp/F+haZtgAyLyNo5QWXpiFXqaR
eU4by2MmXP4SxETPGIqcbCnocSS5ZgZ5EU8fydV88zadiK3RhKg8ugHFEslbc6WdyFAa5DQykGfn
6xEprtAELZnDhdV5jtO4a454rtICMefCc9xj4VwBsZsxw4YAcnqastMspRQhHq00EjXghpYZw1G+
wNDn83okcFN0BJfiDZKO1VgT1IbWMsfyCv+MtXFWNTnw0mZQR/KrBYUTKrxFEjl43sTNdLaiysZy
oLwJ3QLFJPFaQ0yNr0g+auadleJbmlK1bwEH5QnA16ZKZmNQkWDIHNkZwYeoH+WPt5lYlvcaNH4s
1QqOLpbIff771J26M1WE6MBqawRGazM7LNx9vpX6UtRAc5ceBwrNfqjizQ6Fxp/CaalgKlag5COI
NaifqNFUkBzAqNjR4cy8vSi4QCSFff35a+QAcAu+kmLrqTkFDJOCvQA3W0ggSyqhbBgHxzvYajY6
0rnrzEq5NQKsZsAQwLHDL2jYP5c6MNVwUUGeucwZGrOkt5Fc6bFGUhh6/iyhF35n29B3wFo9ejKS
KtXQb/sGkKtvglBTSLMqL+jwl4ca2DixvVZRPI1BEtZKMtDD8ao9g3Sy5KEkVQ939HzrmFsqVLfC
RXPqUlyWiXKUWS6gGvgsejpsqGP/7hbzFO7664AS0hEsUnh4fckWmS+B1jHqFDSd/wSUIbT2wkwg
LxYlV4nfRCrs4avxG1kSuePUSgsFJbr79S5Fq+tcHwp8/KIhViphC90xb0nOWJprjeJIUpTeziK2
BTOKnOoiiHZJ03IAlCFj0ER6hhYWOF59kvIxLz+240Xecz6CzILu9/+tuo4g15oD8EhpOq5NvMSQ
IbmrbxnsDsZXNhOuLJVPX7r9WP4mwRGGVWXEs7ANOnjrtKKdqS6+0hj0xwFzyfWXcCQIwwlIWGBT
r/hz46rni0atGtjC1SD1FwyScrUWCnTv+WYL6jyqOTnvMO3KK83jXQxcjCv1kP4rW8aVGBhMKTwX
kJy64hJfs/fGESJBxyFExE4wzJ8d1YkDX32cQGhAKZIdCP9zQRKciw/vdBlcRNCBxFujntwRB7zq
+WNYVSOBNRF1K29AuiAqA4K4AXQJKA0hdwfDD9YXuqPkfftZ5+caKOkEw8U1XcRy5HZld+UCi+pS
obfN0dPIov5ogratM0U05KgtEcCwguALto6fx9c3o9YiHG7G3Ugd7bUpP+U46UXcMObMfqfFX+CN
iJgl4Y5ULHSi7VDmmwoL96HG38ouLxD37Up+HkLsdm+OOikEytDV5kBw+DjaF7UBHEM0lzrRwJik
kddbNGcwfd5woUusqRlRl8H2DKYg+/3h2Wem9RFo8Ot2irlQ/wzrimA/AADooCGX18W3P7a6ryWv
xiDjPEBgrgwVNnerk0jYKM49nHPtS5QEJ4AMntONtEbl6DMl74AaQ/Brscd9++o7KjLjGj0zPzBw
MSneaSFs2UKYlAi+bUlx8y0DpzkGa+fU7vm/PTIuYALHDzVTSbRvBC1HM/QQOm4fFmZtZoPDQ4ZG
638hlojKTRqPJ8MXsJZz1lvB2BtiFd2oEPXu3RPRysdvjtu0/4PNbEgjx3jVnt3iqTKDIoM0BaCY
PzV/cYNqRic1OkugKauMrhPgmAN6rvcW5vLAyAUUmhQxNQCJU5tHhQobWtZAY8bMtCtgDAJ7c7bU
QhL9k28m7l+rYCzu5D67pi7FTnHL9ZJ7HUgiTR975+w3dvnp2+DFECjO1eTdKzt76D6a1bMy0g1K
o0fJ/Efy1XaDUEF2qGjNmm0xAC2VU3q9dOZHWTiD9dPDppDMBIbL1LfjoPnE44DJFE5MP9ha4hT5
0UlpM8O3V9+soNubQ6F1Xi7hvOuMnuR8cMo4Z/qspWy/4xHHIiqlrf5HDyUt6enorhvzaq1xC5uZ
5KVHbWAmAs6c4xItJZpRYkwfkvbL/sXrJMCMwozBNrYEvvyAEhMlFxTvpfTvyS2OB74xct8bmAl4
x2R3aJDtQKPAgdEbCQ9yFkNo0pxbKtIWaB/jpg/l4RKcgEk7xsjAJAZom2iyWSGkIcBLDBDOSJS8
bpOf7dEcJXoCabuJ++nVL1VTGxm2RtVBr3yuCdvZf67pBxriRoKvCQ70Ovet4NFMUh4qTiUdeouM
dd4V2n+wfC4xEDRPpQWBFBC6B9SXC4TbgrH3anmi8SgwO/hOl1TLWLGjFdHcnRcZHMx4uEfb5STA
UHc+bNIfkJoS4PBW6EAQ5yi6RgHKlRmCK43TRYOg8M4frmmyXxy86u7sq42APfsK+hnuEh35ym7A
jN7QbUFwCojOZ3R1kNFR5bZlzDz6KMKVL9ayevU+KLOTfqx8P6NfKnmXZzAXqg+L1WzuhFb2EnsR
d3VDaIiucZAbviln7xD3/61fJl2KL6cXEm4EUe12FiZus/az6oOOVhRc5jB8J+C/6LpxOi9c7Bv4
rF2lfq7OHbkRv/KOyddjYD/Trvpp3q9rE8dx0Sc6EI9S81k+jjNnfSwZkPA9+WTIWXSL4vdxt2Xg
BcYiWfKzoMT4BFU7u/JRR/ykgVG8xNENzkuReIzllW1frxci61TcRKX83QAgPvR/Zn3/RTd5ScwN
ehKRMblsZrvYILBIqK7BhYPPhqVSmWXZLJn9V62may5Y4KIZHdukzRyPIwDYXDsdwtamsjnsUTCu
I2pkFfzn63E7a7b3CCAyvHxF7dmEj0vAqh79HLPhVHABED7f4N01K96AlW3mRqC9OhBln4ZkGytF
MeEglQwgJIPh4WbLgRxF1A0wJo1CEeFbgJG+wFybgpEKslevNteXD8jK4mgDZTu9AIU5JlJWay22
k3V7kWXT7xUTfFav4Ciu5JIqGHzdCqInSSxfaMmG0IgxXmFVyMbLo2YBPULSfS2v299XOQeKZvLF
XZkwAcKMHY5KS8XzZdfDZHWW3lY7nNnv4nvZbnCgVBUCQdJYxuYuv19bfxW/mWhkjVNakpO7BwXg
0vhVbb7d+GcHCV3c8WXEyTordqzYQIPW1X1Of1gZ177Q0GdcS7moPUfK/PVKWLiyXoGonv0DqLN5
xhB0zmUT3x7rlmY/1rti4cfwvS8uT4pdIZlMcdGUJ9Mwg+8J7eEAyGbrzxtI/ZudpJWDMjpuryfh
68AAAprKV+i/siYC0k9jIwWqmIXFEr4ZtndXf8Ry3ca0F+y40aBASGiv7w5HD4/R+jq/UMmaZfwQ
BdUqrj1jnpWNpT6jm9yb7WLJHlHtgywUzf8XQbme2ijj0zXuuWFPtRv2Sx2HLmmGsZotKUNQ1x22
hiUrcqnNVqhlGUGGWdqlLquFu6nIJjmwFrjEiUxZqOKYvoaC54YDAfrTnrPW3OMgY/H1/SuhTyR6
53ZtJOEYXMAtitkWCzVI8xOAoYS5mm7UYFzHWp961+K61Oi6cFb8k6+IxJteVmYKGcI2ZkF8jekt
q8rUBCLJnC/+6e9MUYzMRddun73jcGWN2UaIw9oAPvb7WWiDtkygEmXlIgZH4SpPMHBaVd78uTfB
YguqCkrxvEu6Jh2spDyqUyhncF03HaH4aqTzWzcPl6oRJBFnp1fC+CUsDJcwZL1/scoXHekonsV7
iDkVzqBH8wuMnvcXVOt+CjUQC83q7J8XVKjppKAKe/COznLuTPVEDMoCrOBJHOR/CRh+ITENHsP1
kkSilW6vucKtgaiQPfNDGkH8g/eTcJkGPCLA+N/X1iE3hpQftaZXvqkEBT6rU3sa69nbk/cU3l5J
xbBNxY9LOiqSeWFMG4t8A0P6MDpKUP1FABd7N+FA9hQih8VKCVKlZEcNijh4yRZzhTGnLdt/NoDL
N4K1V01zqFnxM4dwNMlcd7/SrXhgRFY4tmVQuzFJMt8W+v5QMMXV2PUzmnt/OPAznNizlKYP+G6B
kYLkM0sWXBo1iSJPW/fPs8HVM8YyoKZLreCUl6USjcCFkUq5UPUE5IElMfwzmPQvRih3c6ZW/jsu
VcqboWUUVLyb2PTZhtRS97J/qQRBWXFNDW5Ak3Yz+xDUUYQtQlwAqtZUue4nrUA8mn1FHor5qh43
vP20aKQgY9VTReS8SbHzqtywEJPQOoXpOtKVxPS6iiuosfB70hsNH4xCxSTfaZp1Ezyeuv4D9lKX
Ewl7oIyHg0bvVVreftSOvaGF3U3g4a2Q7/SbmYCTIYqz96rMYs2OvxTRug4v2gJ1EOikOqGxemSB
H2HSRfFQW4XdghvXCv8wHbWVOFSWO2wmUYMn58TrZdAB7GWiFQdZWJi/Ul7LzySxw7QHzv3PEMG7
1PmkRMbeg0O4ZOBRVqnuOtamTYRlgensgUB3LwO0P7nXP2GR/qOEtu9jzZRqzTfLVISufgW/QwNe
1a94R5BsgSoA4eczW2khYrbfCCcZJcwwlR9exqhegja2/oMboeXAdR9f54nVJ0Upgh5LXGgarlr3
ZrgQbjXiVeUmLD/5bWoba8FC8LS7UJ9crDvIir8n4suzrwtGcpbXabDtiFA94lZxox0AuHbH5p9R
FFEEUi3kxKPWNW3SNcgdHmjqKqVUkraqo9SuEtUe2iUwep+QA+yIfdbn6CDdQKaN3I/p/0mhikuB
3HLY+b2hG/F6iNAomh60lFsdGG+Qfcc/L9YbdaCDGb8w9bi8iuaKa8Tgu9lQJ04vimSNG5R9AFS/
gblneFQNNlgOJPGgFxAU5S2MJBqb0fD0Hd4yd0zRprZbTtIsrJsMwQKPr5UNSkm2ARpWH6m5k0Lc
iPD7dcXZp8+nGfoUP/0bFWqufLQ/j1NPmV++LTtNEmRYJB1pulc9zroWEQbPO+lE/0p+lmu0vv0W
j3FizsfIOeJ2P9TkVBVvehKkYTbtDyRMh9Ltp+Tmyd6fUDj2LAvCSegPgQL4y1IAmhgftmJtUWXy
AtK76eksMq+4W99DBogj0Saz6LWtVWSWVGwYcMAZRvmkQ+cEAOkibz1zDKA/psujJE90jBi57Gwq
z4RVZurj5W3QZtWyT3alfnxLa+rHe0RJLZZuRyDWqjKH5/4Kk+2kyGgOhM7THBq/zlwRXf9oLgKT
w/0GDQRHNaFJ0tG10/aK1CcqofeGaf1k9ff4/ZHeMLCCZGDM6V+DIvgGy57KB3s8RRnrYCuP05wr
Z10KdDpUdla54oU2IGpc/T+1Ccn73CkXLbpRdxSCNLNmdQocbRtP5+HclzCtB7YqSgjxDt5XkMEX
VR0mpqz+3tNhBwfxSjuPOA9172dH4zeSp89R1mVLjLr9RXx1RE7S3oK521E3spB0HrmzmHhpg3KL
gFWf89m6w/8ScxsA+xX1SVMM8//RRNmpMlit4jCgBCEB/dwAk8n8283opVX6iYJ/GOIQtahh+KD6
snXB+9eeFmuGoNiCnw+NMvqxI8eSRAQcXRRHf5t73fLEtfAZl13NJ3DX7gbiSlfYMP4yPzQTmACi
W+389UrDoPseLzZOwN/aDvYzDMuliIl6TGD3pWGrJrOttyu3dQ67yrvhAdngcoRqQgHTuBgU3vJW
gCLHLZ0XsSvklGcrg0r7314COggepbQa6mCCUS34JMKAYE8D/SOs1LEvbdgntHP2nuZzdFYPBcTz
NTVboYAMTFMV9l8bOjw13UMNKrrDfJ+UIwA7dxb8CVWAhWPx12HUwVcZCJ3LeAXWv7Y5rinqGWcE
lj1uuv5sfBeosBgZgnNSR8becQVUO7SQNmFVLzwqz0f/O6iqzv3Er/3RIXlwJGzwld+vZ/hrwfpO
NHjufq7T0mRRTxKQZNEp45reUygYvXUGOL9JcJ4kAVf0WzgKW2T2u4Qu+s3u8ElcRWAoN7vTtq8x
Wp+sErJq8rQnSO/lzaf4a0+LbuJW4rDpOOTr0vtbH+cWqUfFJo8VsPxdnM5QFGR3+JcAaSbJIyS2
ZptdLjDPaR8dW0+1a4/3l2+viQAHZOAPecdQr2SrENFs1Prcy85HmCO7aBpZCtXpx7FoCVU09oI6
Tg80yVebPRcLQCtEaRaGHGZUzajTz/HL+zxE0KIpRMUHtlm4YcLVw5XdtFw77J6avXb+TAWPq6o/
Ep5ZgbiHaY0ZHkmFwrSwGeEGHB0SGePuzuqNShdrBpyxa/0iUmlQl0yswnbuxUSU61Vqf1x9qQ+N
0kIi+GmJ4+xPp5DQxa26XSvpOLG7E49nQkHDgYevAGLcvnsXnKhDqVD5tBRBy3NJXbXzLhuT74Ux
T7dgSB+CQHG5KL1Krnvuk+Fjn9aL5l7pMPlOTKQl+VyCb6frHqSJv5s+E/62K8JlGbUXTW4vHf92
cNWaO9D4vtTqhtQqaq4YjkikUDdKE18pJpTINIumHl1UREkRIunGrWAYLy0ILywHu3k0gEW+ELkZ
o74FYI3INwSaZ/wVQwugYMA86gcHbPCIAeC8N4U2uL+M+YjrpRVSjn4BKX9YwUfhaOScv+Q1o2y2
VKZn2xebg1YYgDg+AsoClDn5eO9jMLGy2sIeqdwHGCy4UqtXvp/IK3JV/4biQoUniCNoAMlhMIih
PYDyKeb+skAcRxLxV2nuWmVvPR0g+2ryeNEzJv85c/zSTJZ5AKGvG+1Vo+IF1ZmMklmkjDhT8T/g
wMYl1u2LytfkBc1dOiRaP6PwiVNspK5/DkjBzE115P/CjVafRdfQQXAo64RJXK3LrQO7hCDM6WuL
7qCnOIBTQ/NcK3mKYOlfgP19Ebj4XuqrkAoBLDVJjznZv1e7xSpS6hU+fk4SiYevVifnS/xIYxFV
28ybyPlrd1/kcN7s5rXUsQFmN7x1C8bVIscfSBYW0nuGF4Xheucw5NVm3+AmQBYCK29FzUfO0Sn8
MDSxjQJJf0WH0iERuJJMkx3JEU74myCn2VVKnU+yHebZHaiAnH3ov8OidIKygOzDakxhIQ+VoMNf
4JYuGat0YoLdFTZz8411d/uO44kRh3IQiMfdawIcFd+iGcQ+/0aQb6ddmiMPmI2QuTyKrGWkQgot
WQRkwmRuWJw4G8J2kWL+BJa6nkmyfjINeDisRWzJP1jUA9l4c7KH93HOz6UquSxbtem+xHzMS+/H
B448cCWaXlYCs4lBeuq5WMONlRcTKjA+tdxOiJ9Ad+ikYa3tPWJZs0+RCekia+ktWm3zWNSiiGpC
MwUJHmby8jzRYRB+KihL8+G0cZb5KaR5ybGR+XCn1vn9PK8thK6RNP6ETau5QODtogqkhjHgF67U
p0slwKp0c+xR4PfGaM2lYsQBFu2mpR8SQ/KrdagXYXkpYUqKMfxvPY7o0pDpMYoO2Wim3OlxjQE1
XmDlJL4nYnLPpYBF8wSw+sZPvdGFcV0fpvxEMhT21Nvb4pUgEbcbfN58BksYiB/FXkskO7cfUGEN
tONSGeYpo6jcSj6QY8tSO2OSaRsnhTUxDJezG7IC6KKbpkBR2EAmMIi0dgax0X4QdlZRnBWbWj51
aNslIyL/R+mdPf/VxtpAzQVSnBeR8v+8BMDtWxWCf3MUo0v+GMSUijRcpFEfwMAnssvKnyV2z2kY
XUIM4s5LCcIWgIfpGoyUErCcO2s1OqN5B4s6QRwnCDFobIdPhSdqU5M4lPuIju4KfH6yg5TKeaOX
KwiDHVUQjbaGrmllNZCniiOtYzmMUg9gCwTfL8anSvlyzVeTJbhqgm4bRu5W8drzzTPh2fqjSL9Q
RvwICij3b0WL19GzxEUSeFISJ0QFsygjS1qRb8XXfu6As00iyMCSU2zquRJ8SdDMVY/Ug8Df3+MI
y2YlNNNdJUyceS7OWVVS9E3mncChb76oasr2x1/KCh7tZ3h7O3dFrJ3aK2erW0nkd3o7fXzafwTX
6E1yNL6GN3fVrdMg35RLEPdB4YXFPnrNbGlqIcg7hC0CcGGmP6px4Sezrx03k6qn6iN52vt5/+bv
oc2N8ig61gdwukK+XWI3TuspETvTvhAo6Zp4hov8zMZAsOxvz/yZ/G6iqRe/Cd2Q9/NQ6Kt2FjRc
Ohb1msaf2TRCMB0CmdskQizF0t8SMPrW/bM45KJPnrufYo2xKiTprlcxy0mqx0vXZ1OwPy+N6FmE
3MB9GPuMMxKvtivnx6oBZX4SZPiz8rHjwbhvGmAy2d3oKO0rtvukONz77x2dYSSSaNI4EA41Z2kF
jRzPU0AV46j/94rc2lG1W8M0Fe480SEAz6OgVOo7Z4EMPYBLPEUmMiwzCD/qJkQLQW2pDw/5uiN3
TsG7YMs/2IYQxxX9By87X36IhGX8iFqllcOd52xhZ1Xhr9R1gVSbJYSJtotB6GXH5PvWex06f3TX
eitnhtQnJW+pxpD4Nh4uGvwQAwLYdHj7CspmINmrirPRTAshav3rkRtLxiy/QJ634mbG9XNKYKfK
QSobGmKmJUCQGkIxbXIISAt6yhhncZhvEaZxDZIyFtkBt+pfAZNM1L0wifdCKPTkOEJ8/WtlMzNK
LdD8bqejrsxuLvDxWMCgxnLfKS2GdnhHYgZUD9+b8WOYbC0wbC8JLI4uNqFdcoAgj45c3etanEto
z2bS0LsMTHQigOhqacYgZ7DrA1N/tgKrcaio02KOCmR3p7T4SqJt1Ejk4nC43RkCV38txkZJ7qfg
XIV+ncHxHJIgsmRmR7ZnLzl+Ut/otkPFBTgaIHFokfBEriWIrC/DH2JP6qOuY3BYN7Vm/Uhbit6s
BcYaRH25wqEjrW4pcsXVAFkFfQzQXfrjTwFB3GVl6ca1mw3NTpo4r2xboDv1aJgV0hDQ5JOiPF2F
/yS2+QCvYq/9+qAMBeBiRivjyvCDfXDMwFRCeHrjrBZQ9u1cBAd1SL2IQCZfd1EwWO6sqzeAR4Uz
zw5cxaI+0nXw+jkG3ksYOIQjXGz735quAXKjgZbzpiFiMyTA6gCeuTzVImExSqOkqrMBAQKGeDFD
lYJyXs1bXp801hlVvuZXpkmzJq9IoNUml6RtlyWI0lZWgB4Dohifhh1aGaINRHAqMKlJfeg03ty6
ldJBggiKfcr+NA9wI/sgszGRupDIw2zsLuO8yGOb+vKzC8/FRdtJ5d/rBpRFUrvnL+YCPZMk5Tft
Q9SsNoBb457U7a3WCag8tOebBwQHfO5TWMaOaMzdOsLCo1JObW1DF8bmPCdk2/Wwc2RRN5E1J8hF
57YGozoQWfi54m/5XHhILECkW79NIHOAquPZ7aT3Ol+rbAmlBWHU1prE2n/H0Eaymc0GgjPekXXP
auYjr8dwq9g6lSkNhcgnclDdnnStOrrVdN5oUo0q5cn3gPKuX0GVRoN1+ZsDwXNnfovEGH4cA2RR
/HTzNYBt6kIv8PvH1tZBA4Wpww3J9D5E05E1EEVrjm1/OAlGGUjFu+clE27pig5qjnF+3ZTyoznG
xdfgvhxyQZRYb/b9oQx0b/n8p8BdPA20tbz6qYZ1zei8IWAC0YDAmy/VdPDqcDx8LhvrwNE7wWsd
UTJcU/AKCNMruUP60lqQXqbrsrtkOcRIhgthYLcjtLHKofuvtAIIj36C/Bz+t34KBaOdPuSOKFQL
jo+/hnP0y9/kElTo4DFtOgZubnJppk0DO1/LJ4zmmvfybSXFBcAOGSpAjz/IG12VRbiPCdwDFWzd
lz8vE8PqOMMOw7F9lbyH9Pa7N5dQF7+x/CZwCFn76Hs2dlQBVmd1QlKP8Y1Dm15xYXRW76FX+yBb
d0Od83YLRFBRAE3hOkLzWsBuLZU1ew/CiXcWLq4OOic8X59V/W7MecJuMIZW4LtAV7WRAmMvSNyq
mPDLcOiunRXN0e/Z7IfTA2Aok+EAFWKcY3mm1JSrltxyMCd4hIAZTzOeRjIvtEha7+dPym4zzS3T
oj0Or6b//5erZyPK2Z0PjTXMWOJy9xZel+g8FxZxyRoHIbtP+MlKOIO7s5WKyaFCaFMvDSSgzkIf
/Z2Pc1ZZ5sM8aNiCTNGrR+GTdDxY1VC9VX1FhomDi1awEhrdSCKhY9es7UTIjNN00Ismt3vJ1pDM
ZETXgpBe/uHPFiZdr01c2kQvjVacfimQ5T3JtLPWwXIxqlGh6lwYlvoc30gMuvWel94Yrd67nh2l
WPZdQnyIkZ6emoFxaYFhjAx+SEoqqewqZcTT5xE5LWOg2CXVrNouoTv5HbPW7oz1xb5/4r+zbndy
AR0Sq3z5XA0tWafwOrsRh7sz0TUILb4+3b3HOvmaVCsjsc1PS6meJZQufJXYNwdaeiIS73/vtLrk
sy3PhtLuKHf1Dj0AoQ/Oj535hhJzgxx3djsYoeoGS5UEBb3bIIYV0ELv6xdu2k3SZXXJFjkoVOjh
6sju3xux7BzlQ/m2lgVdCTc0eekU0Um5aoS+MSLJrBbez2CqNXp07gvbolq9qR/cyk3nigI0wQHN
POW4xt46oa0bg2+MJ6ppXBHQA6IyG3aCbOKrfNBjNrIhf9480tDCnRSwxsEgeT4OLyQKtg6BVgQp
r6cO3ot5m6WGfZjdCYgKBenF0quVOn1fAFZFFEfbZktRMFl7CQ3GeWt1J+V1eUsfSEIe2tf5B4M8
HWZHtY6q8yifUdKY53Pi1xlI1MxSECtyrjMGtA61oP44lh2/RuEWW8lqUt6NxCZe3hALdXU4AcLG
OzxI1pi/oGJUQMbuQ5tYz5Y3pjyV0WE5DEWUfwbCKEOURE+NSiWxeicmN7JshN5Qsk7mWqLnzDvr
Pi8dUAvg9hg3EJW88bFJDJZdEz31TlLAZH636vBVjFAamZvUeFZHr5HVBX5wa9bPH2xCCmYln3fe
6sqiokWNHeRsv3QyckbjQIfHL5y9Gl0Hvz9ORfiVLfw2QpBJ22fxCQpVQKSDwydP8kDxU0kvJ4d9
WXHrRTI+xe/pux2hgaFAgKAG56fdq+TiZKa2rIShdgJkfsIxD+mvNm6FoOXuG9oI7nQ8XkrVAnLl
OksnmNpG8KB/2vMCa1XFO8WCsqr7O6HbFW7UNA+MoGdtAVvhupVZNdVVWfQ0Cj/bhjIyYZYwj8ej
KzomwgOagcyzryaVa7vvJjMbXUW6sir0OJQzGAOpjFmP6aAIeU2MWvwqhQ9R453FBUYWWCaFQN7G
B+nGXNwFMDimGFGdp9Oh0Ua2Wylh16Xe0ari+9A8NwDEy8vYPN3WrG7LDLFCHT5Ahp9ZN645BD6H
UtiEQqG3axxQAQlZZbLKWzr8lJcwLsDAst3Kt07sl+kov+tHLEpCX7JoUy1FG7l4750nS835klsX
zY69qCAFe0a1LhJ3TUKKhTkO32r2t2fhRQXfV5uhPxlfg9o7XZJ3s6z61v4lqiE2m07UxIoJfCTD
33RgN3Kfy11U+tJ6pHRd15ScnP8VQsjXIa+9WTiZmctX0oGFJ2D5GpavvkvGfkl+P5ONPQ5nYtRR
FVubYSxCKi5jPVHyXcjvp7NleRfQJoJ4hW9q+JAui2cK7rKJsQoCH5awTv73UTdnRTfXqluY6Kqn
Z5S8lvNhhYiAlO89LnpKeLwsvrwkzUNXdBDXV2b1+d9IoIxv4CH7lJkneHrT/9fIoURU4wbY0++U
FemUsl2E0SJTNogGUg0EdlDjzuzXGRoGUca+MCZ5IcZWiav1mtnmdPuMKtWYbkXVVN19YjaxMj1o
JBl7p/o1czqSvLQoxYloA8bKr0jScZhtkrHRGoBF1xjVDBQJfTaVnX/1DYhT6B2p7RNjjToKGrgX
PcivyanWieVlh+EmXCPk/2UsLpoBbOuSBUNURCVZ5/EXtb1Bl/Hu1RV0dEopvmXZEOJd+/9iU65P
B36o37P804Kfb/22/N3mdR1ldsx+slwOjWvjN8Fr8svYy3CK+m0nqODj/xJhJ/pdmMTpMf/C8y2H
wyrgy94QmkEe+QHtEmIFA7aqWnN4UFsiQvhZSy5WWN68fUw5tgRV/WifiU2QWidw5c0COwEU5fOz
rLhyxLfl5fw//KMoJUNmd3sDUNccUtTMH9Bs2uRhcScSpM5ge1jVIptFX5sE3ZCei14AKtEK0GWk
CLrU0Ka6MhVhUuW7rI3xbJAtrHm8rFKzldoykctL/SQ0CxDKJ7CtECtpVuF9OVvc3pKyWvQ6l8eO
LB8Cz/AgkjT2l8gFSDHci8gvlQlK0ogljdMFxKcLtG1+i3ieizs0mbOQYsdwp06pJU++NrjOo0WK
J3czypVmo9xaKd2UdvbKM+PHwh9qXvJhT9X1suhWMUhXEeI+0/PjmmaOCzkuv/Ew0ED/dM9a7DEk
CWeduXkzmsaLtbfxMTYuSkcsO0tUO28tHnxH/KHBJo2v5BpsgDDbCNYjXFRIdHZ/KlznPKLHOule
5oeWOuqy7vV8oR3z7ceqpJ8e9aHpRb9d3mkq2rSZym3JMqh78xh6hjre0GYCnKKQMecDCjUYtAkT
l6gNyWs0QIccDY0yg6xwL4CTkcovrnhh0vvtSyiYxu/DlQhAmSdKvOpwUwBMm3huvu1+RkhjcM5e
1HSuUYL2h0zYgO6LXJaTkIC8lg8UtDeeigfNSSiLMMLF2TpzsVjaTg3zX/kY2TpjwHNMUd0NWYjQ
nKswqY5XVIj0//oqa4fHGi5a/+bdjEMorHipOrGusNwHEguWpCPP3aMJp3MpFUcFf5isWa9SpDOv
0Qu5vDW/looIRhgvXrt2A38g5QdEWOkwVgD4zMeUo0aIGuReJEbt9Z041NjOFhL379UChAnVYhJY
7CW3H1+jbcxergKbOgRguWa8L2tZHpfcDCcehjWnA//gU+9iZ0ZlAoDI2AqjCY518drB65DCgTeT
ndCnvj7SAUPd43WfNzAM5Sz4RpSSx6GgyRbtwG5LzfeXtynsZV1E1ktwK7XxNxxnL5J84q3tVI7Q
pkDELqboQHY4wE/1lAJ0+ScCi4mMexKV8RI3vCDJcJieRC86hGROvZ8TDEUOenRAIp5IJmC4D4XT
c6FAxILxMNx9oP/R7Om5cRTINeGaar8HM8R5G4YG9QGtT9dWxiiF0oS9b+Rnbk1VeeWlydNlA2l0
ue7nI9lqw3/TxzI4L6w+t6CGKdDryKfi7geJaTowNbQJqc3xWqJ8bAEqlnMxBEz9K251wn5wOY35
YV2CNINjNYnWrc9pvbq05MKfr5vPpAI1PSleJL6jF2t+buPuT1IdTQQzednvQZXq0dX/uaMpNEeD
qW80W4jKE73rDZ+nmvq5SyW4wiVAOySOyHa+Uiuckx2FeZImmwVdkD7/n8BNJbJDlaNbCogs1/a/
9ObTIo22W8H+oJPZjw1/RawQlms+pXAgghyNeaGnUnKLoz5Vqgtnr+n78KgSnEkGf160cPdscQ3l
GbJXfFP4VzRDcLx1uFoSJh4S1ES9LRyh+gZa2CxIr5W2MhHntduko2vYuFJ/uZ1TyhtPsdzjbJcH
5ZJ2WRLj+FkdZfujwNuCMHDUqcpnbpNNlITNUPxRkyF83J5JST9ARSVizWccxzt/+xv2ArKyBNur
2IGhdOcq7r3I8IgYrnL+KoDVrk4fUfFYDat2j4deW9On6jjInVRUPnlkHegU6E0ZLMb4FM04sWC/
Y64NV4mTBj+57FDEWqCSGqSGc1Se5TzvSDsFBbXc+QHWWFoJfwJ+KIUbu4JDiisb12nFYksbYlN/
CWQr7TS12n8CJEUeIWcRZRGOPuXStY2GKHeS12v7K9kY8WRd8yv0SYRtVzafpUvRjZMxEs4tmiF+
YdTICutPr64SXUdpVP1MkUcFgP9NqW//5hax70CV84cexkvAN+Yt6HovBDKDieM2diDKqyiagLUl
gSu8xpDZzYt71Fsphwi10j47v8nXndz/YSViKLru+W5NJ9Nt4h7fL5lQEBifQFWk2ueBKmuqbXt9
J49znzuvBtVVF6+iT1I8fXhNaTdUtd82eEVgINwnHqUpKK9DV+kkboI9CX135F3xYgZaCgVzNtkV
x7lm0S6A/tDMZxgNgrq8nIkm7WR5UYNUIjtLJ6zziGD0ehm3UPPRRIDjcLrpy3yeoYOXBMpiFooO
9Kh3SUyfPBAO2PjMbl4bf8RYdeCyh3YXC1Oq1980p3r/NfAGitEZYS9l9L2I0RcQAVhFmjF6cQ+K
e1Smc85oARHVj87zPFUDioqufrfsvfSsVsbDf1GTtYywX1HHKtE96zjhyJYxxMwNxSioacWHOJKi
RIBpjtJ4kYOW0JIe06mokW5HKRzpAHvHs827wougYlwBt43GYdHhB5aYcFhlGxP3ZwXfABU98JwP
G3YwHPTZvbNTM3G+z//6oR/9qMEJBNE8y9Yv7SWlYAMTFHwGaZRkenzL3wZCjLWRsrlxszmhW8f6
I1WK/4iWM5THwWZXIxZ7xyaJAxZl569CPr8PrskV4LlSzwRQedwW1yXqWFMVIXLdCdLoJuef30kJ
XBvmK894EVEDOVYs9nCoLi4fEHT3B6NROrlleCIlXjvWuFZJPT8n4Jz/s+2x0NGAVJwy0Wq39js4
H/JvJsGGl/78yfjGhqGLSR4DMZXfk6zk0+/411SnXdn6EaViQH/3ng0LWnqjDju+uJbfKNFljz6b
vDPgevi4EqizkZdPsanaS14Btn7IHIYjw50AOUY+5vlSH4mx96quGRXLKdMBVX5uqZ1UhyMyJHbb
KxAvAzdwRgJfOM+wzgneRjNX5tLiK2ox8yPijCZq/cTOC6S3rK+iM0ODi6l7TnsvsSLetzmP3se4
EQTsxUSqaIZLVeK2kZmrKPdM2ZOo8tYmXONuSTUHfCO88+PIBMOs6ZrSTvDesqlaKZw69RB2hT6H
OJG4gpm9U9G6X/GZ0stoisfOXmAjtwM3H7W/TtrM+6t5Jb0kHQeVQ+2uoqR4QWDs1wK2g4aYUoO5
jdhR8O5QhVsLBumqTuAkZD/xu22ak+mDDKDLVGqabd2BeTQzs+7Hgqd15OVQW3Txni5bcWAwGjbP
W8+7cz50uq9oGhvlWRgGw7SqxPoIIgD6FH02lmKTWqm2VeuRS8jpNx8QOfvZEotRygLiMXCUqEsg
Arn3iQDpvmXihn6tWbDfPmBKXrhYDgWONGP2w4EJ4PmsEoDUTYBvni4fblArH/GkDOpNur/6fC6A
g01QV03XhEiaj6nohU/Y3ijZw8q8vFrLp+4NIxbzM78pGQU/+Atz4Zs6zDVDqUim6AcyFqQBu20w
6wNycminlz3XromsTGZSUryyUlshrvpfzkieUIelr0PNXEkIwtFRsC6I9Lk8DtzHLvgSK/bQXNPs
RkNq45OHUy+0wX00pGQzvLB7gzPE6/AzYCItSylha7YoeLwts4Y9Odmjc6MYgKPpJpOB8fu+BwqC
knvLzAa1Wl7q6wwv06QYcamMfx74Azo7JfFyFZ+/ZbXONuxz1RH/SxCZzim/gXk88Juc6CFDRqWI
Fd06FZs64RZXBchUCsDLrWcCviYYbG9HbKBCvUdS3CgF2Hw8wwyKqMSGdzkRJ1XjzzTnirK6akMM
cv7mYRkTFlpahKuorWJsM5f138FAJWTjAENYvF9DYfD4izC74zUTZHfdnYt3bT/iQrekxJRFoF+W
6q5V8hph0vXY2ZE1FyAHAAin3re0MgS8mnse76I4p4qVOvmf7PycPUTcp9OOV+GN7aTEdpUvI8v9
wE5nKEEA9hIRAIXgV3QacCaSZxQSs+nJQ84+j5QdRSjeKoOs2wH2YzEsigkvbrabzPhGa51Eu4gv
hyakdKmsyWT8D+8S1b+TgEjIVoWl5xC7TtGzHFwm+gDDQhCNdDGeI7VW96ZuNPmacFRoFj0zhFee
N9wZlorHDzrXspsCTXkPG0h8MoAhg5W8pzLm0J5J2l12/KAFiTGzIVsh+qdUF9ZfRmMggNN2Tt1n
0F3E980nSEzc8+9ICdctqbC8S7AiaeXexP7syI7z9j9uPiN/Fm5z5dJrUr9b6KtCoQtsFKemOXwT
/Bhy6kLbcmJoLdZVGt+4HJ2aIxa0GYJZUwNevmFEMt5/3dtPYSAQAWSePJ8GODDdjvRWfd88FQ8b
XA1jZRRoWqDck96M61N5t+X9AaKrK0WtIQ1hfqqTH+nX1pSXe8JGE5z0cAIOaD/WTcan5QCffvN7
9wiaIK1eq8SeUJLNquss8LpgNkYahWJXS0IVtZIKnqzX8FJT5vB+vqt+r/LyIH6GpxKBIcj2bcps
ImouR6LbankGlV7HRgRW1l9UBvSx6ZP/wX935O3HgptYooyNQ7g3IadI8RuYyRHfA4YQGhKW+/2m
Qnr3hDt3RuJ9WEfY9XIE7qpbCkHDmZ+LNc4V8SgFVnu2+QjDwRwGry406ebd+8i0b82arxO2tV3K
+1kFXImtsyNIL/sNRWUJs4xi91t7utYqIee48fdPUxrjhdYQcgnkPPSpbeuwme+KQfOphisvY6/Y
m6lZt4qqJk74s2a2E5HrBsVOeNKk3BI7FTujk6f9ozNI5EH5j8+PWrbBVVpO2zi9iB0Ikofri5Bj
WpKwxfr92SF8TSY14epYF7YqOLLnVZMqD2nejt0sNEI/Twzp0gNi2/oJDhY1DaCdzYBBqouD1Jym
s+IMt/tANPpfcU3WWTD2Sygho8IX8zJNj/gPHITe9NP3yQmFdbrPZZpHgVIbCBQaogmMgfR9tYGG
dM3w51tzLLeNdytJO53MRcJc63rKZEiZqx0gN02jjbAJE+Bz6STBKf12QEawZxIr8cCAAJ1stKt3
nOUEGEhB3T2TEDw+enaZTTxHqWjBC++KV+bVtwiwZZdoJ9tAsaDszakjHfKm9rCqhZa9shj04XWh
1hWyc1i8DKNufrCwfcewax5FdSr1qpcAe/Pl68GeHw6hHHwn6Or0TsdwURp0+dPk8Tne+VXyYXaH
+HZ82IJ9OxWgSeVXu9QW9FQkCzsaJxxeLy7uPN0KCjbXcQfmQMmANqNcsvp+m1rn2y4w6QDGf+Zq
pdxlFeYkFHqkCiVRknvY642GcPMQGs1tOXDMTDsLEL2b9bWloleAFYh8MVxa9q1VFOoPEewv96Xg
Bu6yvDI0hXE5pPI7bdNOVnKf+FpOpO5/4DblojqzcbmQTIiHu53JnCLdQsFvh6/zudaJ4eekxt7B
PYEIee5HMyZozApX95YjUvhwg94vMCFO3tY4oKHwZU/7x3SrEOJfE+ULg/mvCouU38SjQiiTqsnv
Tnup9ohdw7AGcAW72M6uSXo70tqY0ZWigk2+7AI/ubYzLsxfnJ19C1/KNby3R+bwTskQKbzedVKn
UsvncZa0qhu/RE7B6FhsqncQ1n01/LGXVopkn++Tqlf5UJVxUY1pFR/gUsSe8/ug62X+27pvNsye
IRgTO1YmlbGU6ab/f9+/QtZWz0bWYxgteq1Ulvh4YBq7DqyBpaRQBnmygaT45ZQ6X1QFZ0nm28cj
4c9olUVliAxoRCWEUmnegg06Wrk5sqqvmhfum154KeGnL1G/L9hj+Ut+9uDYizFKzXOiYUARoMLs
HP9qL73Ax/puDya8Tvn+Tr3FsbY0mItF324tHFH3Ba+q1r6sStLEFtpzn0cYV6lOwBjZSkNUPvYZ
eHtid8Uk+HhWdmx/Ic7CPjWJ2OPvIe4qAXmAF8Uck2RZEO5/NVGD+XzvLAlMBofsdGLSqBT9tJuq
zziSW6af3c0MFOG9LwiIkHd0ymaOB90OFK81jgzn9KS+YOzB4URzoNOfRUygFOnhtxZfjj+zJDPd
2tQAYbBH5PvQtEGBLadRFIRJxs7Z1A5WCKPMz95pVvR4gqh3yqMfzMhR9HcHJykJtfDZW20z6jr6
AUudjTaa/TyaBq1KTaA567Ets4/1AS8bdYeFkpHinBOQf02tL/iVcZE0RrvlFZHa+aJmndRsn9DX
Gq2JoRo964LYil1axPIddTRIyiG/MnlQY0XZjZUo7GZdqdADMhUIWAb1Snh7xWIwRRQJqFL3j3Px
uoJUaj02hReS3w4iwhVq1x1FSGuJMD4dBid7trpkR94kzXgOymWUXN5LaoMzpUe+XcExxPAtUeB7
O/PVa/eBx5mIwAyk5OSbvyBh/eZ6rIAg+DMU46YA+bQ6G5R2YuS2a6I64fP+tiG/OtP8SU898vXc
2XPjEqh450rwT7Ol6d/6c8s+PL0MR+f2sWnJ76tET6BuWgITdsZ/XM/RiMxBqgZMUsJnqCt0h8ih
aieHGVLbeOruE3HZBteT8sRIywe83rhcfMKQ5q+TWGWclFCuYDeI+HkhS/bGnXcFCOTARdsnV586
l3wgdJPLIhTZ4L55fNK47LIM/KB8rRqnl7aweBOz/9eGuXy9Wtt3HYqLwXamrYelz+i0CzIri3WD
ETA5FOjqfDGpjpnDB6Xmnfc0xtJP0ifB77JKVcF5kHochb65beDIy+RmNBPJV4VQQ0u3lFJNuxQG
UVTMH06bJIXIxbcWXHDaZ1PMQDWD7pG9o1z2/3Err+lbbuGQ4hoOVJKvFlU+R79mL4nFnO/zcVTH
cmkdZprvjAfF3SIE1qR7kfllfrelm1vK05Dz+oyDKG9mNQelZhlsj3Hi8iMIMn2HwYnBkR0drKy/
y+cBDXp4XHc2QBrwwATvFKukCeMcDgQHJlpj9WhqopOVp8lDHbiLQ5QLuzCHEG8H6ffEzlDlwuv/
DpCipH6EfVMZx0tQck9hp8eShgzq23vTY8iW7/dI2eXvyI5aISI9lKz2+en6lipE7UvRXi5+d44l
U77vFJaNZ6GSJfY5Y1JET8UnBk5xM94vhtkh7PB6+81JYZ8w/+NDBPnOOidy6+PSNcHgQfMzO04Z
yCogHrN3kcPfzcnxIu6Kh44z2gLgPsi/GmlVnx14d3e0aqql06mx0xLJZew3iMw2A3o9pWBLClq9
NIleF14S3EDgMv71v1nPVnlY1LIexd+ZNRfA/zBGiq96k2ax9/JbzayB5UTpRsfoRRM1F876mzli
I1g11bn09X8xhxrR5ta8urUhjvgyHz95fEjMtamQszD1ntPZSMMvt5L20F6PkFUKhF/+rpO0GXIt
vvTls4qqZghLdc9hJtDpdN9XatfPDXycX8NmnCDUE/VcelmHAmx3tGqqTTRvssN6GMycQCb19D+a
GKCeNrCSiglL0/SWP2tN5fW7CAqSOvX/2ebEgbfRfwZBqmJkV6ygYFPrUOLwgOzhJJqzq4cZoc+A
V6avlbXtErcXVzr8VWHSXiEuWRdXTgnNr7pUpK08YIE/mNKv3Xtwr0T6xy5HJFdifSiqsOKSN8t1
44kE5jye/BtALicdCcTVk5zwhnZcD0ZgzX4Jxd0xqfdHjxQLezaQCt5gCs9gNNQG2DUz6VNPSXAt
8fnAxnCdGKs8R6ncrhLNwcbvYG80ohDwIxbkL7MHgdtJKDBfHUon/gL3gI3nHTGR0G5PKvQNP9ZJ
SUZdiqWkpHZ1lx7akk9m6kfut9pycDmsC1gVzowojk8NqOnz5tLq9Pb5H/i0zE0arxbc6eTCWUr+
ipSakWzIfDkY/l/2KbZfued5q9YJkdjekz9ZK4uQFy8G0ve0sS1hlh1kbBZl6taZszN3oNePpKi+
2R70OXeLv70asZnYOObp2w0MFs6ytqyLySNgudbVDCiME/qMyl7eqGoloySG3mEoQe/RMNYSvCmn
f2ZGHSxJKopwmydgDLB1CVSACzeKhaxumOeF9sb5Ot/5fZAWPr20tF6FOH6Sx8JOcxh16735YfAY
AGpSpAZAHTAd/3roo/8WXjI+0Q1NPx7qiCnwjHRXaHQROKI1IJIAfpIaCHbL6sm4/F0y1KLFZfHg
t5p24c3e5t01RcqZjQ5WLN1bE3cqEKoAatpSX7DuBy2TSF5WR4iXU2KoK1TAiFllDrxFG5a7tUxY
E75a7zQFFuuW5cwwE4GBEmXyVoq+o/3vU+2i1+MGj2BB7OH8P3cQUSOnehlj3D+GCx27m1Q5zaIM
l9T4lSOoime/WEzPTpY3y94hnZ1ytGbDXh21I9ZoJM8+40HNFVJM5P8v1N9IC3H8n9R3BJBLYO5k
aarpef1eM3jxiWDtOmcVHSCWK6hmwyq7eNp5gdx43PV5TWlD4amvw8CJuaj+F75RAietWsmf780M
Dcuu3HyocPpal0mmj6UaeoHjgfA+HTOH4Z0kdAm+fbQhc/KyBfI3QS1xEkOMDNWW9obpl66odU04
u+VNM3+YR1QXQZ6w0N3SjqPqDCaKw/gJ5avqa8ynGHlwEoFvZM0Py5OqEe/3wCdRAH0oMgXbtM5f
GqpwI1y1lEYUFI2xftgaI4FPee3Td5oSkkj/VEgxdq1wBTy0fr5a/RDzTpcS2i8OZVtmsnZkHUao
Z5C4nW0jGknpfQNT2KQWyrgr7C56r335Na/SyfA81nXxncA0K+MvzhjilJw1gYEnvOwkl1yBAb3W
alO9CmG52Qg5A5Xlak4PO1raPKDAuS2895oJg6SmuqYpMiZcAV1dz5IaYf+6bTrZl/PhUvVlYV6i
wgBuSJIxInFNq+0IHmHquBab0nT/u4Ly0FkQ1j58IWQR48Pw1xS9H5WKITMJdXlKnOJljno2Q0/G
pNBXw3XvxRo41zl9hkgJ3Gl79ZMiX3oDzCraMMUSThMyk6Mf0zuTk3hm+eQ9Cbtx6I0FjmxE7akf
X6ru34vrhOo7P9FC0KpfN7N63PIwQmhX5VTSiHdefw0ma8ViDpMebRsbBkRV0zBwVu+3mX2MFmnb
gikc6wRDHlzbxqBJn9n68UIUpzloxErUi6r9By8MkePcFOStTtBqG5Qc1gjAnTupPjg0SgXwWnWs
QkD/LCbri/Qg6FIeSmqBfp6FO/c7kxBQ+kOmypuJpPqWOICTgAKB5YM6H65YPLlZPc6wppEJtmFE
hQsx510ruIFhwNLMcYgtb5pA4Ll1V+LK9sZhAKcJCOcdJpoMykohswpFt09EvptSIT+3aR4glS9t
zkpmdcXS3AkU7ny7g/bmU1+tA8nVITaEn2iEQdV2CfanHrPqZYGuxKO4oqJssuxk1RU9zGxK5yF0
9f5HP3qhSa1+y95m0e5D2pzthYM5QivEkK7D2IT/ZOBeFo7u2YBKdOy6dOdSfU3dxzqAOAfZAITL
wvQ2CezrOk+hI4sKudCkYWvm9HIzO/0jKGFRvMJm0BrGW7+em0cvCqQf/UsQM1S4Hyy3rVKKZyFI
KXezk5vIkBLJamYIaKZcZupF2l2Hjaq4hXvyiU8FI8mcXjkaY9VWsLn0P+9zITHZPRd+smWHqmQq
7gTD8c2OuVzAiY4Sb3JD6b9MuQuLCY4CS2sZ7QPrwS1w1j52/qYqACgs5cOLVwkMQUY6QO8ZcJLb
QWeTowhxQrSHaQjNCl64m4GLFkGH+x7nLduJx2d1/47UzxuvqLYeckeVOjrQ9BkISfpDy6PpB/ix
oTXgVK0caCP/cVzyTftR0F/1zSwWLfh5xsalb5AgHhiSUhrSURWZgTed+bfHANnQ7urkBvk9gCUC
ONA1v+SBuChVUcO5kfRP9rEWqrdDLfyBQYiZOnP/VFRC2UhY0+j1cQoyoI/eXIxbXv2tjEjUK9qL
j+RH4aOgrCRysGiFufnErf+NwWSZDPrnV3VFf5/lGCg6SluqAAXufx9KL5HEwJbCr2T9/UBQmfOM
r/oOnoLtyZvYrCWrEIwXRLOdvLJb12IThkFXvU2OHo8lP9G3JpJ4R0BwHwn3sk3sV1GhE61+K4su
e+BU478/wiB7iujmoKxHZosOIqGSbnXoGutka7nGvK+oKYmdgpHrbgyHOj7kClfCwgl45hRQvJy4
zatq6Be+lDBnFBKRK333TI0x2hWtHBKUZTg2pDGma3rDXukoSjmMn0tSIxZ/ddjHNX9siLDUuD6I
Oo39KCkPisq2y7TOc37N5cyqWxMds2eFddj/3K4s+Ded6ZZcqsq12fywp306Q7k1AxqmBp3nY13H
bFygTI6Sw8oRxd4HLGcTNKNzPldq4O/GZ7Iy5U2B+athtgfPBJzltcVSNlSeC+SohZF9dMXfK5WU
eyMCMPgPC/t0eURbe/t5/eLI00e4/UdSHOPQ3FLusTYCuV9wC7NudWjGjwuSVJCTguKb6pV9Ufh8
o/qwU7n63Pgap1x1YhmBipIxz0r7YPugBsPcZr5V/og3rYSUR9cuPh5DPkLsIVY8PTvxJpE1gsmN
EG1IA+PbIH+CvTV+6VS+QkZLxYsKu7Fs9fruYszUXVSOOWZeBYp7Uw2BIi643dSdnTYBFE3OjYhI
yBi8WqmP9qr8IKo1unzT67ll3TKctn2MZqCwXrJzC7ezqj0akuy6Pz2mhhFeBurcwSSeQnqCiH5A
NzTIXgjv41Jh8i2XIAvUT8PcB0wjJrphwZe9w1Tv1xCYmoPH3ir2NeVRxtRW5xl/ev2sub1ALyyw
OgZcISAJcnUkUQFYOMlARYG9bR7IV/45OLBn/NYkpxAbGOjIdIqj09mu6TOh1v9zBJie6axwQZA5
axk3P6xHSJvKYaY/vc914UgILaaN5td66n3IeHsty6I8Kw5TsPnHrsOwPL3goM02PpRKD4pGZ5lY
ulk9uAdJY5haMqY0ixP6o9g/NubsjjvwEsrg+rtRDqFVzE6CDwtr5jsmGKlFx0u7DScWOPExJo3Y
XgHzWls0BbJxjhL1vCHoJ9NAkrnXSNeHelbBjobBth4hyZMQFw2aOVTgrQ9oS0dOioawmRTT7mz9
EIZ3whkjPkLXPRdPB5cuqvumV2DyI9YL5e1fS9/Y3EcohNm7hwGoJK8r7lPQn8nHWybMACvyW911
PcaBI9l7u5jYAn8KkcsntW8EvHyoHgZ8a/rd0/61m5m+TpzWpQlk2RjXbCcHKfCobqwu7lMOyBs4
uR1+tsLPYYUH9SPvLHenm/RuHZbwSsfbS1bUSC5WXnHBXISfccAjOH9AzR5bgh/EB997kggiD6V+
G6uZpsWYM3ebqKHmtqeLDvmimZfxEiqk2xIGKcEG7qFUQDcXBCjGKppsIaCK4DEpjJNb5rMXEDnf
3Bb36uMOmtt4gq4/j6ZHBRx5gkmQ/xQapelVu01ZJk0yCagj2Yw5JNiSqwakOZFW8EstqwHZ6C21
DpSHSh2njQGAMe5WcOsYxBLP7ZkGZEtysx/K8Tocen8IRMheZIw6Vg065VVvKhyD//zTOCwd7MSl
L6jrzdQisBAUkvIcWn1YY3zuBZ6E6Q2CS8aOeZImtxRuKCWjU68h2O9H+nUiGRlC3wdagUqzXmoS
PLZwFElyVo1zH44D6vMBN/kD9X1Gd7BbEf1GuqD9cr99/8P6ept2q/pqZhYMGz3miT7dIlA0iiD6
5yz7JD7lPOvWg81M5I+BUANK2fWP/H0zQM1cQaojemAwv1ZJEQ+wJ4FGSyv0LL/Ox+OkifzCyf3j
zFYkfgXld/yiZanBdTmjoqyTWUDiFP/Jpzr/tgaxfOvXapyS4YcfjllUipu9qZ2TB8Zr8gmYSrSb
NOVQAK4oeI4DxYGPWztrGDuKgSY6jXSh1ga8Fai5RuoZYjM1kTwxdlo30zr++N0+Lv3XI6KONrnM
sAK6wKsLEYUqmDLfmrFSflmXsZCfZ/XKhffxi8uMmbz/OJxeR5+cVQed/yarUUrKzHgeg/limzVa
3+FBMgykOKPp8gI0WqaRRNpySwDdXNDN0/rvOoln9Oo7hRDC/mukSHneJOoPl+iuzEflpnKGlV1S
7CSNtMHwefa7GgllRs0eCaSrcSwG/RjPf2Qz/8cxvBF9v5yvcziuaaPbXuQnH79zhW2bLrnTTVzN
SecLFcA5goEMwNBxPlhuNvvhCZR09QAFAE8dRcaPzi0mBUqLNLM9tRnga5YZd1zc05/RSX31NgkG
ZEuprdwd/gblnUxiyTTD21eogidonaCxunJ7ze2ce/NXxfhjnEFZcj70q6OL8dgLDPvW5nAdLFUd
YhgZpTLqdTeqGLYuxp6CNP3fTmycL7avE8XMR6pszZWqIf9PnZEpBPRDYifzoSmUINi8RKi3NCWx
ltYFRjYmSVYXY03h9c84CVlZLKcTN08b73xkyvu/yID0Fft6FBi84GkvlvvgjnMVs0x9oTK62nb2
GtGovGDe/FldI6stvQL4ZtOkYc1Ehuj0PQ1bU8qZoKThreYuOARqX/5zEYtQcJySky3ylsqs1k/1
seMoGlpFLLG8GB6njDwvKqTY+oB7lcFPAN6FbvDnkQs0oUllJmEno1tmk78GEk8bO/BW9W+9phsU
0faadB4Ujoxr8UEIspp0i8jifimDimnXTQHa4RL3K3HWMyicBAEB9z9P7/hfnTPdHi2+l+7vsGuE
17J+xGrx9mSg540EdgaSUBGgBtV3HE5JobLlE4vChSH5MNzylA5rRhUcKZgioete/XDJoD/eVxcj
LmzfKcmuB7Lep8X4vdaeybjxsghno6PFD6in0+3AAnm2+V8zwHONV8aDbUdOprVo99IXELDwzDR8
c9S2GwSnDbgpHDopQIfN17LRkKiZ73ztPa8pQTvVulJc9i7hS/q8QINdoPye5IOHLPB+5MvU1WN9
0+H+lsdKsjVv543znmK012ukbuTFWPJq2VKWpVSTGmJOkRKnxLRaI8wulj+1lnyPTXP1ZbVpA5FF
ciYXiFOyR1fj9J+BdP1DLxcmDOp4e8vYu+ptv3VlbahYNdEei7BomcUumveVOEk+ikd9Eoz7s4P5
SQrwg9/fcxxiu4Gx664XcN8MurnaHHVqxsTZ/Js4u/BUaUMAMMNXpOiL+RIOWwNG+HFSgG3fWSI1
WgO9ZA4RwvNJ3cXP1UDadYf1uGvUmYPfDRcPmFN0V7ZjaDoLXiJ8bL0wn6H6zYhczInu2efSL6k+
g49IN7ls0Ze8NI9O2tJIFD8OJkY5Qqwr3vRbsMFs8YYztBxfbUtm7eTpWG/sMytOPEu90JRoW1vZ
8l7aGAfkXCt6sSWE9FQ2/RdZ2GXGnRwwueQHhD8grgtVHGNUhzccwy77eQGFVYn8N9+6L4BAE66x
VFatY3uh+K8L0/0ezraKkzExzI5nmlgntbcysG78iTbI62EijwQOedr2w2jyziVfPIWfp9yY6mk5
T8cAFSvwG3jOsyOgc1HBoYvPKo29FVYbSHS+bVo3RPMkgWVNG4KoDsnP1z0q+vl3Aj0w0s73FZFd
rxIvmDMR9dxkN8aeOgXS9Z4a3XMHIFqWIS8PZ2c6cG0dir9Ag4LiQyjURuc2zHIZjN4sJqBiHftU
njkuBXi6JihPYhtk1bFLda2olmChs/JAp7FUzaPA3Aip/kD7pVhZxEO9Ta+b1phQzaXqiAWQpvQ6
WeRlfzEE3JRFPrr+Y1c3J9BHkieUtrOevmrngMBVvC3tstEa+gx36+9ZiM1ppuYkp0YCz10bHV45
U0pWr2/IP97hDBuECNLglA+H+Zt9KWM4dxvmKm+x+dOTqtvG8fQswb84RIVXpVR8dcNcfC9U9yIV
jLd+ZU/cVIPGauzsuvhaHlFHr2wrkdPZNuVbg/cB1zXVQFasl7Ur5ip/Q4+0uXjJYibSbGvXXVuE
JoRkCXQNGbHbSM3i+i2uEj5VWKgjVoTgW0E9UNUF8+LiCdiz+rKHN5I5kDsvE2ONU6uUV24Dd4WW
nNHeE8Ql1B3hCkP+LHGNhP10oFoB4hiFVnHCWQ2iw8Fa0PlMO77Mo3fD5Lye+oid/HkKf0pIEzhV
IocwgONjbfkxbMqmJoxHIf1Jska0wNWIZzhPuIt/z4mPiOrFlzGXeQURtZaYM79PdzeIBGYSkKEF
0f50t3BFK5oOy6ACtvRVezxsTyQksmBEmDwgDpTmjl4duIBeJasL6VsTCs9qky3iJUoZry2elZVC
MDthHX5lwd8fBknA1LKZua4A14mIMo431ch1IUtHel+pEhI4brJsCrVU+PDxkYN6onjYAH0ZQfWg
NVK+aIlzMT4HnhGHU86exD5guGCFp4ZcZvl9qj2JS4DelmoA4pzueMfbAmUv4DmJ9nvzyyAMGPth
2yWk1braZ2kjaLSk5ErR7W8L2j+iAw8PexmQNnzMNru0cWHui1FqUgb6tCrWOgOjoRqSH8SiL3Tg
dn8LBAbz276uhyxjFoCFno8NXY1b87ZCm1WqM1jA2KnGlaS7rM2MZ5/kZMmM4LtZCKezw3thc0P7
10b0WzGjStxcQL01pdTEhY10/sGqjHoY9sZ3hmUH/UML7V9ZZ42+okC5PRL4gppzZjgzLDJCDznR
EWahmAXfb3PSwVlV3MuBJB6u3C86vDe9bAe88Q3ada7QNwIYPtZ37zNvBLSjVSdbQmfcdn/1TGl1
x/EZGMFVSH2816pN9WtGuSuHc5A0CGTjzbml9wczvGjwgwLRKYsazVtBQtiw6cqeKX0HH3n261AG
judKZ3vqdHYWfpxfIkAqUGOrKg1+iywkzmqiaufwOxlw3E45qOW0bGzLi/Lv/FzkOziTbmjhWcZW
yT9WXFVs6oxBldTb9btvVUY3FoTyN79Vw4VTYPnHg41rgrl37RD98Ulb7tv1bLhZulQQ9TiHheTQ
ai1uB2XqGHOzeJh6+Yiuc6NdyK0kHVg9SaZGe8ZaWlctZ4S21T93OS2SfIz02BemmAfYeyPNyasA
tzhYdxc+coHL0BK4E4cRuPyyr7IGg7TT+IDfwvc3rMOrxeZZbF36Eqm+l8Dd5F7Vr6jWGOM5FWnL
9lJarm6LKtuk+w87/D/Sb66WZrGIiwLRqbOPX8Hr2D3BIgNCR0wi/PofCSxuSKk57LGNJORux7dJ
NjkNC8qmFCjewkWQF8JlDHRkUbe53Nmw/3AVHm9CMS8LnaF+6fcsbBEHQi1O0n0c4BrVQXyD6eB+
GoFQ2EldtviHSs/QgpNjeSNW/GKQylbB6f9uaktVNJnsBrXNPevgurLEXMBMHb36Hg0WG/u+tfYA
WKTNCqf00eIZBnqvZXaEBDNtVAbovlB8BZDta4iWdNLznhtbEtl+IXcVqIyuu1LEL98nUOmMJeeP
NewbVvTyBpSB7ynJn86lgih2WXn+bflHzANkI7UQIkqOdurrYdSPraGTwm25+myGN8B2LacLe0+D
Sst/NYYc/VIfEyBCsBJCp7pj7Ur+Q2OZU4uV55mG6TXN0QrGbor9OhWeYYWl0VWTluHYx6ppcBLz
qUo50I5YdmbKFeKqJBY4W563vrT3DhTK+N5zjQ8R0fEvljLFhqcDM2XGResf7FfIVN17y44Y/7Lw
w0L+HR9+7808Udt/Wv1aI+fTybWofCP9hAoQRg7wBb/dmzQoeBAcgJr6Gq/3bcRfdAgCC07G/zTn
7CQtILoNViOmBtz6E+zJzmY/R6cnRbn0semehha1t4ET65vN0L2NuwhO2QzpTQVzInq48asBRFKI
z7XnTo0S/Dz6/3s1mkV1xN+sYFng7KsweWJxF2dGgnCll3WFIjqqyTf9ywaNdUYqk54QEYz7DnX9
ItWgsDDmX/eLekkmeRMJ50Dj/iGM8XQsz7yxwDZa7tve8HSYQKTk8iE9G0qtnP2/mOJhzgNCyT/x
2v+vCJ/bpnpm0abaqsFv4/lX7NUiY3UaY2Rh4sV4cQCDetB0UqsAqY5BaDnpXBKCwU5x7evqvDoK
DCzcQ3EbL1yFBQB2L+Y5lpJRhcpXHMQNPCVYOJconRx2KHmxxNq7IlI7pAYw0kgyxPbCm5CTeHaK
4E+2HJmR2iynzny3tGUI8sE4NBUPy0vBkpLXKas8ivMbgSQJsXNOacmrxKWKnYnfYk7M+SUfcTwn
yuSftz2ch8XlLdO6h+IhWpCws6i87zzOMMfYwvgFTHRLcWTEtQTZWoFzdoMJ3vny+MyZKJlc7VpS
pKV46x4xW1mLLrzmrIAf4T/1jZPph8IVoci+qjO/XHSDT5VAyL3EX3YRqiYODdKL7fH4fzi7NT1L
s2ELcJn9SGM4nbAqAsrxRclQFALQrSZe8A35xRHBfO1sBh07XWYHxaUXl75oFPZMLfjHDjebp9RT
eyhlBu9Z5fG/LqIZyG9iuMGm1oQ0VPa245H/dzWY40NMvFTdScHVhoJSpBqo9UgUj0lkeU8+X+fR
Tvu3wstj2+bsLZH448rcdLEwP3TxGvTM3PFnZmwJP0s+C/yZYKnniHlbbhu2myqZsZxO05B03kAU
z+Aur5+QssQUWYzqMGzIloj5vH8pxcOmGfO/IN1Zf7Ob3Pmog6To8T0RyaQcb3uIvl6Ig0VwgdPJ
f99nFuIACxwWtivd8aPQ9c83np8kyy0YgjtayDI3Q1x05m/iFtBZ1araxzfN28bIaqriHKarWQPl
ZmSHEkyz7qMV45Qxq0DRYCyhA5myGgMLs0kIjVR/bAeiSXpbtQOzuddoeONkvIQOhyU7dGOfmdyx
MAHmrGO1dbWCZ0Ow/67TVnEsAdofR0v6lUFXZN4pfCVM2gXWa6pSX7taAL2rHeiblU1rLsJzUfTa
oGaYVAi1FBAVOukrzJxg4MYIt40zuXy2vE4H+bgA4DVP7ombpKAP2whze9Z8bLiJeDcyIV7uIkr5
sA/5P+yEjhe2WtKIPVtEOmmkWZ7y7AGpxkf9maDrxIdHqeyyM6uP3mIeENlbLL/F0TQ4j+HitKVc
z1jIxenhQXXS1Z0FO7dCxfEwmaPJIFd+WPvIIiPCbygAeHmZU35i3b1bVeDCpv/rtsB81K43UQlQ
ttpecLZ/r8TyXXMYna+MiEJYzBa+HMP0uM+9o2irM8HUuuqY+o/UMGfwpvw9tCfHx7tUiRQVrI48
UiCnF1zeifoENUp/ypF1V0GvNwMHh+K5yEzX8QMnarFfnf9ZQAk4CptPHR2aR9IjhPMIMyJBAFc2
w2NMNSt13W9poYdih+fRLjGYric3VxlT64ydOEBu0Q4L2Ip2CDUhU26ReGMVyHHw6MD2j3G3m4pu
udQ2KSby/Pbd2+HGjDr00iKSULUvASTjcsRwvojMgO+UpLBw1PJdqqwZs655QdGFq3pX0muefjkN
wygoLsPXhC3KzL8siRJjOlqsXXiANfXqNkQt9bvS7090KiieFqZbLmfVzNh3k97kQ/Y2IdLD6Yab
pwxzqvkE71Ig79jd+9+q3k1cARcWUJV7YNGHOBtycsr3vplXfps5rqe4VlL+pwqj1vrdN/O5QyOK
9OU5H6AryqhqOWvV1lJ58jQhS0gNviiwWspYuqdF1WgjdsYeL172BPGOQLlPY3sPnErLhxxHAPKh
yKRuAYKq08CHynDMbREuT1ScbJYMB281Ol+3P6jaaHE2KFrkFri+GhdduZYxt99Mz5TT2UdENh1w
JCwRaErfZniQ037aspMMVOmzAzU2HXiWVKaUD4kvlW8kopR/3dtvGqDsf5eriLDuxDN4si/XujoS
A6QBYpzT3ltm62yaG71AcMbELnCgoiPoptBrDeA2w3ojUOotEmaZFnfxxBbv1g7onXKA5pkvVShD
kMYSK5+Dqjo0hitIlZUxWBExXzW1e8Fw6opiCxYCRJ0E02xWt2+1cGehRmg+rBiFVDlON+u3cown
K16YxrLHL7kPm7A97s/AkE1d0ND68RpHt+NRPZ1TK2vt/higfiduuu41hYuqxNkpKWjMp8kf5GY/
HLST+mGjvCrJN/WSzTh98eruikI2DVN0wO2/Jm5V6Vto4iBcxh+UpUvI5A0QgRB+tcKjubIvozey
VNr/14BL0SxOysk13wfp0UpAyLyEoWvy7bS6hcz86oirzsoiBs+LU22AjrAQQs79hOxClDTukHYK
nVJLPnxa0dK2C2hU9o0ff3m7bh+CtiJdImd/FN9ZEwX8vUR2W8AkuApHJLvUXReV/YfmglSEawk0
lSYX3m+rRWcSXAqpgor3F8Pq2cbETep9pyrabpzb4zpzHqDS8dKDZq5HdYxSosjGlxBgWsPq52DB
4r+xC7XKIgYtTd83VcCf6rwzdXg+4fiiUdsiB3QsujyZIYMHVr6dvEjb4p5b+STB+cjssIHwmPbN
FucIDUNRHDSa+v2zUaiqJEVP29oryr2rPGy37SAWqfQSTjZGfe0Y4WGAL77QBhvsjQg8Yi38JNMS
uun+h+vU6GE/uFG4cPmACnv2xv5KgdJQrVab8m6NW4BleBrNdFcOiBN3YmKmzq+fUEMjWlOWmJFa
s4uURTf6EdX2E+xJrTqInrUcjSctrB2PJbrOIu9cbXOJuuj1B/Mydx+tNAIyMYbWGDJ7KZ5KA4v5
AWzL+9LF2/nyaPlY8+rHwJ4MKezyIyREerPiTufAsmJOr97FCH/dNhuHp7ieuhp7BHnnNNxGMLur
IO5GWVd9cJF7NU4LbjcLIQYIl2iWeVcN1DJl3LWrKHEMYw0+EAJYye70F6Z3/p8O2W6t8fXd4MFq
Qe4w5byCFPhZ/I1WH8Q8jkULOsTPhF5myijmf9EafahNBBzZ5oJ+2QZxfxBeN4itz7tDmaZvr3LD
laFVcrGUQOlJifdVjfK45oBg73WK4qQJtsQL4Z5Wd3DUFv3tidrYmE51kAlAhBNeALnF0Kmr26hp
BevD6sbj+JOJqzgWZ938slS0VGiOwPojTJkG3jQY1Q+pEPVjQukebcT7UXCLd9j9fmrHqbrlgabO
+Im/3NT3Mu5lI6Gy5SFi4epJY8xV5I1+mRSntfsVlcFhEtmvJyGLPAScqOdGQuyd/NwyNIwsRAum
RmDL1To+2F/V3PPmi0IlAC/k2duu8ruiQWABCAcXh1kfy0Ct55xBSzmt62ypqlC+UFZgYG1zBXLr
j2IhZKlxUcBG6DlCiKwWWmDifmifpjmzpOF1yFDA8cUKqgKIXdP5hLfZPz9LYmzYb9J2mz0tEsPD
hxIGgwO1y6Y/k+LGQPBIjNBXcuR6CdoLqrLFHw8u2EvOl3pxlUt0tfLi7m6Ylbfd6/yf+MNr1yFi
yFtOSiW3DZh3+2KfJWfM/7vVNuM7EwtPFCUwb7pV9wlmPMEmCLa90yLooqqgiCuf/RM2/lyAESGF
zfmr2W37Ko5i5XcRM9xCPV/Fy21uGQU5L34P2GSGHVVENmMcA9wsWX2zPZfZ5x0LN3YMhu00lR7S
/C4PV/eUTXT4DYSHWylG40jUCoiFHGWbO5aoSXwe9h0V443BxUP15h0rAY4qCPTLrwKgiseAyili
FRJLVTddfc4rsAjKiqtYQn2CZPOVemeXu8+bA/QvmEP+IzK0nkpwyzV0oyLTOdVOXzS/3A0cUDQk
NI1C1xBWyau+sgE5d/G1WIVSZsP6gtvBB7PqzC49gKcFsH8maLH2TASsiPMR7z569Y5Tyw7jLXbb
nGoy8lR0KN9lzOAwUdGK4175rztZtEYUXPQLxd6SQ8kM06w0Xq8MMYtDhjfyBps23bW9OQ1hsRU3
Jf77K4MmwAiFcXfFtfHpAryLFUJpAx+eqtZQqp8eQ61jK7uvWSuFS8xO1t/EgRNPx4bE35y2rSe5
S0z0HJoW1j9uoC6cQAPwTiQz8k6uD+nEFSPAtJa2QTKGsqmYJe+D/vx0+iaiK/8f7SB0KkKXKq0y
xM0Kx/+0xBWyICXwAxsFojSD3vcezt2RAczwR8n47pH6znj72MAdQZSB7dY+GemEE3wwxvo2gUns
WOse42VNh+HQlsGSaaxWkByBy2jLRNxOa0pCIIs0TAah8wb1iN3YPvkH14BAtpLw/9Tt0N++I3cp
gk8pKuBekqnlOjLcjn7m+uoSxL+5VwVCaSyx3ynfYjjF7Xrbc4SWpCB77ZNyTAMgbs+AuxU8jkgg
hkgrZyEuBVml1Yhy+mgWPkFXkrvsGg5KxKQufxJ+htKrsOlxhV8pVGNcoOzHROCqUp/271SBAh71
dHKQbVG3gBTX7iXCRetOn+SSlFOE23ry60jYENcKqZgegGnIevBDKpjmMuuX/MeCsfCfVEl1xJI1
Imy9SjHXE+KvNEt5YQcKSiTzaZWmM8GVJ9VxjFOK+PlIvLzDMBEk229nJwT76Hc5t5ohMlQpgWHo
F2l2kOidfQrV6m/KPN4OmvWg7utMt2IeUl54HkalDJuT2onY9yS1miqKu/ku8UC6Rt4bo0hYviCa
6JU1XBBujWa/OTqhRJ4jh/VAB341/GwIBAAeg7X366m1vMc99aid5nBi5YfFAqnFjjZz6T48P5uk
aDLloHkjUvWQNZ/iMtFJoF4ErTPE1jjvB1iEvOKgiuKJcrlYOX0cmiGNLrQM0Aqrgq1bMniU09S/
z3KuyV5grJXeEvCXgHTVFtxsSHwDN6xpMfxQKBvcpaWewS1No9e0qfl7x0/7q+GYq4xajcYEdEXZ
4Vbj4ma5svigIJpgck3C2p90ITHeLh7hj47YMxrhHCr7OuQGQ4TiqGSyRHL7hlRbjncKe4BHb74z
DKIJmgCcGH81TJhRkz0XSRonggXYZJb169/Fd4CD1v2uPgx1qB0+xObXVvnTbJoQJ/rP12BQd+/8
GZl7ZmmaSmw263Hp60g5dadDFYbHQabTatViiBJNwct4qv0C+y8BGeOIhGQdJrLTDeihSZJeJJrc
htomCci+2iqYX83AvcGADtAc50XemSE8OdZPn9Do7US1+DJmmo+uOexCW9QN3+b7HcCUcEhN1LW9
IwZOmPhyjG3kKVjLVx1d3dm/PMmNwX4L6AdvUB9hjCvScTlKDE5enxe7g6CUYvaHqvmvEmGit0rh
tlyjdgcICFpxLMrWE2/5wXfBo4vhNoUhMdPQi+Zgmc7smytujgH9G9drPq5iLrJ9AWLhU0MiL/KQ
4PMhmZ/1Xrarmc1wDHV1AuemOXkBvgEQ8rQDNmrqRQoNsd7eNUTaiaMCLv+2cJ7DFMNI1Rl+hEqQ
3CnEfJ2qnhjBWEKOV19ZHkjRSA9wn9lLfYyxfXk7wBWyG90DpHIpRcmb6yrVZy8Ctoxf8sbxlpb0
53NvuXtaSu+4p5kIlgkniaVRF6D/NrN+S87ZBXwX1IDcHJ79JpB4KAtlNfgyoGBSfGSKpQZ/QzSb
DX7bi2T4YTwq3KeSRtkvcrW/+FtpV/aTNlmoVK7WHdvzAEvthv8lCeL+eBni7lo0jdJKd6/748iP
foQuCjsvOC4jkODr51ynLJl9NYTX9jThUe0DeUAA4Mx9LiDSoCEXYtS4SxZP3adAOnc1XtVs5P4o
vX6cdJOgfujYznPc4yDD+1bmZh8U2+2qS8eZkPax+TLompruQIzhdjg7DEmQ7d/sLQH851i9kKPf
2NF6gPv6pOZS4T5SlRI0zu1cxV8Oa/vtM1bbFQ/QvpXzbEzxo3zWqKY0rFa8IL/l7Fy5KRqeYe2u
divzclLiEWk2Bhxi0/T7f2fjfZS3v2UtVMOf2vXJYiugfug4VKB/5yZlcISmglLnjd7TtFQfS0I/
/kA0euX2znPJRZIkKT2SM4zoG1Jg9s10mT5owgoSKkUMOeZUv3mH+S94vwpovBpgbdpBOBeUrK81
oE9x5sOWXY4KXyXA1DspEwRVdSZOpahFYMZkIcB88BSYMy5mxMzDoETRxNwuvWqiQlOQUU/YDT3k
dkP9m+KvStVfN3FPi39yiPwCz7cR8rHwBOakrSOu7LxcRBfZRyUPMv8h30ObyYQdiMX7TU2Rrk1e
zWcxJjxUkNu9Zy08+t1dpnCGSP4jcoPShmos7JzHCBK/nXShPlQQX4g/gG1uzVcVe8JNBCcVjrgT
+Ag7/dqn1/CrY/6RnK/P6XI9lQPRywPQHtc72unl1oewRBkAMnwiE7ujarFUVoooTRNWL37QiBPP
SecN6/65TCuonx+2Mt8dIlRoim2okJebVsOYKlpcIDCIFP5ny6/TAuypAGAMJrJ8RF0Pavxd6IXL
tSIZ38RBPQMnAfJJjQmgVSTy4N9eS54mj15S6yeDF8OvnkHJLiVmbEvJ3k57tT+QJM8i0R6dwKu2
G+s7BMepgzuYZ5VCXKfX/oCkZ0FDhhn2FhS+SNx7zGeVPX8qgV6U1rxPFkt3Ll9J8hnKlikZCmdu
WSINagq82ATnhnJYaG5/oq8PjXQ0+8QPvOYTG4AGCbF6IaRvTmZTD1Ck3aatCGYFw9rwcfuiSE+V
3rwiHx4e4UtFg84Kp1AhWM7HBNJW++i6jCmKPm6MCyrFxZ8xRkIuiUZo3NVRBljPmBzK6/j4fAB4
8kfIdBG/KkLcXAJ3gaqC2gL85o7qJiwxGJWiVjW7AeK7Foy4QfG7FIvMvqOgH58j1E/MbWspqoBI
bOkkcS8zHsNkVd6bL2NNs8u3WH72IQMdb76YNk8hC5ddQcnXBs5udTnkFP+A/A1fR5fiKWNSrtKO
b3gufpLQ/DV2XPdtt0vn8KmUk8uHFgDyGmHK142GCt1wZL+LmJb5DmBMdlgHbF/W9x0H/D43Uu6Q
6BcOI4U8eSBNh1cF27CY1dpLe6+oLbYRc9/y94hgnhZ5STCgSk1pzYvgfvUN8/4fVp2Qpk0q/52e
9W1Q6yBlNUUx3Yf/Qc5uTAl9lhs5UuIbs/6e/5O0KnxNkgXLBqv0V79fIVK2IFvPSbNpBhlA6vA8
roXp3gQzwbbhc/fvjograOTaGUdqw24svfND75yAWrpIQ5Zwirddz/kdmxasmAywrl32gwMFVI11
2Sw4cy5pReAoTfsNE0mxHtzaY37HIpOpC46Nbb99L6WWliZqxYXVcC1JvhUxKYrIsHordyrVmvtU
LrNiJji0JSoIUNym3UQAKuSMEXyDCIIei7mtQLDEWa+v7++0QrQ/O1/Au7wMkDlsiQ/jEW/zrHdR
mxeElkyG7ubKHYm0+nht1K0VMPBG72y46yWoOJ5THhAule21ev5ZPXARJHReVscGZzK1q96BouCh
HA6YDOe2MZx7EKP7WBOoW5H4R9L5U3dgtUiSeFv/rjeHUzBccUINcfBoffLer8qtc8j8GNicInfq
K62a6X9p0DUe6SSGXl8Ou/f3HdXDaAt9ws+cSeEu3JwB7j1V+VQ2JYebG2YKmpvC3NxkHn5EcotJ
Hts32gq1UgjXyAm0+CJgyYjiTZuy1/ACQMd0LVPBB28Ct9D5zvEhSmX5QqanqDZHXTvUfZqKO7fv
+Dnb1m2GOlxK34k+ZmGm82Kgx0dNtp0Qtgj2uTYkF/UNqMpP+j9z9Izj4Lcs4YLXGbm6kVfeAN9l
s6OBXN/e1SFpX2PA8RiI2M8RAQwlT/b59wI48J/pxn0qE5CNCuIwwK0/V/6ezHDHaElMthyPH4dj
UiLV+U1Uc3YH7T1Nc3HtN9cUYF2jEMm72JWKgJ1leT/y0aQj9lEz3Qo9KQ7vae8GFNIufQuQWZ8B
5Prm9qGXlgtaBVMhsSRIs0Swhfc6fob63UK8vuOM+tviLA9PWP1XWVcgGlIGVhRWwe++IVLpD6Zm
EjeJgW8auxjQE53aE7hjNe3xfEubEv1oeftkBwf7xK3VrnVSeLF/6zcS1qzsLi4AvgvFaxzvJPHC
0g8gV7aSqrgBpzbKm7G3daJSFsEvey1Ng6KquJMQ54P4LzeJXFWhRcnL1vgsq51nSsRc9VUoP6L4
O1O/rb2b6paDQbEtdmBdl/J65GMdbCvWYWU3Ky0UXaIJrnCAdfMz+VKfIfXg+0YpSmvzpKdxXdW/
7Nh8Hsu5/xFWTqTCVBf9KuintJbp6GrHq6RvNJ2ZAbmKNRqaNo6f7vP7ddb1D+VxZLtqtThn4dE0
Bv0vrSO2E1lfUcxfjZoarXw1Jn2UqJSO0FvSgeTamijO0BOpEZ6cT5A2HuhdxJnwRoMUbAW10DMg
c4gwljZkfJCcokqw9BvKzrbKDluRPnmH8ylF4cGiAQ/oPdHDWHcwACpo8f8gGV5WPQQGCTQBGxvY
I4vYwSwrRSbSvaOZJqCKWHFUQ5EGxV8h9jEvrB1WgV0Qa2H7iSELcBQes6dwzjsQ815LANS4T4K/
7LWlWd/ylZjdX5wCNjV+MZOB73+6DdECk/gdJ6LOOnjCbraORoW+K201RV5WEEqlJTMo9u9q1THU
4QApsFBc4cC+2sfcX1lMhIiviS4+xdqntFljwu2kxaccH7wHwyZdNZWNY1LHj/H1fg6EJWuO33HG
aycUNccqJYKvq8yu/fZyT889aaxjqhCoXMOz0OBh5aj5qdYGPYUDZpP0ez+aqVm317UkC+z2UN98
2iHICILmJ09P6LBy/c9ffDzH3XkP/A0iMqMPpN7Yoa+kuEzPD6dhVmf1IPn/2HPgFJGWbl9bD36F
Cb6xQAC0+PpvqGH+1rwU5RgXP9KfUjtgeCU8C1jFbZmofRWBbcRliUuNikgqPCvwQATacACFAJXb
4vSMHAZ7FLZsTpJDUiWjK1nnXPSgv0VR4otieFngqeDzjHhtKps1JdaIWULLDJO4aZfrWzPL3Xo1
kELtjmQeFCYjFk0crn+V4s3YXbugKrgP8tOb+viqhjGC9IkquODVK3MTvPy8yghG0/wxNNn6GYUw
GGgC8MiiVrcsOY8pokYxO4ekqkfP8zHYbE0hN2dxAijwcSuFCKqoCcyUJ3HV6j8ZVjbsNR7gGkE0
HmJBVSBTfLuQS9PpZJR5Aa2cgyLhUR6sGCqpctzVaFxXwNi5pwlDVc+YvH9fFAHV7Eb+8S6wwEYw
N8KSEiVPH4G6+MdsigUGGIM5a2k1Qw1PaaWbKTedDVgC3cWD3lKSRNrkXkGkMWuzd+aWMsT40RWj
LI/57vJzBAyuAPNt2fMxx9dzKoouTeg5gvDHH8av3/cUGf36HzOLv0pMxrYWqBZGnFbFgiXo7KLW
xINjmFSgu+eUvnnL5P7jvVBoK3jozjNqdtga2fNW+GfTHAixhDR8R+XhZ+aJhnqftoHCC3pGg+gR
SJLsN6inFTm6n8fBHBsCTmhIF65q9mOmBXxS7DexFZrlUvkQhbn2bTFYtew59Uia9WiZznWqgnoL
W1HEQhg/hsp0MAPZ8CTFoiYh7IR03IFrChCjYqoumfZsZ+D0upwyUWQLH67PYzolr5HA+jR5U8MO
5y03RImXM3E06dypp4p/djl5zCxTfaiUMBZgTqltEKgDlVEEZlMenf4Lk/Cgm+6yrsxvd6r2zOKg
zqX0+7tNMteUQfB1VxWCsTgzcd0D654I+MG5y71QIS7SosOuhAQWvYWXbDTSS4zq/1XsEYfhjlF7
E3fpwHSQdav3NIEuHzlXAyIOreC89da/kJUb8vuQo8czTlG2cNdQuyhRD1enImustpl9Qpi53mY4
exFOpMIVyl0aZjFvJORRt40newtKIpfxPoDn8DFlFItXlS88wiNqZKDzu9dHtEB7milMtRU2VGxn
fgmTPCiZP0Kla9UgSO+Up1+VL7PpDWhIlJ2cd/TYu0ea8JrcNkbUG9Jk9WaQUJ7tRdEZb2Iu/IQ2
hhHw+7z7XlcE+1Ju+5wssJWofcZ8FWCdhNUZlTOJMH9Upm40VL/RJnAKwMzd/ZiE4p1Rmebgs0//
7gb119SucONDLuDWwFYIFhpji91iFxWcdYuRue+36xEFfyvKjhRJwEc9gHIbuM4WM+Qk35orAeSX
fpN/ht1TfZnoKrMukwaZCgR8KpHrAKx18cfJ2KWJR6sg0508osuSUI/R0t4AAMAGCgA0MG50sdTt
6irtgmaxo6ff9iiNv38QmAb74V4tmqG78T1e2CiIGsNHAFBkKVPq52iNS0YF77BnT10XkNwZxUoz
adu8JPtv86q4vHGD64GOlhH5p6Z2q/8ndz9ZU8CYYzBkK1NN3i1TNwafKTVih0wizB8aEszUNQMc
62ruhDO93Aa3KkqyigtyWjE6UUd0FRMxBqgPXIe9W4ljDnVZDm9N0WvyOCTPiaPPL4pWNR3VGppI
gQM8mUixfpvuZ/zpBtOW+UBFmXKNcJVTyr0AkcvrlsyzAcGiM06S/bKOS052gndnzPhmoewmGQcS
vGrQ0gUInfmlZ+55IVaXeeIvojD31gwdvmcvNrWMX0qxyLc4Pok7k0Uz7Uf4HA+voFEFZCfyPfZr
i8kCGpLJnGeaSEK+/FEb144RUZaMWiPfHU8GSWktG/9/39eSrIDs/zHVR9ELNdgksjKBgroaXV8o
/2mPbU0YeJ+yQpizeNLC8swqaeoNQ4aSDkH9tsJTo/IwQMOSnrHAqwHAFE8/Pfg+RUQL1pKqKt9v
129vW79Z7XSBhoAAH8QyolNew8kna1FxMnPmIDOrnJQmQCewkVwukVX7Mp0nZqvGUkyvv1v/Jzvd
dDwjNF5POTdTa7+cSq/wtioA+KDB5fWXaI83KPvHwqfw0+At3vvcS1mdNSsdI0tlmSA6x/R1AtUN
Jj9e9CE5lBu0dMO3LSf7v0MWojJiNnFNn5cASt2thKI/9pOAYYacwaC5OcOIQV4ZEqQVEvdaQbmO
y1QTuQLdK7laYiXuYSJxyBxRimmilu/OhUNimBhxaTAZ7Aps8P48zqsEPQScHLpgwq9qaFMtLdh+
xNa6pHp918W5jAe+eUB6STfZCqG09lnR2EmkvfSgwXjeLV0hb2MXaKYrO4gU0WLGyme7OMlmRFYZ
GAEoVZEezAoO9YmcwBVgi0SS+SIkT1GQdOHNxQwIxAeJ+tPW/1yg3+aC2t/mqsInaxl7zSQSCQUM
OcbTAc2sN4tGzJH7DmZ04IIDkedCBo7jsXY5qgTG+tVnrQcPx+OXZRzkdcUabZjCxtCWUBi7rRZD
zbHa/V+sij92XeZigrhOzOFqKiPNsMi/TmntzDhW9qR74a45mL7BliGp6ouaoN4AewpaXH6NmEbS
4HBf25PojF3qGXMdvML+wqVQ1O/rm9O29uy+KrWEOGy/Ehd6JgXVIM3Wx3XT7YXyWT3AYUbAqaNa
e1RoQf8ql7ZhMTbTuxzL6n0g6y3B2D/iy2SV/9p0kkPxGMvyCae6rwLyI3AycX4OnAuehXV9A7RQ
o05Ogx/CIONIDgn/BNf2z7lSNr+xL+QYovsSucxQfrWgKn+zopqd/PsrUFs/zN3G6Jz3pQmhH3ow
aRrus9tay9MMJAGQ4EBsMckaWFwZYbkwUZf3PhPwEeihKehQX0fU9vDQi5unWdWMSBqXUYULJDW9
IeBs1IF35mB9WQ9BDLwStoKmBu/vDMMu+Cr+Z8ewz7R96/jLgAup2dJVSvPQjW2Fz60tNaBAh/M5
rzvwdj7dyVxMsOYReGVxq6+m3iCe4dBTH8yRonbMAgE9G6BuDEuSS3Q9gmVdEpHTSqgy7Cmq5+8w
beT3HxAhvgwuMNL0vkdICEjL/kwNVrc2mxv5S+ZTjsq6xbcHZJjeJTPZRdYeMPMmvvKjTFusPwmL
VYVv+Mbr3lRqju4JVQcg+DnKlxeNTnqUAWeoEYHBkC3wVOa8Rm/eCUnvkZ79KpKTyGSb/Jazd9RT
Q5EHCFk56GN1S0CZN6DaGNX2NpuZtti3bc3cG9wTuyKTO4zx5RFF5BC/GIlzzB9KWLeK7vXf46jz
vtkPglRiN0l9Pwcrd7RElsmGUKizVYjK0TMaZ4DKXVLhW/nxotRQVio4BvoBrTjQl7Vj8WCxcXhg
N7Aq9QU5PlrSRRwZD5piPJvI7mPdmwlSKA5oR5zWw88l44SdgkE+kuk8/Z4YjgqDRH4q8LzFxasO
66JkxlKaBx9b5Au/nHCFa8EN7z++kpFOrADuD03o1gHR6Iy2dR6HIs+XupJmo0H5i5unqdbpM0mn
ySsnnksnGZgTgfVJTW8tc63QXlT1YZiN7UEGw4uiQoq9rAc4PqX+E2ufNX5w5d6fn2qe0MwksRwI
IvW5KUt6OI7sVXbI7X3eAa2LnV78tHHmSZCs1ShG4GOYOb8SaQoiQXvIg2BIcCEdhE88znrAW8TG
7sRWrTYz0P5I9wDZrAs8ZF5eA++eI3cbOltC468xVXK1R/GsFlZJcfkfuBTWnO5i45waOYmWDHRL
vrK2Nrv3iOP1PC3AKLIr+Fdz1xTv58/H8nVsqLuL6Dm5ySIYoDtfzE1CKdxAhYqVfjcWBqeZWPNn
sjkNPXAWklTpPLo90YbLKkTENl0CY6LlvlZ4g6W9cNADic7BUrkJbhDjrWx1Q4bsVTy4+5KpLcBj
a4bgL6SqGtkpZ0HMbt9z/tudcdxawdMLTMcPm9DQKj/PSCwK6wOirivttS6/inMsHnzB20wzv/H7
7MVacdcbsQLNXWB9Kakn6Kbh6jTrpq/ckITs8GrwKLaD+4cTlVD/tMmcTuj2Poy+EAkIT2wH+68s
ZJj3YF0t55OzG2yD0D6TWKTRdIo0bhyCLaNAkGiYRSZyJLgab+jWuYpoa6ngoQtwQcX7W8K/bYkj
lsAe+LfIn/Ij+sa4IU626DDpX1A560i6Sreevc3kX3daC4cAbG0WdG2Dd39Hti8V9f02aYq0iG1A
BRlg9ODOcIj3A8JScsHNQWa9TBrPA18joW5AuOgTxIOfd2CLeEB7UVzJSBdTdkiqYunO1MQuETL6
bcBvOumiWNfeTDNIG8evIu1kCjOQn5ZnZYWH23mSJV/OxdPRQdSNnCD5SZc9zdrjrjNu+RqSnj77
QVbMkEhp5QRkcL+FzMVYk8J1V+2KzRiR/HmRTTwdRYG14SZwE0xwzH1kt5BYvTMcMC+Q7pHX9mUS
vkAo11A3CQrTjVs9xMvldQrjtcLiSS1pIXX+1AxgX4n66q+YCuiOxDYP+HUCja5tC5xrWJ+keTB8
8DEuMvcn2snr6t9kQqFTXSDWM6H/VBwevZXo+ekuXCnv7wBdUvOt2PPgcNZs4CpmKQDPmb4Kv4wi
KCRGUxFiNeuzvHsRtsQrj5Krc35g/5pvzq9VPbYL3/tHgO0aLB6GqH1rB8RtLYvhiUNxeZ0rgtax
H/IFjWMssx1PYN8u9q7JujXYJfeX7ttEmunHZdfOMLeXrJRSg9rXEgwGCiYGi0JWedkT4mg0Cb90
MvcD0qrK7zk6UWCH5LkTz/GOt1glIXG9fE8cbsQe2nEOEv16en4r7Kev6TDCJ64z0dpF2kivGJ8Y
M1zj241ubzEJvgJQG5hvTS5mBNMvZikTRTuGTqDZVQyyBhc1V4aqGXr7NnC0OAlzMh7rt9P7GqOQ
+sKvYI8/tuthogaSx7ZpLPc4TRn9U+uvESWzkTubkcIvkqT9HiWutpd1+8aovRJegHeM+nKsqXKv
Oe8b62ahN098iflc8sYGpWWX0DeFAymHzpA6hSBjpditcYKeEYTJjclHIgeOV1Ma1mCt4b3QLkzp
dzD/8BLjSRXpmweMy2VocuhrYlRU184ie7gW7ym7pNefd+MPRYKIigi8s4o5VmBF804QPcpVI138
8tGukc82Q+UCvDN2zxdjhNQW9WuxZbkR/z2wak2KbSvG+XVKevbOPM8EoCRNDmtatq4XtqwPokD9
OBusy6AaaZsEaaMas3BUHsy1hLlfyBE+Ct6BSTPPE6/25sfx1AhuwKLUB3bQosIq1kbtQW+AubLu
jqpeiDiBl9kUusJOc2CwlmR+fcXaVrNW1SHrtiF+f5E5Ok4LAOXhr0AolsO1GqnA5IiFSXzFx86L
D/52p3Hwm0p0vasp8dD+Oez9crPH0AdOe16FablS1jco5t9llP9wf93MnKkiB1gF+qVDxovBH3aq
BRUHV0TpIs+Hf8V3LW069ty7oTwI02rIqqzKd+lrVwHAOOmGZXYq0wv1XjSWe40RywHBW5ziivab
vztaCQCFXZ1A7EueArGBYbANgp/rU/qjZUGL4X2inZYY0LVftE4xFpfxLurqGzN2dm3WtE18dPlL
yHyYKmgJj6YiPGfYK7Tl7KyV2hS4ZMxIqUeIZSkVyxDpErZRZ3aYfZuU0EhIg77FzfJN7IBb55qh
FpeHqfo4AqIFBnExelIYvkYfjC7GITis+lWzLCA7A2eEWWJOBR6aw7mSWCCHLU1WBEbI7qikl4z7
QJJSnH1EfUl3h4p6KkP1ELBh/fJ+D/QuByE+TjZyEgKluKZ1xddPOpZEqK5rDcQbvG9ovi4MU00E
McqIf7/maYek7xudPjxWPKYmUnJ7IyTgRYnGZhZdH0foJAY3t8aBLt51m+taWkoZNgiYVj+avKDy
8tEsggD00+jf8fqc+Mc92It9q460zPgpL3rO/1cN2wPWfJ1Qwy0zL6bG0dvuZfrHu85aOjyhJdp4
VLiTRSO5umULn1U+Ljs0zHHNnqv+BQsO6vMXfT0YiGLeNdjFNYrSZYa7/qtDq8yM4K0Ydn+CJOe8
MVmGdtzd602HkiEESy3g+AABNywI5jJ8YfEYEnGKh6iIZ+P/uRtyg89Wi3Hj0bEkcIMVVHbDLt43
S6IUmWy4aBGMGKbLiYVoXVlZNaf5U8qxuyH/iGkfuInBm5uzaEmYrBBPaF1ickU4eRVQ680KQ7xJ
XUmQLCNMtEFIZ9UwYvDP95Ik8lkU2v8tvG5wVvuhHyQnNwRm9hkentJajFPDR8nK4XZ5XjUVc8oJ
pqRt8MV5LDFQDAqZdZn6EkYxfWw/B/H0o3XhYgCjheAOfaFwAdC023z0SyToMA1Qhn+hrdOf3fV2
HUJSqlYe9ksR96faC11GVIkzGXre3/fOHo0ePoNbBvWynEd1qXot6Sm5obSULhyhbTZp1YadEamz
qwcQ1FNwgxOVZE7nwZWwz5nKLXsbUVGejK8HGGjgn9lDsBw04k1jgxNYxlMWQVjRCzvtRHfNy/tg
oOlU9KrHuurU4Abt475yiWeXShyf+zFi9gzxIMByxW1aNt4hMixV2Ll3aYKrcV3RSCyaUWzv7xDp
zVDUhN38f3ardaCFwACyPS9zqvjEelEtXrrj6+yc3g9u9tJW7345HqVFsVYn086nyDat36cdJSCd
0gt0yIabcJjojncXBvBkDWD8dna3753ViBILiyGAEgDRECjnb7bBvzJaD8ZGMrg56LHYyGjg75Ag
rvu3O5SgplN2Vdqf4CGPeoitxjMW7gVoDj0qz6D2aoL7AThWVdstCrtc+AQ2OoHFsILomYscPosw
6UYkeF0kZd7dAiM/FJwUsdTX4rWr0TlOwUaCLtMH6z2hwhVHoci7BIaqQF//xSgQkaZLH1PTj2Rb
IFM/lcvoe203HAyMSBWBsMYTfaq7HJn82YKp7WHI5Cae3QwcOyGbDPWcvViYXm6onuywtrvgxRf2
omVWtnWCw/Z84ydxWzP94X6Jxhx9y+W1oTdZxuUzGgEEq1hXmSSz+XtaL3vXWcMdaQ7cFPsRUeXW
3Av/v21q6EH8fJotoKT4bFGR8eK5mcF2zLdoOLcm7xLjv5KomKbz3Rte5jsIeLEMMHBaV8IdheEu
vvW3scKoRyCsHNGmjI1lz6EJQZtZ/u4UyXdrUXIByzmUctfFbTeQGumkyBMRR21jGuS/JtOkdqGa
SuwqY1ao3pMpjtfTI1jD/T7Szz0AhboXIvJ4oKsqnUaD0ZUJI1ZxJfH/A+wZrZDJ6VLcKdInDsPm
AtggL+5vLtlhLwzmUBdALfzPTr7azhyYb072AvauC2A8Qsw9pZXmNdMo6fRUP5jNglbKpyz/5PKa
EctwJvj0BUb9G7mX4U6TqglP2Aa2knYdnMK/BIObVP8erTH5pleBVBegE8l1g5l5k7dgcefSEOOv
Qd1sQo14RaZDUd4igy7Np5W54ZsONAZXZbVJhKW3nOFg3nFuLhz4eI5k5bE0wKM0LHI3OAzaXhEE
FHOcTdk9FA5M6++Vf98JvfnkTD7qnVK0NvlUjkp272/C5/FUrVAedPXqLfG4e8KdvAj3B1Re5oub
v0Mo78CUGuupdEXnWY/5d+oam983o8xuQy7oZ4P+C3QF4jT2om1uQVX7IAnqHkX82mfYr2soEK7F
nY94KOd8yEx4clKcq5BtoSeXicsxnubIi1MCdgb14j01/ApQyYt0mCDlPTeEjuhhOu93UpR5Me2+
uZWGvjCrkhzh5ZobFh0fU61gfRAkkW1DZ6kLpYXe3iy1BwECj1DW0MmjKFmtRyRR5FZYWUEz7Llr
1SYnpmk439zcjvZAODVXUK8VqeN4sjfx4+zwLUfVV4tYr6/EbHdK1m547T2pGtrMWkN71DylAkHu
uTlz1MDH36axdT9EJH8yBrVDAfVbpeKI1KHM5CcVva6kD8az6gNbU/ApLe09CXv6WkCwX+LhGZTT
+BrC5NNxgWnrF0I5CVKoakAzWSoV/r1XRPvaxh/SXbcBET4CfhI0aRsR7NLMI2ML43pGw/f4BZNj
vPMp7aPYDFqA8nzV0Skkkg8p8LRhA69aRqXaOuTM0v84GzzpnICuao3ZIrWnRijSdDoibrjDIoCE
Sa0GRhCdiLCqXkgtrvXkoXT/JsHnd4raq5UEsjbA7zSUQ+MUc3nyrCpLcYqPFTI1UIDa4L53TDn4
+DGbukrGjL9tjohRlN/UG+kv7uEMC3BkqjqEMd7kUKWwl5UDo5cFO2DSXPhDmmQgrT3HQzdZcvLf
yV1PEyeNTHSfJ0MXYLHr6AIEVbFKV22gL6CZmAECSuMqFuZ1Sh3hZooBxv3xBFR5k+vCXHDvSbk+
QZ70au4/5YmhbinQ8spDCeNp424imBXi+RZzQ1dhaH/fcLyfhLonaVy74R2Wy4ENTauhW0WBGUdL
jT3RpYYJh4PPVOS+4vkzeu78SIeTyVbUFhJ/nSIhmMhqmbr6vCgkD3CkDX/c+bHhjukYEeeCKh6Y
BLO0bKNeeysn6u1DV+DBBOYNJffOpPdULLYrAuPJGbvpnXY/FAov0zZkuOZ9SEmRI8hY4XgXqjLe
4CEB/iJSswoFNu9bRIGjRhaSQyMOMGnWUrZUJkgUlz+t9zxEe8c8MCqId65UC68U6RoNhkiKnjJO
3tSRJGgvsTLVKHf71L80/L62SA5JvXGQmKGqDaNHI9DDVRHnMTr1gvp9a9lb36ZJDqV0bP1RIaum
jqPv4V15oxwaTUiscth42Ijjy4hVUMUouMFp4+fOaAgc73btGettN/pyxvaDT3BqELsSufsIZOyY
o01fOWFohjfYuoXhj7F+8QwytGIO8yTw+yLZHKrJDOAf9WpyIpWcGyYBcmZUTXgVxjp7kRV5kffA
HzfrPMnjK7Tj0vkZlF7GbMXHWbrGlVMCNm0DBqHKdhCn0f38NpvPKfCQB50Yfj55gBNQpvCkuwgB
yxSGxUt49ccqJhl2QkUKLieGWzAJqtYiphjCW0UAzQ0YwcjpB1o2X9uhnTzgw/KLTjNAJ1joYB0H
qwm4LLdoDIMwIjaSq3ESvtlqOBdtNaFxqHoKXFcaGTD2DI9As3Y3J3dMeKviZ87c0an0QEsYpYEb
ZWgNfZnkI6kbujP94nXQEohFjrQ/D20P+spMDsBmgCsRA2VqFcIX8u92mzCrniddkoHO2hq5pYgK
A/G8bOxQO0nBT+4Vl9rK96Pc4EXPK3PAkewVDM85Qe0ACP6blXvytgbvNK+jKJhcK10JKxDTHXLd
eKo5GIJnkX26UISeUXuZ3Ok9qneuoh6TDlKoMUI1HtYZHjTtMM4OQs2Wc2n9KtXKqUD82DlAaJJi
CTiXNmefWN7Zq+PDTA1JV18Q3b5gPtUi4ipA8pghEBlFKkTVG19M8RDID3m6cM/ycaHoQLaxHjJH
OHU+uw85WyvlyMRREvyabGeo6OlCpWVM4t+kpfgBb3WBd+GWmF+9vVBWSYG1l8uctfJE8+fjuoEY
RK8VrlCnLRdn9DA3qFMJ+zODKIe35NPQOiOoGT+Wr+w/hmCsOB9hYbLGd6s2kqU+IQkAcUfOLGd/
CrTD4BjA2/ruF0JSh+Avqw+a5BN0rVr6DmBwBFK24CHJJGUQg7Mqazh0ZtVvCRhs3Db2Ljybzjj+
Pzy9n8W3Ki69lg2C2Mj+wgqkdxx76FY9SrctOX2ZNbD4qzpda3emHJrb4DHgYZXflT774K6BQ79D
2TVav7w7awGJFJ1a/g9I9wfYz0dzDwW88GcIOCL0nWdCqqjbDV8qwrx6SWw8h216IJg6R7JEVZYt
RaXQ3xzsjoYOw1vPikO/Dun8PR77n4kRNONXDi+BEhEu008weT44Pz5923b45+CILlKREv1PAEU5
9YG1TKpfOKtP0MYIBsAXF2GYR4iANkCADVKZL/KuyWrgjeP9hC3FGXxwn+FmZGOk+n1sJb5pc3Sh
sLw9YyyzER+gJy/VyYnlbShV0RPgIA+gS+Hzy5rFZHs+gjeljvm2G22csPJT307AfA2qFR3ZHYz6
gfyyPJ3o7doVjfkbEfCtzAz4dQlXxIEs3i5vU4qHVFtQsGxK+c1EI+cTRa+Kdd6C1ljfJmIEJweJ
e3MOWknzb/GlmQLKaUZYwihwmF9yx2/F3ppzBK87jvweLtSU8M1Vpmkx/cPPi8Jf0YffBuFwnjU5
K3FI3wX6Ji+dWunLCvqY4FKk1qMj6KALm9bXSLGFZFiArsLzoegGRenQTOcq+sMyDASvhiC49SnV
bECmlTAEd8I2YGffcGWdH4o081M1IZ5eCiWVv+6Vea436u1whPcNRU6gbtF/AQCv1KJgn9dtCSO8
s+UEzi3GHTB035OeouaZ3LpgNrzMreSOgBLnqjS6mOKDCE49xBeTZE1ZooYuprXN5aTzXM7P9zff
9k+Y/RLBAz3vDRjXPJ1ZgAAkV6tW6KaDP4Gn4X95pRP/rOSXwP4yHGWKcwDNrIY0q0b89E8VM22U
GGFCc3VxB6grFfatfRKHoILlyj08B0Ldj3prb0tJDewFjd8S7lk94K9MWnsqEdF7vXIoPNUthJgA
tBbbPpxlHimYT81u1XuK+9+Ugbar81CX853rsYrla1wgFiRbC3KADxTvkisiZc1D7b89HSXjVY/D
ZuCAw935jRYbC1baoool1r52yPJ4jk/gXWaSI+u4TKuPR72hNM9EkKnvoz6P3r5+eYO/VN59q6dx
M7VEbDcY3G6hkW6W1kTjkJtl9od7QWQ3P/F4GtW/+o39KFpBWDUbnlV5/9uJnrFcTgWHlxbE4MGf
ATkYwbGQ+d9HcWB2cisCEczG1TdmmRIlRI0aiagXQ/ZGkS48qnEWOxVpHl6tWw6JGQcmom3XNi9y
O4W4phlhRwa0xbcYiqGHLFBnUoYDCPskzXb3hyimQK2UahsDN6GSJ2l9kr3cx8OsuhpL98loUnCK
TWT1cPzFWdyZpYdaMAlsgd9vsTdgg3r+zq8YuGn6BgrZ3Sq/ztSBVOZT9xW2n/XdoNn+zPILuzbO
4j2OEo9AE4gUD2D15XzMcIahwR5nLRpDrKBJX36qoys5s60IHVfA9eNN/pYB1TAe9weOmWPpl+KJ
3CcOOnbmM7qBzHyroPK0X1tAtq3Wj41l08VjD2twf5QSLRfhcYeV+FqaOR0TAzsiNGzZXjWsaA4o
mhSgFKlbRTZr131TG10TwdVfJ7CN0Z2tElAQwQsPQARHidT53fNuE+BP8L5nWu3omZVthnsbuRpd
Ql6kC/85O19vWt4DlQ7Nt8v8k5gxIw8Id3O9zGr8tsDTZkV9t7Il0TxcQ88t1wL7Pr/SlD3UBj0W
eExdpG7MIv1TtExD3JIyjg7pPLsHl2XxT4Wvm+bn9CY4DM2ujAsaxFeGttUqCYBS/JSyZ9pJfqnA
15cnvWvCFV9eMslaJzwjWq6aQCviWdNaxMhE7HpKThmfcafROl8aqJ1WUoMHTWCRWCYZzpQF9RVZ
pZlxu82p33XJkFF4En56G3YPFgsRm1IcDWquDRUnvnhsYahlo+M7/sBs2ziJXWogb+wyCjBdlIFy
lMr51h3i+yRHC4d05wLiWerQ959tYKN8kIbP73WJwHhK7BTtUAgolfP9Uch8j6w4lqfFRRVwhcrW
em8YA/GX6kUVmGm82rfoY2EUL4WmGLyBWa0nRSUdcqh3113MtwMfa86LCkdtZWHAo6ZDl+LP4aAf
goR5qILQH5hOHl2+6/uEoWt5SHtELBRbj4VCvSDQ/czOV2Is8V9XMdhskarQS+tZh4i3r9nVMGSE
oomlBHErnbMR9i2CNfQdE/r9ThLUgwuxsicXSbK/C57AAEdPcXt7EG81I8ZQJyNI7wg3S1SKoOn2
wecRBLgqirhGibPjA/Re964QKvFl1Muun8NAHtKTh4fOWjwZ7r02rxRSXxXATF5rw31ylEcDjcTN
nNxicl5hPJWGUzAZpmQHsQ9yg6XobpPiWuBtyzdRC+/KO32OsaOBDgjy9OllcMu9QmbT7ctY+DtY
Tp8zTf5xwGzqRIECs+UJiqTMjMYqndT8AaDMW/j2NRhCMCZ3VwBbmlwrOr7c6ZJPVofhdFnJ//EL
x3OP4Hur8NL7b4e6sfegCT/qwm0L818U8ssypAowP7hCcX2R8dyUNVc/DQnmdHQqrY5zIhrLwtli
VESJfyRmj6xER/iB9ZUex1xFcwSqFWBd8+B+WW/q2HpF+6+e0wO1braZ8D4AhpxAxIx5zf00hL3L
jvAolJDJScPe5ZuGEcP4zd0CcthJ5Ld0Ov9smBIWAclKRFCvw1Lv7gOfUf1Xv5tHkWIrexGMJOUQ
tKZv4ExYelE7A1Ml7/QDPZf0j7WroN5KgGF5Ke6fV7EIJiWl870r1uTxpr32yiuZcyAFcqsF2UdO
kW00aiAcaGO5WbcKu2s37uTBMjx2NjJiOsxTYqqCDYA8ex8H4VmXAqlQ11r6taGxdZVShnN5rR81
hJPNIROcSVwDQJWatuKwUKUClLt8++XD62nbx28XHZlX12bH/HlJbhmzBT38JhYz3wTJRjpQQIYg
WfdkHk1BGO3YCJKIggsaJdj/diCGXE3ubCMv4Eb+rF3bkqhceh9AsCQpvOGlJk5fgW4k/UlEILDC
+Yr2Fji0LK1Ea0V6mA6hTrFwmEA7HSfPxZSmlzqqVA2X5C19raKno/tNdnQpDae3fRQmXOBlvJmD
VZjl2hrMQJ2gTfottSvkcmmzsQWTVFmrc0v8oVV+zDtifcyRv+dLtwRD1zGE6q7QuihlPv/D22Xf
iYhpGNTec8pbhp+tckyiqUS/+11qc1cADzSKzHbHYcEZo595QUUeoRTV0SeIJSTWQLETF09TxFzN
Gg34sVmlK9X0AMdY++8GvBlNtiQSZkqH1DccWWGFv2FRQByOiZRqO9xkedmSLzYzn/kRANuoJmxF
Jic1CTd91dwwV/VMP++t5UD37NzqnXfHD2Mta8TzdjUzr0wUeVWp4A/3/PASt85kQLlLzWYtnoa5
ii1FYCNGlddfZA8XShNFAlwH+8fg/rdL1vO+4vpKUjMK4cCoVzae3kNaocoe6/zv+nAeYmXbKi94
oHly3RyBdxwm6/3Wm6GdMf9hbxL6hy757sGrenFXbkfNceWty/JX8suhC3Q5nBaen3L04DV0WO4Z
dF1kY0PfF1LTqHo0WRbE3GoJLmEkddOVtJPhdkoggi2JUC7N3T/qhuVk+2Isn+nh/OpZntPyW/J3
GYLK8hgwsonVPFQ+7fHa3h5GwlyaooIlGGiL4uWK/Bm+CfjRReDlmV9wn3c/cVppb9Jk1h4JtYHo
gXeWOMF3cEHBVWXrGsoSSZOxSVvqfyhk+XxCjJ8NThda6Rw08Hgj6fCSQVtaefrOF6ad0K+m1Z4l
mMv/awxuwUem7RIuzj9oXO0gh0n6CkXtauf9PqqoQBipqgsJyD6odMfpz05paHAi5bV0TLOfASCg
zFNVtQgJpHdFXYUCtgTJCrjj7VvAZzUWhlMH2tflSA6wLczaHSFU8b2nPR+jKkBNjI/lEnO+94Eb
bU38PGesMfVQMAyEWvVyp/F5TBZ5z2W+CdeEbzs3ZtfMIdf544Z7qn4ZCO67OLO8Zg0J7khlYDNa
Q9o4P/kD+trAqYhqQF6AIicTV4Mt4xabRBwZgh/srOMzVcZQF9FcNKxGgxggTD2Y2/+hYNWgTxts
jI1AS4+tF8KvGFlw486WCEmgqF6k1L3c0ow8rWg3CswxkX8AN2fc+wFm7TBBGC+mtCPlGebzZ3Ou
vVlv4dLXkRaOB+cFmQgzcdMqWLQnDbZFHTcEmHhF9DalNOVnXFRfl4Mk2twwwrMR9YKuj2bZUQM7
RqDbdw6ki+4gfMxujKD3W+n52zW2z0WTcgAp+0zzb5aoKER9QMrWTaRrfYlHY7Q8DWm/nBnHI0tV
PD5qBDXP+sWFOHVFhgs8+s2mEepnZxMdE055s+izqUSPBLV5YxSYpbyxSNL38Kb0XLXga4Q6Krgh
QF/DkMo4bvED3MzHf8Lyumwrh8jgDfcegpP+/p+cJMTVRX1wmzPAoklBVFYDbEiy3vuEF2tASdtl
DqNcjjS38YPBLqOgaDA9+T4plLI1OIuR6f/QLvXkNuygrfZ2G/2h8efWlKpx2i76m+0DcyI30iB6
9unIABs+FXJ4M5UeYsPnBK04V8DXYghzyDu1RXCYpfslUUF5LnFivmqLouQJMHTV5pKQrUSantJz
bqaHubRgdD1dZwmc4CN916OfhDbS38CThR2GojoYKQX0/JLhdCdp/lk6dU+rwIfpp8uDBBtDTQ0P
Wwv2HUgqAsFIaKzFutMIw44Q+mjC33k7qXrVZYkaus+N8JuE9BIn52e4eV4dgHFt1Kvu2Rba/leQ
tS6Y3brimnSqLYVXigaXQA9OLSco82F8TeCDok55WvTep4juLRvFlWgIUZ5E6zBH7dYOR1/dGUH5
9FMhY/FjVkWrVwlAhGm320rCFG11TH1YcMOJCrcxpvNK1177dW7/NyBWHOUVo7hW0sXTifbpOWrY
VwVKgOAwyZDz0P11wpXxez923Sk6+Kvz3MCAaYJgPZr/3KA5J/UVTXPNMSznH9HKtQbO3khPm2Ik
6qCpPAfJNxDmvICwUmkh4ofofiB1Of0Ez+v9f1ZqdUtVITGhiGDB0xoo0IWSb3jOu3+uVnelt9ci
K1Ierg5TGZU9US8oc8jTNPaQUQISZe7n7ItAo9l1fVnORKxYcUBm3WvUWPHJISg0SHxvaRdwCI2u
dEDEdQgoVOf2A+8Fw5yyeLvEG+sPeY/lu93HLLCCw3jR2h6/73lcCZP/cOWF2HfcW7YFwv9t+yIu
R7iv3vSBCOOuBXl3nFLt6AB7N3hQ5/sgRjy/3wlyCF6qPJVaZ/1IWdnjc+mPNekNJJ674VnfRiA4
/aSczA96epXs5EZuv3b7HVlIeXVZGYR4epx+YS7ciJ0qOjKisOaNl0qCdzTEZMKTHIsZA4FKkZVP
TqWQmsWjw9ZwR0TT51LPKcGWKuDYbKBduk8bwwbeaiNwlsSvxvJ35v1VppT8JM6ITEAqVTynOFQQ
m9oGLMmla44C/TGTzxdyFnJaTWJ0Q8X1mIjP/jxbm1/bdoOvlaz5X9aEseArl5Q/jjZmBjQeqM7d
/dDMEKbDvxAZTzF/X/noHLaT0HMdxrsMxSjxvMnznQQ42oezcclCk/n6ZTOWcbyrKIlvkr9MYDGC
kvxVAVBC9sTI2rb25pProJZdSl2VM5KE6BP0gBObr83ZxRJdgyrHlLQEBpX9/V7Cilfdsn+jD2G+
UaX4GSI/oX2KZ4+g7+A7LLmUgTJh4HVTtnTAGb+jcIJ3s+lvXbhsEn4+P3fzBdKJTO0XNmSuGbzG
Mhqlq1kCjjwDJvTfwLPRjBbi4BlSlJYD8qVdMrJsnmrmvkg/DtvOYEPetszU0o/O8A7/WSkVJzrs
3uCJan7LMRpkudK1aAzn2c+xbySwBuDufjH4Imu8BRVyxcf6zmi0i/N3+GNGh6IRJgtqC+ELAAOM
iueg1/XvSU+8nyTc7/Hb6mP8NjF4RB7B9CYURqVAz13E8UKNKxbnBBKGIenz5R5ycswz2J8qHsBw
/cywrXUdMP0NPykNSJVz2tBa7XDpcHGX28GMGEK1M9QLeFfrLrKf+TpnPgVnKkzcbiiiwHzZn60t
4h3DSN6qbMS9MbiHWsSdMqtSmNgH2H+jPAL1Hld1ykjY+DeasHFT0PmbfFNwuzgldh4r6rS0UIAl
CGCn2TEIREYH+ddxtCK5vNbt7WVdTWuAyb2ZqVU39HBxcUmY6Fq0PKz3CtV+1PpKD6WXSZNg5obg
qHbV3KOhyi3V4g/115AeCQT4Thac+Hx2wTTK5C5JakC92492/1kq5eBLjh+ZONd2ZzIySN7nqUBs
ofd9ib/qdjsUu8xkd+ZnvhbV4L401mnrTzox9L8LyV2wJqIA7a1pkjl8OyeWp/q5C+LWWaT9ySdK
nloQyxlkoGr9/cbu/a8+Jjzr315rMTJFv2ivl1rD4pW7gANJCyNSns6A8bU51JmIeOYf1hBU1TUJ
Ov3NJZsUDzhwR00eH+nxKouBqgGqkr3bTBRqSZ4XUFQxZMVAfQ8AhoF2O/I1WN4juagXH4aFbmM0
2qAn9qHDPon5x9MyaJmQpsJNlk0aJDNpJjaXUDApvq8IxRp4Dfs6mxDkjj+tW8YPp6ZRRMYaK4aE
DHdgKOQQmLVlkkXA10VI5ZH8cFNhGUm5syUYaLn8+9UXFgF6NDsRUPXInNfPp1+XfJc6HblMcGxI
2YK1KrBpDb5ub7tQ8kZ4knE+rgY+slmnRKBnkHC+6Sgn7XKiYvszyPR10GOUXyUX3yO5zBlOY4Fq
LolTaMsgsWafWqqOd2yH1JwpthP4QN6QFhADOafU7nXKwzz2iu/MVvFZXIkmfnBt4MJEDqIfK+PF
RVWi/hjYRP94PiDQFgC2+TR7C18gJKG4s+15bQxTcrOubjfKMRQAcQ6sM0EYH255jl2GJTHbwrQi
+09N12gvJVua4gKpMhczBlF9sAci2HhB3fJduMDN1vYKcB8v3bcJbISZi3X6x19uwkYSS1yKipyv
P/gzwZ710s8Q5XpBVdhtJAQJxy+f45fjL5cOyEX2ltQA0RBwbTd1dBKVPGRYWFGFusGkyiMujRoc
mbeSexDrR140KaHbbLSgJir4PA3ZGMetpmDXwQF0FiSTqUeRf3SNirzypHX8v7hlCTybd/dY09Ha
xWqpe2W5ksywjZm40iCTzcs7HCRu5JTXTffpDFfgYhPK3RCetWt9tANrxwIm2IVICV3cWVTBMB9w
94egxcyI0K+HNfmTVljevNflQvGxqFoc4zmMz80oW8Jtcy8OI6lOlmT1LLEbryeoPCXix0x1Exmn
kgZo5ygfUCHiWzyX0NLVpcDnQrrb6nI16Ay+VP7Lm33R7tp9dVkXjFSOUU9x6yi1koJyIXhy2Y7M
LzNsVVT8luLuT9VvsXgXN/w7hbDZWQfDF6UozsTb0R8bEkb6/E2AstctO/HhW0o1Qy+mmZcInBzh
SV4COw8QR+3hXxT1ZATQNDOVBED1PfOLpgbwUDPfQmMpL/Zf7OG5VgVqHnsGWh6GQpU4NHuwxyz2
pfpPbOcFweSBI/4utAntQCNB9zA/KpfN/ZA7zKU24FTS5UXEdM734RbiXnidIVE6Hm+9cv7RMOFG
o3bJT8eIcSONZl6Xv1BpoTmfy8YYezUHXVW/8sAUg8+8POYubQU8ANhy+wWVrXBwIT5k2vCupqSr
wy8ijfpfjGrTmBn80UDRZv9oipMDdgiWwz4Ax9LSIvrHuw0k/5oAJ2u3/VbZ5D1pAoPPnc+5hQb9
+sCwS/q+ocgzOlDmgQsb5bX19UK8kP+yqWD2hJDzmX0KJZ6vtfMDWKBFrpTv42OZWH7w0g7H7pQd
b1bViyADW3+y8TEFoDPg3c/6DHdgS3ojpqJOzFs1QBLyyE+WDlDxhsSbTDGtDjIDS8mQFeHF0/3n
ujv0j/qBvrP/WlzWjEHqZsm2qXd/Ck2/DVZpsqS14m9JEBFeBCVj82S3Ak1ZMq6goVtMl4YrhpWY
Lv3/BR2NBEkLhJs/KM0UNF+DVci+phsE/RE1gZ/2VEtAkmCPUgu/yqmHHRsG5r8xACswYYO43QRY
WTvTtUKOs5+BB/B4KqySfETDTNfqL3fvd/8yChAwxxG19GcVQsoc4mENe/v1GNJu3Imx7gqRPboZ
jkeV3JonGh44H7HgdFJ4rddTNifqugioucmedY12PyyfFSEQRRSCK8u1FP7pwAvONtL0/g8wXprh
V8siUu9nHPBjjyZkY+jSUAbfVgk/alXdnOY+BPqIwHsPPYHy7nhWKK2+nPWHmBs8n7bvhKUICDRr
pngxfABLW/6mBoKFtkS7HCod1OGLs9RNH9CMiMJzrVqV/XdLX2yni9YDIH4QwbXtsb2Mgoxl9e+f
dGeGQtQosyiy0Z+8b1Y7Rzo2CkvxW1ZyPTHX9kfqFocUT16SSafiPAvVCEo3RvIJtGgbAqYcyhnd
Ii/HSBt+ICrM2DsELG8BKT3Gd4bQI7DPG3hRAPrxpDE+WwPiHWdOHYOPiFqgOjiPrDY0ohPHjWhK
1cclGI2dYeT8C91juMYJFAnStssIE6XwU6O9RL6IvQfjEY4Duphz5swA/ji04VhnXPXDB9ppuciF
21QOKDrc4lAQxxbTA9oWZ+0wYaiVRNjjIY8VcWgGHd+S/sZhs82lIQeKaZeFHMxhXadybC15YXrl
D7MomVTg0RrcXPbDVPC9dBHpp8mL5Jes+BWQeQf/Q2lnRV1bChuK6jBUwEKBGtptaAVSSO8Ps6W4
2W6fL+RqOu2WQGH0y25ieh7wArvLvhx4FOFt8qOMi4ozvnnlkZxzyWXRUaPcuBHrrhNThxgVAik/
uKDl+Q4QnN3xLzyGPW7FFaZQ0V5gYiDslH0/mA0pm837ejT98BW9TN9D/dbGR4iQoN8ejxjrVojM
KlIwWz+9PjOf/3+lGXTFpecyeARWNqSQOQuQZOLblTSj8LM6gZ4J2Co6KEr6SRGky2pqd6cOwVBo
TettBjRMkfAdoeaXDrVbOKfs0eqXCcPu0/5edZdXYDxAHYs2zTahbkqkODgDecWipc6wiueBYEWy
+HFwoGJCvclVji3oZ/dfM42RvM7bAu9IhNvzTBY3Zvn6/EfUHeGtyuB4/SQoOgL4fxWx4wNYI5fL
hGhVJkd3VBKLwBqEDoiKZEYjaIDw+++oJtSbcr7dmnWod1+6LZPLVD7Jnkr83MG9+SPGwlezPLCq
33KzeLwPL2NfJZ+/CjQaSJlamoBn/GdKS3Zs2G5QV+1e7ns/Hvuqhjx4EkCilJ/peVdf1CFoqU9R
Hcr1jb3SMVPykXpvsnTVZpwwCCBCLLv0Gka77bdYpOGDJIO/NkAYgUfeWUeOUkIYbetJBzUgfBbu
fISd3GeTXJysTeGbqhQF8Ya3IPhIqR18swhwDysyk2MEr7Ut8bq7H5Qas9yQgWrS2v0FQEj+m+FP
+IouiAZ1q0lOYKh31KGIRKnw2h5byyaxlJ3Rz7hX5CHjXVkdGrP5hafgPdfWk9eqomj9SeE23828
P3MIi7nxkmT5IHUVMebufIYMR4ijbolh6ayxwdPRp2bDf6kcKiPoeNcF4cJKnGkEfCFgmMW2UKWr
ZScRk5GgnxDPXxCrZ2e/XiMHcpEmH1a3wzXs314GXxOPem9wou6ltEnVw4O0DhC6VyLHQiEGaL7a
6ghePfJvzqhSHeHQTrNWRLBIjTcf2c7tyb3MZ+Vm1ntTfwbIPWzzKBrJ2feo25Zq6mRAjWBbeY+i
bd7ywwnvrb53HU03INRMro4kvBYA0xExIjx3VnBVfDdodqwG0hUYo2dlnSQDaykpyAQNCJgdFp8B
l+gmQzBIyUUhcwQWH4IN0ipUbgFntNnKe3yrnBltBqW7iFp91NAsYeT7IAUpdRM2D9g9XIN8z8Bq
oLehbmKy6LHfqxngz/re5mYfmKyjzgoG8Gs79VKLj675X7J5bcXrtn7vUkryc3LqEgufPdyc2/RB
Nz2f1UA2rzCG6G01Ju9o89qx1VvQlG5Bo7AFkdsf+qkxCufpHnp3/q+F5VvcgJv3hZth3v9N9jzL
gCbJ9pKejdOQDnXW0wI5X8QY4Iohljnd1N3yJwIbI92u2zQB2Bfm4uOBPbdz8PGLNRq7yeUwhG4c
wluUpchkeriL0+PwZqHveNNE9c1i3y3NNM5HV/OeA/JIbAViKsnRTAMS+B8sAV0FudDqWZtZblIS
9XZMoYZaLs1gPGeLHbS5D2txolfMrvopo7H5vIav6S2k9mSCzC8Zws1pS9tvyHLJpaSwx9FnU7OP
EZU/NlAoVZ5VJpGyJHf3EQI4CtE3E3ynIgF5TOq9N+NcH40xOgJYIJ/YTwEVhXtACR/3+qdGoiuk
NnD4FgKLlf9eqbq0XsoD9TV+tdFobNz9XgGEtMB67UtbU5hHelUXAQP5eAVxeOF8DSrncpdfnWXZ
cOzzgvlRs1DKQd9Uk3Ji9KghpfjC57PrPkyrksu5OVvdAlBbtj0UO+y1mkuU9VEpMqzMTsI/pvgh
PPHyrBZyNPm4l8qgx3w0t5+IDgHZ+RXMD5AeJPjRgbAxzwvFmdWpfS3kGXhbETARYBIk83dftYrc
+zZltTd8ONmAhi89z+YIKP6hoB38T9vwxM8e5aE6yZVm09JYqQokcs31Nomy8F6Z5/mBBb6w6ipv
i6nElwkFv6Zoi5EEnk0Mcfu9pp6G7Hi9sa5fGdtTig1cNUVxOuEWp2FTQvQAbn2uXvD2Rqpr2y5z
IFYr6mgmzbCZZ7FGoS0za5mOWNH+F4fayffuopok8Jqj+xyIODt7R37hbYhkExYZ9QACq6qKK4Y5
WzHjksYonJfTqhdOFe3vSdgILNz40cN+b7yPDV7eIJaP0dl3X7f+1JCDu0CbbBy3han+Shfuq0fu
KDeTbIbQ/b97RHEGtAt9IWaMjim5f5t4jU62sFtouBeBASHH9+5TLYjfuhgGVH+A29/uC3bLCVZu
D3nUNkMtgaySBuFILtzFqOBLZTuC89iwMie76Kk9RHdnak2f7090ELVWAv/MpDkmHTcCfA5FTetq
XBFkFSk8OFJL+ZwEFNxMFXoRZWgDgEVKAWgvKvavwEDe5kiFxsZnviEdq5yyvIRwHJyIlHRkSrBP
6+8EuNIg3y0tyvGWP39b1u7C+5KkD9FbjuNEe+WMEuKrgxX3PsqYM/HsDTbQatjCLpDnCUanLBco
7loq/9iNgIXfeh+L29bpOtO/ZW3HlGqUrel74J0CU7JxTrdWvDLMK3FJiz5vpn6Sz48ZheQDva8M
6xiN411rBlC74fGnb41KpPHfrsQ3rY2VRN/rBfAcAdvYk7DVkXTyAwpgYpJAZG5gaSGeiBpqADdy
9Sy8pdtats9KcJ97ht+59DPXELYTDeMPI3H0eW+BbFqn38pxEXh2rIJFGhgU2nGv+RUULg28wAlS
AR2wcIJWJdOzcX2L6IVg2884WK2GHyhYPC3X+s3rcHnj0C0YM86MvE6+aT7J/Ut9qexKkbMGVJ6u
y6EYlkrwslHpH8MXAdWHSfVZ4A5bvTYYXAZZn6SKLRORQdEB8pQ9sdDEMqhSheXCwztFtzsvGhMA
hvRB61yrsOSeAJQKOA7fWLIwPWT0Zpt+3HDzPd6ZV09d/d3t//wyHV9aRG9ATl58K78Gr6CD/JUL
dbDCaJ1G4AQn7pU7OkggQmZens1CngE2b0xuXP/GH67Gks2QDAwwFIJvWzf07SAl5x1vyZ+Od6Pj
sDJyNqQXAjBXnDKBnLZBIAgLFlsPCcXbObYYIQFsQBmS/AjU+wLUJk/jBxkPWdJRxACrkPAjvYdZ
vfyPbHGY/7ErD+ID/Gm5UR0o0uEfxkBzLSfOkjeNisgZsl1vkFwuSts6MLUzbuKX43P9jzE1y85g
8bk1NxHVnTfhKQQwJv4iv0rqJc+Ewkg0NUCU0xTzqSqUbEocQWImKu/tjJWJSqiOsrk+0fWgCbdE
TCIh7Xw0S7BHuXPwXfc6uFC3i55F4Dtq1Jkhjtt5mWmueQOMBFPt9KRWZXifdeKgbnwLiJtlpcou
RHbVvxYldyMJjcZ72kXhz40CEUNxvdny4XEU3VfmQicVPBqoL43GxGeMLqaulvg5iQ+f6kxywlAF
lqyR+7KoWdpRzfenhljdS6fvafuVasDFaY1dv2GHWJuaWyl6TM4ea66otluhwnzujtcjgNlOeo33
wb2BE8xhX3Xsi2bDuHZwnnsjRYp9m/sjVwTWDqKwuE2nOvIqPK6nO8mamT7LDx0t0PuFHW54LGjR
F+VObtKOKrD8Lp+0YdOnxTeZ5FdYY0seUPqsTKtjwaDJCXqC0YceEk6B2jZ0aE/QarWTSqMajQOU
61hb9HFh5FKrKXucdpvKAyOLn8epD0YcTVkzXtiX019JdxUH/kvesdAedS7cwqPwI26HlcD7LbAZ
A7bwtxMqXTZlfbuUAhnxB4LGFIghh23elt0cNWEfW163NIqEhl5R+7ah8woRf9lucNCV98guutIU
wDCVKxJyJeRkWbIrttFjVV20poqhxASOvPIwaa9KQbgvK4LV8Dt1aBEctk0dA3hB9pnL7WLzTYzp
QeJQ4uvR0c4Ggtou6B6Ljq4iJ2YqROnBSHGAuMs0WObGTotgJaXGqYzXY0fo0y0CPTKgjrNzIVty
hNvBgsVOVJQWhKqKB0OR89V6r4Q+A+sBXTlqkcN0kAHbrwmp0pFLsO5Nl37k/fYnVIgkNjNd85i2
7mSITHYZAZeqIQDQJGQP5pGQvifeGaYH/xWQboBRXbXUnu+OVSKbKkFpDgEiQoiR0BtH/KHNht/m
VsdTtzp+SrC+pdecN/u42NhPXIINopxuKUAahIjgnnwi0kj3MUtdQTBj1JKJDuy/kkbkyjmpEz2g
viJq6SpReJWIkH8QEL1LJ68uGCmdsX3nZeEPq9WJrB2/NQYUHokiD4fWO6J69eZx5kmCwvqYCGUT
TE309sapLBguQYRHoHQuzmeDCwgpI4fKNFPOJ6yOxuwMroBYDbkAooAa54owv6rpNbhu+vWOcZ75
UVvn5ErrqX4hhy8tATKTifNBt1pezt6pxXFHyJBbUrbRrAB2Agw2ft1pRwT5BOQd3+MoVBsoQBC3
98ZY83VII7Qi1Z3+f4V/ePnMejJuMgstzDWI+mqoZJ0aHiqMnFoB7P9Rp6GHRdzRunAVT62eAk/V
CpMmL2LttY6VW7QSICMuGpSLizyTYL9ykcgWlJHSN+eDo1EkTa0SfNf8c7C61EawUqxD5dfJ49jY
m07G4F4HhyeroROikSI1GKZV6bxU4GxiSzMIr2ym1O7O9dz1rnbS5Kqyg2iUvINxoHq9zSLipRAP
YTZabaTumSfPvVz0ok1BxH7/agKU/pSWhAL6kzpqaOcBvNUl7K2JztVg9Vp9RUD+qjyn9vyI71o7
Wgnkp3j37+JW20RpJJMM91l1yJ16Gl7WBtr3NcxQE4SjsvOKQhLGurom3ndlM3wswU+1lxSGvuEJ
nxIfwc/Da24jnS8FwHiTjWi7hdfBt7BKyrYz2Mdgj+Js8bsGTGQZhwmPQoiMUly5BvlF2FqCxorf
XbJYFV9+SR2QHvTZhWcJ6RKsGh2wb0RZ2eUVk1rjkQ3hVuDq8RisZUxb+LGVPh666j7O4AyzPpfv
ZvXxFP6hBbFVtJeBbyYhiBpP+ozIrRgJ16MVjB05Qq1xaPr5FZTazYS3pWzMWcdrufmf50Dr+OmG
97TV6Cbe0uQ1kRJrLtYu8GrxNHtIJNOMQapbqPc4c3cK1cPTjJ8XMtCPGsprezpjiPIflHjoNmZR
JPS9czFmGdPkHMpkssd8uEMTF3Uoe4EvYiSt7ypRrawpUFlWj5WpzIm9QHnmHCYV9bhHNeg5VXGB
J4dMx4cJXaqEzK9hOes+RtuBj+hKL4pHOJNOYhD1sj9WhKGebB1G2ScN/8tP/I94iOsPHv0am2vG
VLA+ycuV0J1CRM8j2CgjTu9LVqNy/ReWX8ad1DBscN5lMNMGEtoneE1kEPTSwGlRN1lgR/i4NdmT
3vhOm7hUO/KK/lOv05uURTzIM7Vzj51l+BpWCUNd2vwUriMoGZNylu6JEJCIqiBMO6RYjP5B8W9+
cb+JUW3jwSc/SB1v5k9vCK9AybUAEr4q2NC8J3sFvQ2oyRYna+hHopT4PION+cj+DNA3O6BcRMI6
JKLyizHz8Am5Rrsi+d8km70UQPZLT0CaHLRTPQSNrUTvYAjJkL32wfOOW8OmD4H0e8xjlrq7nBQm
O8k5WQ2CBxj2lckYBFCDtdKrSObg62uToEgF8eOpvbJJqFkVnX3YaQctvz8I22cwT9KSCdwS52KU
hRBMXMdeY/IZmhepRVKqSAD/lWcRa8G9t58/0iTfoF8Dt+mxlpunB6om+tkr8ruMx1Q87z5K3VqP
Qsdr518gSrIgMQzU7C4eS18kPOYq8LsYzSAPciMccnTwt4tki4Nu7gWIeO97oMRBBCbAH0h+Xrzn
tfIrhkQ2UrZEdeScZkx7FCL/3Clg74+yzcAKLMNmw0Po/IlUDniezmTu3ZxSnOZa9WzpnsHttXCR
qL+nbaQvhrvL2b10TUbcLrogNJG/t5vYcQ7Iuublc67dNOuL1FZHD7c9PyCrH0FKE3my7DBYVJ7f
nI5DwUrDjtjnOGsFkMfIIGmba7PfL7Ygt+gMaiXVtkjQEglKxN16t2ZSvLkXYJv5qZZVhoh5HuJ+
TDoIIzFg5E0ZANJvsfQZPzYRqEFN1gt7xB5o2DINb0T4rExWdLwqS//bBo4K0BotyfzRdh6Ski5Q
UoRi/WoG4B14VC5GYtgK5quQMvJn54SaIShJhlelA8jenidh/sYm33IQ/rZNB4pEK3MaYM6JmnqM
mvavaxSjFNIzMJdd6L7Zr7D5LOZxitbt5gLXN81YFnfOL/1ek5iOBd2u31XZIgMJCIDGP/PxJMpk
WibejieojGl9aMhWd/ElmsLdrBuPMzxodc1ORSlCUI5/Ol23sdNozaa2lwZyVWYFIBqLCyhSaxAu
YvVuf0t3LMY9NAhHTjagQWPO+iCw1aXsDb0ilUI5Vf/Wn9mV8dbaBPLWCMx2bRWVR88sAlLMATqm
H4R7MfkDmMiJoEDRyWjHzTe6sFIoCIIRQLHyh919WH3KLB+T2iUO92XMy/AdIPoGIJPFryXxcFTk
gG1AmK2tygtLK+Mf1WH1yvCk0MKGzYX+BCCrMuWuENWqyexDtgx9eEnBtRYfTmULKPblcVwbgKkB
bnEL3u4DtEi7iiBt83+GtdzJubE6V+Eia0N7n280KbpqQd8piwBrdLQ0ejuYzYR9xeP5sDNevjmx
z+wXxfzVBs07CxeaWsCj/m8yn2b0IrU1nh+RWt5aPXBivvT5w54z2RDCliRbvwJ1x9RPOoKv/HhD
LtjTM90cN1u69oKfy4EWsyJKLmF6Eqjf+Xw0SPWRucwGNeOpgzBC+usjNex1FZW4sR/89kaQI+CU
EcB/ne6lmNGUWNQsQDTY/96PZlQg7ZG7kzhWAnAlyY/Zt07usKEn38gvVlC7bRdguxNDOHpvYZ45
ywYY605g/ZxBdKwmFkYQcpPZz947Bm12mmJ6l56cQh0MR5uPiWnc5OPccl/f8QArmOZiQ5nqX8vK
cZavr2uXEp44M4XW2D6UAHP4Jdz76fG2aExF3HiSbd0cDMTDmNkNhDQ2SGB+1igHqGVXP5ivzamF
c2sKffUDEjWFiiUrl47EmgoppyWIZIKjSZLDFFNfhXn8CSQqrdH67Irx09mcRIFkOdJTR8wTQymu
o/ycZAsVo8i4mbcYzg/ylLj+TNQXWgBK9zeJt6B8WWgPzk/XP7JDKyp3zMgMPV9UGiosyKp77o50
XkQ18AtWrzMMMw++B7RraGTJPcNkBQQkmDx/UBDXILfaLNu2A50+86IWEcNxR4JJnTLGKzIqJCbq
wmMVnTLjdm7PN05gn3XaPBzu1eyOXXrkWnGW7ldt5LBjVQTvSTTcgso8xMMJtlprih99smVjgTjV
myfkVgOTdpXappzPdAUaPrvbml9+Yyq/Cz+qv+UHyjUhpxCz6ZpdD7ofeDum+v3h3Prw8OvLLoHD
TQnwJxkARbVnhHvroweOeSFbIuh8IY8I3Pv5pxo/Sa2fomyi8esswsPto3zhDgw1U4GdwLczoXzm
yXQ1RI86pnPVEX2MDZbUJ3vvcqeO2JC/8/BV89LPqiBPZDPUfBSryqwAWt151OlgtrKZU12Lorcl
M37sUMnLEs8mVhYbFGNriH7YMo3nDk0yz9TdLsx/F7lsfxv99SGgA58CE019ykJkWqBcE+oRzIvt
x7LRJvigM6zdykdFM93a/uVKDNvUh51EnqPbTRk47tYrrkyUHqzzbsPERNaMzkiv4v40kBKMg2XV
HnppG7EKJpTa+Lc01CNAdBnZHv68xBA2jgwchdOAEq0+lbIX98gxxTeOViQ5MViV86778t9fA21/
jV3Y11MM3UJ4yFqkZG5v5zjL+RjfAvuMLJfFUED+CXxmeIvR7Cz1+89MkWUwndUKHykL8Kin8SY6
oYEe058w2lUSxxbxfU5ndvvnBdu7XrSbhfbUPqD4fdRJVnkn9xNJa0FhdLhttOOEJ2mchILGLdVK
gayQJdLYMvFOge4zlB70kbxgjpWDRarKoO/xED7VPz0RxLrXb+WfXO3OVaU82z76EjxaKBFWy9Ce
/O73pZVRs7cguJy2fMAW0IPHD2cKA7IdxZz/nrjwnznBjLYd2L9J1kENzymBphzjdB7v10nJSpzE
CWhqym+38oWKnp1daz6UOH79Ofc7qefI9d7groodbLx0/658g3ccjbtG/VO6O1VY+9JFJ2gGzr3j
TIdNO9ZuZ+wGNVXYZ0aN1kgE3EMdf64eb72oJGPaz0N9uEx25GKvMiDmtuFUftkvkMtyhUgzWBJP
ijjmWxslNn5osAmYZYQ3SxmNTLXJRN8aakE7edCNIEymIzTo535zgZB1RfyK80hc15Dt591bqVfD
Y9BMm9uHaBNzImuza4geKXzdmLlkIsLVkuvUlFIX5EgXpKoAqh/YyByOPhUnBAj6m5SRarj9IMp1
2CMQ5G9EilzGGoREh7gppWKltJVZcW8OsZG5YlNfbmlIW8MPCtztIvhQR0uE+2SZKL1rikwFZWR4
aTrrf94IanJx0YpQvyiqXbX6rVH9krJKkH/zrLQOHUYfOm12p6jrHieENYe2yQP40XnLw6oq+VwM
kt64as6Gg+AvwtY3y20R1iEz+6bn7pEZWMTwBaVDFUoBWRuAYdQQD0JS2HDI4mV3qE1TNu0YFuEw
DTMDWwZv+8qzAj+y0agkqq3z0t+YCPeYTNWWbm5e4feTy+loQmOEtsrXmcysoPmz8o27kf663OLt
FjBvjFHFlfaR2fHcfArEKvdFrVzainelnfALDkkpKqvgJxja3VFIJuXEqKbyAdjNp57Lfao1Zcij
JsS2Py4kGOTgiQIGqNYFclqIPaMQEpfnHza2SF6JqY7GJojTP8RICjAgAvdCW2Z/KPiCPCNad4vm
wxioYCbu42UfUFVUVCNyiEVHC2T14X4idE+upeyk7EM4am+tHetyMI+VOhLbgwRwVxDep4E3t4XA
93JAKHlO5AsPlrL6bMnzBBiYWBWW5Z4FadcpYsYANitcYXS2Tr72/VCyHx4nGu0LxyV0LwuMBP5C
wM4i+Kn48Aqc7GlxF1iUo0qZSfq4iLOPavHrrpk3EwVwemo/qk8j0jqlXvR8FyAO73BLE4VUUVZU
tc2rUek1ZL7g1359H/yphrzNt7Ym47ttnB2yMVBUhq6nfdCL53QKchbvXQBrkJIasi4MnFqeCq/K
P/xXrOy3lKojEY/SIOgDD6G88J0sLYqF4RXD6SuBmhhE5j3Rgit6ZxyShxTPlKD6nvntyj4pOjdz
tAe2ZPXbwp1OXy1mXUFcl+UNND5nHe0VyZs+1sNwmO4zC2uzKRFzzw0kq9VrzLLvc0wnz3Hz5s6V
EV91IWGJoUBlnAWIlLxeld6HbuVect5vfoI9Un3o14GuFGz4c/ZEg0+8BaGp7cKISg/3VQze55Kr
FluQ3cKYrkZUelB6mmTYP/yieOgxcAJX58GTXgIcbNUm+iQFEIPxsWxV3tZuOd9Ma7d/st3ZjoU2
kHzdX6HxdS2hzUSwRqpEoVDswqgEk54MucF1v6/xWt5vPBjmxuu1ntRIL81VpcPLFbknbZlmb5RN
7/T8Yk0sT8X0MQrtOJ/iEkdtcd0IfgcXYu8g8kZtvZwR3BTnEeJIc95Al5G7Dea/9zlsw71pOfuB
tW+wPHZZHJmTAasGM9yIRVmB7IUDkM8lI1z8qs81HNCUc2XEnx1n/VdNw+7fkpMK+uUATtz5iYvG
DL+YT9drgDN1pxOOF6rLCuAlJ4AZPKIgu+IQGJt6xTpVjPFaqdVhRRY7kxYBkOHc70p0uxj1J443
5iLBrHrkMKuDwKrx7OkbvunAi7emsNz7sGMsTCiEMK18eo2R79b8xUCJ7LDiDT+hAWArLKUxNvhi
bcKbloNXK25UK8W6RSnu+NvOo77lM76+A2wHZJnSubwag22HRXkf1pyhg9ICq+xS1Ijm4wrf5fdy
745h6OEyEhdEMMfe3nL+00HdqL0Zee1REFj/vGNyMYUpPm6JgyJP3R2/k5JL1f3Cmou3mHw6g3Nv
CjK4GUAG6A/i6KYsl+jx9nlBqkY0wVT/N9RJjmNynZU7IsC6jf/pf+jv4TM76nE5rsBJVycj+aSb
5iq0/sazD5pOthUbCOH9uQqjPBGf3e/GarbT2VUxeGn9SgN1CaeQJc+7/IjLtwFUb1Dvi6WyrUXL
c2qbbYGUmz4Np4nu33Hi6o6Wk2aT1xVkbejrQq6ZX9rGhsFTgSbs+UwqBSUpDTRRGAnYNgUc8cU1
cv72zmRYD3dlSNdahfPVxCHMUhRLpdY2bbmO6WLXPCGLuLTu8Wk37pSlBBvH5Tio8NXUSlDMxDQa
i0EiAlPUyDRYPIpZygEXkwcNZxampzRwBB4BjNyTfyjziDEDRRXBnK4WxJNxRNjB1YfUHgrU15NC
mwCcSucSiyJwNtcDdtg5NGBcPJ+m81r1hAP5F0HWtXS+9oEaZOS+XtL7P7eNxhtOphxmJKnPdgej
ihJvbunv8PyIPUUmwegd/ct1HNfVV26K/3voge6e7o5jcQn5ZU6ismvMDJ436xnOO/Y7OrQ10OEn
FpF6Nwvc3Mc+mCgl2/w11LQOuP6VZgIVItlTq5xYC1CVFYACOuNFeJ8iQeK/8XAqO6mrHOQkA3as
z7OJsOEmQ8WMi7s3DHpkpNp2WJzwJ5YaHY0qQKEuVqb+mnEnE5TvtNxKK+aiLITAG6pe6BPz+Xht
W1Wl0acUrnUiXA62/POmHkdAoFnIlg/xhUz0LOiFZCLCPIIJ0rS3lmOdsjFh/ylrGVPqYfVYvNoL
MVZmViQt56VSuV+GS06uPoTunYQfryuugUdPT2vFkesHgRuvf1CMmKJqd52hfPAydW89EbbuQtsD
SyxzgoiHcEqhE6jB0SCwJmTE9SnfVVzzPfOWenkHwM5Id//hoLVDCAAJIFBVzWl3/7GVNoWnXBr8
eKOl54gIa9krHyrsx9QV5FXbzUOQrta+qV8Tp2Tp11V/9STVnZzjtbkdkEpVw4RsKu8uifcuYXEN
oYf91jqF+51PkORea5SxOYEUwdmcPKo1J91z6mNgCGlK3WgyrQy2kJa3vCAU8JpCeCqnIgK3FTdk
wlo/AQf1kcN8iGReA2kru1+yb0B7cHKZ55Ltrs4XPYhbftuXiwq4IbjIj6iwbRvlJyXDatzhSFwU
d9ndgZJdLx2Q/telv8RcsC9qff6hFJ7pX464X6i4Tlic9iDbUnUOKyVqIeW2X57G7tOCbbfHssAf
UnSIEl6p8V9Ph+83AHJSGFJOT0iZmXBMx8a1OQBSwUmvbNAOPdy4Ie2prhQiC3ycTfYQzRFsQtvA
cEwX0jWgZb1C1JmfmENrgPs+6Sce9F5+hyKMJBLO6suE3qM4XH0n5O9noh5iHEjeOL4hFDCniQhA
jmB9goHRtuzUI/1HBcEwnJ9bWVEgxe4FsXr/x4D/eR0u7XeuuNfUvsfh7ovn8DGgU+3Gtr4LYEEd
fuyC70HNHH4ndw0IzV/al1M6CNyeJ1Wd9suvuhlJkKqWxPoMeSptchm50rjHl0mCx0eR0OUvPUzD
HonntTylVcWz5lj+cqL6mBGLoh84U9ukotmJuIc0IRaqDg+R4iZ7/lZUEpwlPyzvi3imMLK2EOmZ
QSl6rfSxy64zO5UkHwOoNgG7DpIwkBDoTlpARc/DD0cFoRJumKQSmXSdwjdM2qRbwWANZ0ptQPyT
KuwykrE/HrP0m/DUKSqlocrObCDEm/9vonKQuQRpw/w76/V3xrwbK7y8sIwRCQHWRS4mqqyzOhd8
eDjugWPdHMu8Ympvm11PVANAPi6E7avg2om3Z4FjDjy2Ea7OWfR2LOW5OtT3C1R/NSRqlQhPGN4F
o7timRGweOkbzySRy084bHT7zGZGS8+NnJpvkhp0wDMJQ1+nHMHIpnhmqnlmjJUJSIRddT5te8UZ
RPPFi8ByoZX4eeRNn/bmSmFdWuEz0Lts+JmDYjkEwKau1BrQzTl2bF9Sw2WiVJmNJWCwjtUbZOxO
sibWzNeMUUB1q+f9eI/arZTU7ucIopkDsMxuSoN/0HQVz93LrEtVvTrieZ0Ji8kXKn/NTz5KHtId
IGnr2/xdAKHp8/Z1mNdRoBvm9g0ApKroIHGhoIucy/dHyzEIDx6KVS2qGJ78UFu8gQ8IgxOuJlkK
aDANE/W1N77JS09hQsYPr58qavlYx50TRbEGgfhVPmPddstSn/Y4LbMDK9wjfJUjie22yW/+UGsQ
LywZbSNk9PrE7yQc+j7cJ/qCLXAx71ETu90mvRRGpkH+igiGSt4Zxi/1w9CdqCx6qjgWw/kPfvjc
G0/eyN41+aSAahSAkykz7oeHnSCUXwzffyOyYmOannPMRWcnACOICYL9xj9C/3XidKJ2jbPJoucm
zC7zgA3ToO/BfonVYD3DzwHloihKPIQIKybvDw77J468g6T3L9Lh/5MnhEH4Nn+NtDAI70zckblm
7M9HBFyCvAwszY8YQf69+b8SkLPmUDbzjADKs8veD0NNpxDh4WflFsoi4XOnC2NcKKChf79zG4aq
zi9ag4bZka/WvSe+OKHDkeDtfTZkMpF9usWb1oEtQ63GVaaD627et9RHYSO8vdIk0nt0DxwaI6uO
O3NSRzmqSI4KQ/StvVz1Lrh7Ba1NRM1eLXLo/aPdO//a9sWBFfn3DqKfS8w28vxeekC++iwGEHdT
vw/fPJ7YZW0bUqg2yyxiisY1GR1eSaWTvZVsrNbBn0tRYH1iqm0vfK+i0iM7ITGbkUimxgnPFkm+
LaNCSa3jhz/NDUfqVwmnec8okW7dDiPsc9QbWYhBvS9p5OOl/YClFl+k26rYYdnE0mSPakbH7m0C
dLHZuh5UPhd+ACGGdyf7jmcVmTb2ro45XbiyWIw0a2unOU0JBdPQF1mZV+nPdlbzvYuXp+E/xSgA
Q1ihdi/soxJ6Sk9IpzIbPQ9yqKDY+GbqxnHs2el1sg08srMpr5RHXJY+tjUMWkjhg3t+TCXLvrD6
DhswEW+CDobyK3PCuKXAzaoikDOd/1GF3ovctyrEqa9J3WxZVDSkJ8JJVIxwPeWGN2Bfet1fqEzr
OghcjzlbplTaYlJw+FvcU803jX/6l9iYvEwY1vKTVbMqBGdDhRmSOwXBJBvYAOX4imaAAVk8LjC+
sXFdZgCjA7DJWtA0SvCxooydCh9CU2encs6WTb7kwiMmW+XYx/Xgw5mjxH61EpbsXw7CODcZ+jkH
K0RaOOcPoIBLKAddxMBs+V3qD6+ArNpt2qZn0bQ+KXJWQCrJeboUW2oUBNm7fORJSu6m0nN6eAr2
V0TCU663fAfJWTXY+CFzzGjxKYA89qQziWfrCmuNoFUaG2qTdqo3fIu8qzmW4T2NqHM3uzcspU8B
GG6UCTE+ASkU386Zpg2mJtQzXgWaebL9U8kW6CtFMme9kyTn4VhJihNrPNYl1rc1RL06BmGvu5tc
MTOQ1MtJvM3H35rTJYwnb0Qx4s6aiBVTf6jcFmpyn/fnXRkjekpSPgo2QCsH15mgvUFj3vA7QdRH
pCRyBAakmD+odHQ6HAuw6+g5zKJWcahFmlTM2lTgRB1pgakw40m96Xs2yeaaXX3WS9IOVkddP8I/
IFk1xHcLKCDsbiQy9VhzKauRIRMfMrYL2Rf0rQx5W/WkQ68kgeLCXVN7D3clgXvuIoZ90XZuTU38
hU7aErfpT2BObPM3IPfpPbzffR7HQ03rCC/7cgLfU3rwkF+SU01Nj12v3J6OLelZRNX3EYyGjdQK
aPoi3AmYO9mC31xjHnkM39qKxobzDI12uc1MxG76tGwmWQYEVc7vMWY7nPJ2fKtFTcZKfjw/Oxqf
P7hzsGwYnvS1V3L23rbXgVOZmNlOkbVGytDxDAJnWw0/q1oC7mYEgEEVOICs07xo3o7ThJjU5h93
VjoIOZ9aELx+FahdZ4zJ4m2YOLJLjcQZTmWzCFZmQ6NVO9T5HnvH38S/dLFmrzAbyvtcpXOfFn5X
upOZ+lNh76pgE7c9oBvrVcEF6qI+HXXftb8zmFcBAWq5RB/+DhWyybJWpWrXCLVf6DMxFW1IppKV
doXJsdu5mUiQhETctuCOHVG3LOKs+tn6VR1y02uUiomItTYYQsOD2OvWxwrpoqPiwk9sJT2fziFJ
TeYrix2WTOlYnosxgJyy1JqZ3WZsusrvWki/FSyxKYzh++LpzkNd13WX1hK5RBlRRmmjsrKiUVPU
+t/os5HjnbNQ8IwtIcCZDk7T3XJYenNq4RkOgPIpD/ASMbmIcmkAHxium+5nWS77RXrpb5uiXYF/
S5PYaOW0Ruw+VNIygLbe8NfkmBuy/zCQK9JUCsG006elaSep6IQZRcHaPY//zn88mO0ctxnPJtKS
mmzNH66rrCaUPPnZHhtvEcZGeLp2Ydq/zbsKBi4FWXhI6xIFvg/Uru8aQwO65efTmEGmd7FGNn8P
cEKJXHclIzRI4wDs4n7Vjpi20d5QdZ7BfM7s36p8KjgcheWG+BdV1RvJCQZeOXG3HEz8ogMGaYtg
jUo7sYlUL7A0JB9r5V+7wYLMAzeaAOjvSrZdkO2fAyNaHyEXHpR2qGLcyCsyVyIbFwepCsGUV8EF
vYCw9SNLcuZBbAhjl26JtcKJM+DKm5fTGRsPDT+xchsiDZJJI5BQqe7OrAf/A5m8xEi1LAfArGUc
vv82w9sxeZzLtWLzEhxuIiq2JpcztN10rd6YFkEgaSwFesGUhrw7sXYCkfx0O0/sQkP/c4y5hl/y
5+avUXkNJby+ZJ+PHgnnu8t8hc3DRqitQVyhi3TIXY3U/UMMv4Cr+lq4nxaCE3zf9qsPxnt5Sn7g
ocDyoyc5Ff29zjt5B59ei3eH87ZCp5R+k4brm/fKqEzeTEeXVwyUx1rBAV3rtvPIoD+s91Y2IAtL
IRaFV0EaSV4If7Yrht9lHoX7D/y8MGnO1kASOdf5X1zS02ZgxefTgrhVxl/yasbCTb7+xQPh4hdT
H9zs4Bc1ylTXUqlFgf2xOqDehDoRsroaAIW7aTmtYLE+jdrsrOJzadQK/VwFKmwZFEk874FVtyA9
8rHHqspu8BMOKuaMlx/PcEiCPD00hXeAQKihLkbUNYbbX96ZH4d7DUykzIcFXgDEO0wP3G2RtXf/
ZwByTGGV7r+o6n5w9xC/LTTbTWbeCTSt+/5t6teSNRPxDKM5X+uF3OfMjtHEUxZf2Q7Cxihg/G33
vwJX9HtWCjk8EYaVulc8EHpeTHvX5DYXNjwCnILTtuzxwLSXnr1rObZfhZIWaC/yhyLiDJ85Jo9Q
jibCMyEj8SjUYzghEmEX/+lmkdArnSmHuTaFUX3jtYWnPSo2TsGFnwkVNzXYsPywSeNsGZvnQy/W
we6KJBQLCRxQf2swMiZqPW6er/UC20aN/1MYdk1qZLs20ctvj4b7FhNfVdkjfhYhAvdpVIRRSiGR
I0CAToYl46JUE1RpcTpByeqZAYwLbtiyzaZe9QbG73v4TuKfrj5jLytGDnpJBc7j2t/XfwMJotbx
jSL0NJTzptp4PA71QzhuFtlQhAnII0VrNKuC6aQthykOmHMw8Rtm2L8LZEhlZj1CLLYwJB4Eug4I
KmQAQY6W130KXIEjTJt3qTpfMmgiTfZobl2G3HVF4gLrBi4I6jp/7RuSpHr2rJ3wks8Vlcp84jbr
GnzasRu+anatS2IXL0TbQXq9zX4l8rZoAFXaCum9YRGau02E+iXT4MAYkf3ofx3HeE6EHfA4T0yS
69zq00SO5ZZOner348RyL/kt6xJcrVa3F6uoF1eB/uwAaBwhc0yxNOvJEP0+4G776+fnfgr28CTq
arxysFIIj8rKCThu4sDvbsATFoEahl4KHO4wbu7FcBhM0Wn1N77+7CBpMtnXSsyDsFueiREBhez1
BlEv8KDix8pjutWMZg8G31VOn4n5j1QLqxi74vhBVopde3oIQzT5OLsnAgtBh3Rg7SAsbMqMpuqT
kOilZN6RF/37iiLQc2e+b40GhGPKZt6+Aj5IFK093ybgdNxQbRMZU4hM7onKYdr7MtxMb/LUBb4E
k7dmFIzJJopVMxLw8DevXwI8FcrXo55Bf7n59VYyN21M+5bddiYWGDh8ce64CJSRBBUJ3LjKfmvG
vuqy5mZuv62MDNjiOznn6ocf8sPjSKkyll/WZjGC4HW61MmKQrZe8VsHzMEXFnNWHXKjor2XOemb
cVlhSjteiB+Ze0XwfOV1Ff9AtS4TYGVECeaJ667kltcCiXSuJgt4NVHAOUht6SlzWXhbsXDbE3uQ
yGG2oglVMqYJfKrLRM0WsgJ3Jwg2tsoaIwxLjTRucI/9P4l+oYDV9FwFCqjV/w3GFzs/+yY5glD8
fWGcj1cK3QeZyYkYfR66BZBCURAP/pdCeDALOrOfuDwiIVyy3I1PI4zBAnkMZOfgReVByAF7gP/S
o9ONonQLPbFBK0LQYdQpZnyjXKyI4ltvYDRz31wHmvFoR9BjAZussBWhQN/zZ3MCMMVRRsKJUcwU
q6JIExoHRR6RvzRW1q5kpu1W/N1YWZdPOWd30aiWmhAwyRoJFGWC6G07NRshN+Hh2Z9vq6Tt2DCL
91DIq5NpliwzVGvWc/bC9B9dTnN0GZfXXUGFjIBycM/7zn836wcIhjYumJ2qr7LLwEGW16hbIXjw
9/kFax6jPrQQp/biBt6xtmECwGUpbwQdrvs2Df0VRRTziIbNZWYUE5H6Zz4i2kbuR1o2q/h1wI5C
4oUiW5VVbkb46WXZZVEhSBM/J15wEL6fxPz7uoIhz99hR+sYD97JOXvY/T6WJdj04MYK0r9b65F5
M0jknteKJkW/JLHVjIQRher0j/UwSbU/Q69+Q0p7OsQqFuy5vMgTmtBmjgie7kdOGXRk+2jpiZn0
dvhyqL6/q9xF7NzIxMTFg7aNDR3YV/Sk71lP+vyRfCU9Yx9VrQan3smxtR2G/EhyZHTelzG7ZPDI
Vn1cQ7xPEXIkV3/TX+ZP9CiPHmk9EIcBG+youhc7YneRdH0arUWnCLLoAOI8ILYQbqkVMnKRRa+Z
VeFcBhUBc8M/11RTY9qfBQ6D2tN7Y2lQYogz4ysqzb+kFTve9PpCJf8oBX19kQl7Kx3HWSpNTB7g
ByIM1RJ63JYmrfxJTTNPBBdbIzP5b6ysT+VYldxixEWu3bdhv0oWlogFh3fqDaxOws67v0zTKnTo
j0xP0YEkwODl72NPxeNM53bMWFCDuL+7BzXpFbjugcYWczCeV3jPEaAVg8gde5uzFszK1QYs69ju
f+78Jy3mkMfYujG9DftI4OdSLwgjldb5IoYnqpdMRONuRCgT9ZAQv/LVwbh/NumZttccvLj8L69B
fbwO8zMfFt396UAL+uwodpgzuygLq795okw9e8PeCvNlVcPUeenNqKk4ocHmZEnFOoN+a1Cw0FG6
mZssw6BxskEcb+zvLI8VVVNNrRF+Bbydm1lgirEeC/XpR6yCMEuk/wJYpg3TN69sxaXDWsjJijQZ
GIkcnT8r44hIanwdc2F2m5FbLGEt1Su2H8gxNuFBep1/bqMV6XsgZvtietPsGaBOEP//9u9TFtXp
nd4lgDE7HXnKsDvvLivI4O/Xu0troV+3xi3jDNfVSrjpctHYj5htkEm0nsvMaIXXDUQjgaMKwfOf
d9D2Pbi7gC0CTDBoYrpEC2OkAGpkpXZa5EOH+b5ojSIof21sZwmHfR0LppLI8cFxfXCGvLkeZi21
Szl3C8zpUJ37eC9kokJUKjkoXmncByR8Il6JptDpkv0nJgukNwlzuBWyx8XZgWywpW6XqAoBRp+q
vESJ2ojtMfo9gVWrDGbH0WvIeFiicslB4wliU1ig4onbNTCVRkZP5XeAs7mDwnJyg/qwQsrAQ5ZR
lKVxjx9M0TCPlXr3BxcErLuu4j7bLRbr6NzEPxr9QTOMMOOGWI6dCK0g3xcJTmi/6bGIAik3mRoM
WBvxtSgbT6+jVCDwN1irpKN4IPXjk9/XVjl2yYdiaMDoI1dZaxJdf3lDB+oT5gFdlIuIUEcI3kwx
cbFWLXTueYVo23iz1pjgCPYk8NkgUOK9CTHskpuy7VTJqVGT790xhScGQlL2AV1j5iY/KseRjeU5
CmLg+fDpFoHB5x7Dk6ra5opihMBGsvWWiF/Ebkibj7YTxfIJc+EMDKM3TH5mmL6/Dj9y63f4MHrR
Z7soGTtGqxz9hXy+4AqEPwppApxejF5NH9A6I0dyzlbPH16NaaXrVeYAlcBA2o/J7k2qzkEPnjvT
qMimjv8hPXn22KHG737JKRjvuEdMlkfRxLQ826UmQtOLGSN//NLXiW7nwVP/CByzNd2YzTEaFTiS
Ia59ks7Dfoszyq5oakxkh224WVaeKVYS74JW7Eorb0BZhrvUQehpwW8qDNjH+kr2867T1n/FzDrY
/Zh+fIRLf0Eip6Kil2OZWSLfZYamH31K8uZGrpDHl1QSiLtLnpqsa14X42G7pe9tdhuQ22X6TIH2
AEuqYhKEHzL8aSzaIbkNqA914tMJwconkbHvfuXc0/ZgxBBdTnzmyqTf8HZozgJViWoXn9PGXl7N
IDvKi+aytmnf6u1d6k4XJi44qN0ggJ1Bh9pSdTXVcj2s07sgAzEEADvY6bE/KWM+CmpKG8BzX3qL
2kMjj6J++8B4e5hj2RuaMq27ZTluqJolrborw6XFk2r7iqNbbxXEn9et8GlajGa3hq53cah8aJo+
4SqXn26gffP3TqnYg8+y72aGYhVV9zS9LRk/Z3QTjTstkEfsiV3/m4nIuKZ2SrQwM2nJ6oQmbYVU
c+RJKMymDnlJwFMFqq0A9j5q7GhQJkYvYLgaIEMMG61JiAKP66TAnY44cWoG54MygMuJYzSrdG5n
drn1//ZvA+6YZHpf1ABWW9qhsfmCIB1GNqrAE6rvQwhU59qpzyiguPmj3P4SR7TuMUNck9WLdxie
RgV+Hb3hzL4Uo2YdtrjsFBF2UIaEMKLC6zXt7IdXlQwb04DHVJQs09N0h8nY2RXW9YjWyCgl88lA
mlxuFgP5gQiVQUN0mdcBHXiVVmJtz5phAmPbW5cT9Ym3txacWNf93amTuYruggZ6pjoapfSD+2C4
3bMdyQb5v7DlfUbqxfoGs9gyotaFlgCXC+wfGueXEHdBn5b1XCSoz/rGMfygioJ+8EAHBRQlL/Ji
/xWZzUvu0OPPyGNOIFEqjIKWIRYjB6KbPNVZKN81Fy/Rk0QiM2tvcT6wXQh9IlKLGZH31TSBymBG
JcMOkXhINNv5tvAN5aoe6AAKWj5CJnA7E3SHhqlASLfXY2CaCKY1gAoCNfKbO9Qny8bQ+PCa+WVk
sfFtDqQWBsVSHew3G2fz0VZ8DZ1Hv6GT8FkYLfQ1lv6FR867HNwR+QI/JrW0OFoN6kWe12zwVdkn
zzPTctoAcFZsGcE0K3HT9fKBqzbrIchMuYSrbxz0ih1vySTMLQMvd5Bb4SBkqUg1mL4XojONgE7u
wtOOrPUTUqmxJQ9CdHhAeOOs6CVh7nkOMt0/x+xZzen/tYYtr6eWrbwx+W5o2SWaQ+8tdctE/5gE
6phsmjmLDkuWlTbEbNZCKCsZeyEmmUmoThM3fLYIWTah0EejqWt7xdWhjg5oOULPLWc6Y2bkaHNu
JBKXBHmiWBBCgHJ26GgolslXhFsxQWEZqboQoL/UUgiwV+/r6QqmoeZxwNU1nTFVwr5iSh7qgR3a
uvuysVUL9RIz+rYFgMoX+mUiSrv+Zk/QkNRpbDLTciAhpuyP2k1tsPe8K07Tii1BmDwxnyw/dmX8
8ewhHz5tY261qoHOv9Fo7M1W3AVxXFwwv4i44fz0nXzTsb5Y4pzMWtYc1W/U/V3lhIxeCjBumm51
IPepTjYy+QNm0ETEZfLDglMnrUl0xW5SAt6CIG4M71J6y9kW5aAc7tzUbsR46kHOLelGfbvgEF9Z
B24Pztxuxp4zKBweaviF+dplddSG+H6QNmDej/G3sZrhy2ytkBCEjGJUZKFcNhhivd0hWgDqCvrZ
gF8aetxbazK7t3qq0NDkOQbXbkhO/PBlVkwm2vGJFM18kAjovRgxUocmTI7ET3VhmxWM+3lnc4Bv
XkLOaZ3WokNX8sqjYI1Czj75wqPuuFxekKhAA2l5HVG19byO7ivoTYLOKOb4PYAa2AGUuMv4cdh0
v2So7IJJlpOAGgsYu6Z7QVIXXsLKthO1jTTFA3Ss85/lZ/I2kZGxK+dlxvguNtoxuCHyo7KV7BvS
2WsGHoQOhQ6hMTbTD+aFbNizJpgoza1Z+ly16lBhaKCBVeDmR2Wfq4Zaom7Uuqqp4lE6Zk/6QoY2
wsCWmBT9s1fTv5OUYJDUIFz8kKuqkhnExkf803qDCiRhB7k5EifRJiqvyrrZdL9Fa8w7tK0YGI81
2DxRq7EyQ3ATAjhFX7TfsGebpSTb4Nu9j2IWhWuQFYkpgyIithAiZd2SKGkz28jxLXRNLBRcSvBC
Uild3XivT/IJ3SOnNKBBgfv63p6MpiLQ5wz4GSaRFsIw0V2EACZH15fSOoWleljBP1mlofJGZ0jV
EZuqiZUwILZKSQO3Lz2ih+UzR1Gow3FPeN6Ynqpx+bSHL8GpLp+7Fg8KrMxmKO3eBr/TOYAEBl1V
/T0jQf2BN15XDqf0OgUmwWrNpkRzSl3yNjr1BjHaHWfZdiIevoCqs1v7fY1+o0m7Owrk3sRhbXAb
8HyjvIoARhIk7tHHP8wKpUTSmZgjVz3xGOwl0H5d4ZiI+QldSWABF1d3YLERqKR8XM4jvcLxKcZh
BTTembQGB9l4a1x91n0IBsXVHQvDfEYypXwIjsqU9dl3tqUdB6+dhwGGmfAdsMcjoVZ+rjKwhRI6
A1PIPlkMWxndHIXWsfjorq4KvIjqEY7FRBCoMj5D3PFHTO+SaaKs7aR3url2MCLPyepUj7LWM7c0
4t9ceDb8kT0f8l6GYJiaH+sTJLmh7xG+YMQQKnivDxXcglIURzHjSVIoOTxAo8Tt+nR023JHoGAW
0Ijow8QgdG1FnzpBfbN6vvNVfatc2+k8YPmqwznYGB5ocvPB0BoePeKFDlsXstpv9jIBDmwlePgh
UFnO9IdNVT5gWX6YJg49yiwcSxW0Mv0z3XaMzxBiQwr09Fjq42vVIXQpFDzXKGz2OeHUUK7/dbgz
kd+2sBBT8gUwmwCr5vS9KDLyBE5HEJwXwwcnJ5OoLQU5SUFuNlSbPpU4O5Kbc6ubn2zY4OrnNBia
Ifb9uymZXYqrpJppJtyHh7B1+b9M2+zs+3jzvbY1gBPjZjMzjWwZh02GkLaQnPUHhOR2LKys9Qe7
eLlY/bcFo19jOezXfI/uunxeCoQyqDPeno3yopNxiYuzxRvmZkTd6a5hz+LeRklSIpU+nJhIUkLJ
XKL0CmLaj1c0anNA6/ARMrUk2Isj2q76PvnSVpcIKlRKWsfbp/1wdhe6PPbLr22adaPm551eEcgL
pXfH5k/eXxxvnO6R/mkTxrL5m23sIqnUv9lOtzhjt1u8rdSWne8W1KGEnGcZdiROnz//57NaXEY7
IdwIf1YYHdWFFzRdhxo8wHnrxI539JPTfE5lvq+mEemPgZyi3ZhEqneWLN3DAOjVrDhc0wqvCcDU
wFhQejNv8xsonAyzh2U5A9vZMBYzyUVuAkQPzXLAYTLRyuGBQOfhrWDzkgac6OF07tTZpGbLoCZS
PbZefH/9Ynny0c0EYjZKwMY1czOBdO+y713CCmvZ0Gw9B2Pg2RDrzjdlq72J2ZDWyhrHH8RCKW+7
l5hZaAplqOjC2/2CJiYYbGLPWhKLaCrKuENebx47dgLauEpxPRAZAtOhYUu1HmLu73n+PZsU81PJ
RT89s/FHbD1IIriEGPp9cGZCIEYx2exRYj8TKhGyxtdgio/Fkd0+XJJcdIwjZ/YvKOE8Pnz+Nzp3
rSvJfgiYdPbFNX+OD2dVQVHrCXR1ejBJnOWFNDJM7OVndUPIphtdYUzi4miTeBIBV/FNnUCjQCMX
5RgZxgWUzQP/6TB9GFs6pfzhyjWkZp+VPPuPii7FkgO7ESlE5vwoJj8faA95N5jj/2Cov3HEhx0B
uabycGwYFbBrc/VeI/JPcAlce1hz8jgjor0hkT3hPaz6IFScA1gAmM6EDNAlAtvJDZmKoDXUdDww
8yCyeh6G6LA2m/1sqy0yGsj54Yz8/kNgKTs5361N5l0O6+SSTMpbP859Pzjut60Irzma4NTHlV6T
EkBSW7B4rPR1BnyhVjDbzcf2DMfJ4r1hUHeJ353aWCtyjf+Mj4tVWBtFXZJstCwvbNllQ+gRFS7e
DxSSLBRLeG2BoYWP+FSm4QAVfwKqvk48qcHO+zLUccZ7/bDLyWyq8bwMjyYYIRk+FekC+Id1VndO
WUMWOLS3cCboe8rnC8zienb0/ezLP9rNhqHWtRjqC3DGygVnfQwldyhyhckK9LBPYxqjamNLEyBV
35rg5lqkM2QXFsj/r45bIWT5tR0Hl3HLXTu3WbaC+NX3E9csow27OlBptYdNtjKMz9iq+IOsNkUk
GIqMPtEjl3tJerwX61tTx+ejoiPjhRKx87aWf9bKP9dgNQ69XSUh5avJ/d3Ef9Ah//v7OkmFIb/O
ObSMWlZoMVl55mgn+hwebccek5v/k1GaLyF8wxgTBN9waVMX8a/Aj6jxir5rZ4Ena0d1Y30F3wix
Fn+ManBovyQR/1ENduHc+IPiM66BizaFtEdNEc+LQh75GD6aHMNbpnyejRPvLquCSAGEP3ggr8Vo
IoG4j2pN0PuKYoTq6c/Zacs/qLUUnPL0b3MioayKH+I+U0ItDgJ/BAz6GorMyynLx0qbNZ2R0J2f
FoILN3MtyvxdcxvbcK/Q+S081n2oQSu7L1oP2ts03HGCK5P+Iu/3/rgoHuwsRfb0uOVmygMT6Rte
IE75LjKMBnDKytJvAQGYbFY3Hd5VUGAlAKdRDY4pR4LYsSw4OxRc3Cj+80CT64FP/UoowwkGMBtd
cyBSbNCuPE68ixbPLT85iN8dcgmNX0tDo4kj6GRt8J0z6H5GhF2F5xjzd1HYrmuOjR5HUsYPR0x4
lpyOk2pm2ahenfUEkVYZ+9/eqmDVfFwTLBcwcJBWipulrTLeOVDcT3yqPYZhmM9xwWh5jrQHxj41
Kxgq0hllumGIy8lFOpqT2DdZIJ3UNPZp1qrHSDZoh7Cuhg+tR710yAoBxQHlz2n+sZboJUJTOtj6
1yfSnW74V8gXsd/shIdKUrf3Y5unfHSl2T9HSf1ReyJtDS/yps2oS8YT+EmgBLKCOpy2ZCEDo0AQ
TjtFV9qfYsXaQQU2F4F65s5r6kL6TvzKjDiVPOZsrJ9ymQnD/qKSArOhs/2v+bSWqgOMupnSXiTl
R+XFz0yJWRSeH9wEkS83F/22VO2Aq/f55gkSugnFnCXYDjYagvm9eFVPOZ5zO+e+7K0JePHpRR43
PSgJJFoFOxZ7fVLR+44nw5ohCtQ/sT/wAvPogvr1zDkgdrYK3nMTk3AoEMfnMOibb5WC3qJpu0WL
0s4DdpXZhj/PIGy2P8L2O8nUdFc0LkAMINmr6A6XJXvfEW0OBDib8dPp07egbqwG6VKNr9zOHSXy
lrdhfe3hzQeZwdt1aor1UyUyk/q/8uXnE6CxF5e/m/zSQqIQnO+oNcixFO2KF+lHn+i+WSUfa1d5
rC7HMXGOEp+6I03wd+/5g54J5TpBdaHWnq/pFR+Y4llixFrUauWkp1OR8diPLK6Zz0kpHi0MQ/1Z
W+kfdJgWCgl4vkRVxtF+d35Cx/OvWc4G3YbS9FZ2n8BFzHFOyuySRIviMncZijwTL/NCMYFYaBRG
tES4/LNlaBUP67+nDtOsuseAPxWKDd1AjQWp4Pko9Z4xMCvRwfjdO74vLWmWQBLQQhErlYB8HoqY
1BVZh++q3s8JYQO7Vy8iCk165inrK4gjymO9TaXHenmVGW0JId2NbcxC5y4/+jFFqHUGPrrkD1hr
f1yOSzLJWdXy6DuiwhiVtbpZxMTQDIodZnYbZa0fz2w2Hc1hmOKUjdXdFFjGzZUidRirAK1odvud
Dpn1plVa6RA2ZPZB94PsYb/6Ccr/6xgE1xuN6/c0xUfYcF7nM/1DenLjxdFEB6riubEXHWvCKuSq
kUBi9jniXKbJpmTBYTLd7+HOKge1zsRSF0khLNFYV3cTDtu36HJ251FMW8qXX1frC1nMEAniptVI
KYCCZF0PLg5T9xtRmtoicrvzNveoM1/24kBnaP27gMWLgI2POGpeq4Iwdn93g1zX+PNQk9J9/MKa
u1a7CAD24gd/un3VA5Eh0Zi4pcmfjmdobGaXrQXvOejJuo2QcvbveQgIQUeVlv9k+FsBLr2Zd2Zh
LszE8ApbK+gj3T1Koc1FBkcgX+VUJp0uk1/iDGGoiJwQh5jYAX+i5/w/Gmq5YL2uW3V1PITQiOcM
WCg3TR/QjSj4VGpnU57oSiMKeauclwsy17S2CN++NtPMpelBop9D5pZNvlQ69QW+HsD2W+So5pN2
vlrn+/fKPJFhiJH1q/5TCG5uwSs5AjjfIFT3T74sI4b6UGC/hxdU2OxcbRpTo2cjwmoG4dCy7mcG
0/b9cAryJ8kHLdqQT3Kf1wfBBRj0nKh83Six/Mwl+Szb3qF+EEH9xd8HbDx6PQedfm1CEvkqfzYi
w6zC0JS8Ez5yQ5+/DmOuKW8nm904TsUYsW71ATCG4RLWDmnsYqa/KCC3UpGfa9ALl/tvjleoXKyk
ZPH+wj9ixsODYIZoyHicrDrKroBIZhG38CdqNLEVDZQvCsAxnoZ4w4x5fFT7ueY3Q+JlUB3tDXQU
qz0gVYhNFpT5BGVDs9GOAI5L8svUNenFERvnpTe2CGFjuaieAFCPZNBRWhkSR7VqLmAjPQQ8ULUz
pk7sKI/ZwpJHrnxOQXcErAED45EJRkxvAKCY6gdYXwxOirQbSdQRYcK7rPeKlsz56FU/cc4uTkuv
gPF+Jvuk/3v9mT7P30eKLZfQVefxFT5dYGfPSBroCdHQMsr9q23FvQBlJ82ufFumo8IHXutBr5zw
QdbSlc6EhY72HVoCKJCWF4seVE8P3zlB0hpq5OzuVg5NdMrv6cnO+33h5h+IZKwsa190RFoirpJZ
PuRXbKGUgXQXVxCt8TO5r94bold+IWxjCxYKs5+ia08IohtfwuHDe7kv3+KD6EtGf2eWUXO95cxc
UVU5QI+8Tp6Ek4j8dCDD2wsEoG6NvVhYQUL2Di5bxnbTn+ud2tWOxiHT1w8n1NFtVcOwkM00Bpau
x9XDf0OTn6gA2uk/35f44jkbrAeormiYaBwlYfOFTSvNqW0sFsC3RuNu2tod+yiiooR6eNaMCdHd
jy2HXZEBqx0Q7PxfeX4Y3RCTtaR0DFA6XdVbMM/IGaqfmS7lrfayMiKlqtvBKDby+Sslyz01MEnm
a6xcGWkne2RP2x8IHuLdTtolYyCg3ouUiHwjU/Mb/GXHnFF/UXBV93ChwJa0bazX876vPo8Eg4XU
6GLQGnAqpwHmQC/JdRoxVhhcVxyPsQvUTmSOqkiSHJOXHfiZVKpWufOtu6yLV4hr7SWSKvNHw3s6
KAARWb5tt1tCC2STve0A9ne0Posj2f+0j1uJ1evIf9GGlAxDe5zdfgnYqNEmNb/zQUW+h//megin
nadYCdgZXs/v7QshLX5jIgvwr8fPhCXKikBzA9aX3nk4M6ZlkPAAH5xbpkHXOD8L/szi1MI9XSBI
EnptR649aO/ZB8Uyt3fJpFgm5tsEx7VKBMt7bc/MUjI3ICp3VxjhHGI617WX/3X6cK127dvV8KaI
9cHXzJ356tlXM9uw3rsd4vlbeHAbuKFsaf0VcjFRPK8OQMHCeep5P28t4qoN3Z+NIDRXQcaAwvXh
6x10ouSO2aefgbx16ePS3Cw7Bqhp07eYdkWigxlzejNgjBz5WYsHYtDrtHj3RberlxaVqDm/5N8t
t7uJWMOKDvZKAhx3vFeR391yOA0CxvbufArcq8RQS0liN1sKkJ5e3JBv9QSALHRaXNgZv9Blzhlj
hG7yxJ9mfqMSVdBmc/TLKkO+114a0/TwdTllG9+ApLLGwwbG6iiEispJ3SD32VjOWmPgSAqm2IZ4
vISbGSG6wqEQ7+Q6/Klrol524CGElvovI6s0uVD1X9P/852RVD7+4J38Vo46GCHadQyFC77EYex/
rkeiS/D8NJVhMjF8gC294YPUKNWp7Vr1cEZfeOPoCIviWqAKqBdmOOlX7xv8/tKmIhB1Vpl1dxk8
e7+XS/4UK0OgC3ppxKGvvpYRVL6kGI8078ugPOMbGYH5idygE66vX87nGPgDT9u2UBEO6DlyfzFU
9AgOMBQcw75/4PPKSpaFkfdjJuFgqs2V+r6RA3L56CRnH7DXfsJev905DmhCh/eXYqbbCmmv8GxD
NBJl8ziSPIyic7Y8rgO6OtQZSXP2iYOIUWpJUcktNbr9c6/IzipmM27kax9xWyMBQPJ1XKUxMXHP
y6sR9S/TT/mfQ4DLpGx8LTER4qymNQQkhxjV6LobDpFRKK5cs2TnSB8d9Bx8XRuA5+9PhMfrev6r
ecBjQArnhX/S5z7awS5dSTCokrekFrk0Emyvn/ZtpUkjAofAnkyndzZyBn9UtPallcDM6T19qq8T
DpjUusb0HiDO0rAGgDFJf8PUV+lF+k6qlybBqbGSTMqZ7Cmhttgf/Ez3Wsu9IDP6xLoRagPAOs+p
2aTM2PwfibU5EFIKlgmvgGAO9B1+r7pXeNRecoZhjeoxGN811f8An/L5xAjtXiZl7yVIoNT9G3Vg
pPu5X0/fKQIBpdXc+InqNX2Uhh9SwiBs3R1tCxun96vVsk2C4RePGfs1N4BjxjxvXi5yWWnRI4+0
2QGnyrRgRKmdoFozt87b8YVBqXi3SBfCBB/qORztbUZlZg3bhkNxy13OQjawG4x5ecMoYCcQmukD
/WEjHpIQ4CpyMjd7gurAp7vCINBJ7oUSYsB3Ky/SD88Yzcale8lvhszvCSRBgXXELXzzyjxGF7Xr
9OtgtZOHGveiHw3Khbg3eIYjR31kPE+9apCui/OpYJf9nhgp5WTMIeGLM3MmbyW3Y6O3kZltrC1M
H9Ys29bvKf0eWJENNblRWPRB3d0w1+Hf2pvckCNVN/98Ekc9dQU6e1nwpHHUbl/1HBfc0BIJa0lw
8NT3ab7gJk6u8LPgdSN325svsK8paETpwqLwlkEgtSPNOu+dsY3nlHBSocfIUwx4m2QENLoYKlgZ
0QqWpvB22WPHogOBIEHdVSEuEkwCKjdlO1Y+FyB6URyACGEtP7ILWgz/Y9dKKvihqXfAdAnzm0er
oGrCXKXcqfsHs1Gu68fLkWHryEhgM+Zo2tD+dUZjOJZORn0sKn/ufS8nXs2n8bLkMG/8yyIdaZn3
PkkeGbG/TVhi6LLHalEZ6WBUXg5lHpv4pdOmnDbuzJuW/qGYzp2g+UZnVKkYrcc6VKtMpm+YiPJi
Jpdv9waPO9KrHS/6DGJDE6FxppVwcyFeesOuQfhHAl6N254jWZNDY6Ba7y+9CujdlEYkMC7ukTVX
4ZGKKfH44D5/mN0yGY5D9W67n03mvqNF7wMTjvIoAPXp07vcqVrFpQk0ITl/pe8rKs84g3h+sdo3
zbeqjnIJ9oxXFAg1GhF6j9aZBriU0xEG+eUXfjcj9rBKG23mpWSU3EvbcfvIiMWFZtyim7b8vfsT
2HoyeC2+fpjvx7v2Hsynwv+aql1I9wbTlEM8Ij6WS+zoTPHX+MDBtJ6ar9wrCMlj+r3eNrkZIwFt
EgXFaGWLZBQoveyESRud9jiDUTAbJWt5fPyIPsWtbp9ZlHs6mfbBrcyap/4J8iL0MYjH+z41r2DN
izLlP7L7fr1jx+rsyoRafLNw43JYRE3gThbTk54gfLXR63/UUTIiQ4lXwr5KXiJbQzRJ5VwBt64J
J5yXJ/60DEWPHqD53rVvJ7hl/gOs+NkaSP9oh5vHEj3jSDYYU+lSIiwgNTqoZPU4C8MJxsmRLRhT
3WEidTnYzgoKXUN/tnlxmYrtCRdBRItwn4evOvshlYWHrhOEwDr5XQMvgwAQz+qEh6BtpBwn1ZmK
sYKwCa7xy7gulJM6cytJEqp9VtgxICDgvCUBl3BSPqicI8iV5oKPSz371phdWoMRsjnvw1c2QX4L
IrqQFNUpvmE8OvqdQrN33x5HvjfrDpp+mSmaRKgebe+TgKsulH0FYaCaefXHkd9tVrvnGXnoojbL
qSQ6JqjLKb0AGd37w7laegOishlQYsGp/IUoH83tBpSDp6qxsdhkmZfURIwsk2czBtljKpU9Mve0
jNzxHvswXijiWtn4hfjJf61UMSDMiUGN68MJzsmnUpyKqwR6pi1Bh3fAzb/d8vgo6RlUQ6XO1u7X
tEhQTfAksaJc83IcphKfaL1ag4kSZGsle9FMU+7bjNcvSxHxvu9BZShVkaRIBTLTq51wx2/nb39A
hWNXRSbvRcsLkzc+B0BgSz/LDVDLAnd6iJSi9dH/ZKGTzMaHHkUOQyFsyveQBM6ntqtpKOMeVqKB
bb1UDWBmIepGmLraGPGQbhviztzhbdRQ5dZmZUKxDiPpFr9c4alhdS0Ct4LOB0SE+78faFeosiOg
9QokHsYEtrEbaoX3AM+WeXb/TuYSs/MD9eRrAMa5MwApqp4qs83HAnKfYimgAcxJ3nOhlSG3fOE8
Ve+ZBB2C5tvYCS9LlsPu3W/4DyiVTTS5irZj+zP36SEOZTGP04i2xqzkm3lpM6FL70Hlrt0YZL+l
L2WCh3YsJkRtIOnjU8t3bzNmAijJ/0fpVAlL69v+xfrb0wvRSJfFvAvgIAXAQ6nDR1SRkuEgVbPN
67w2QzJem24n4gdt+0J8YFqx8w5Z0TXaVkNw3Ex7jNIzqBDk+OERGZ414jRXFxqyhHEvva47YuA2
UtuagyP0Wqrwe0OSl5M6fsNDm3WN/Tp44UkZ8r01yS5RstRRe5lL0M9pkCbqDBh8h71VvtcaZx/u
FVwQxIv7mLXuxDW+BxbAWkOSLqQdJM9PF3QXc57jx6hqMIaeJm+hkXzGGEALtKkiMi7HQq851y5T
StahGsaEPymWJTLmHrAxQZBctqcP8iEKTv4oi3YeciqPsDr+DvxHRIjsMlRnrL/jQF2TioVC/fcL
YCTvMNslM9M3YL9GmKdNw/CsYhtW/ryLzYNiwatVmFEtsR1ee2sDYmRCoyHheFvnD/DNQptA+4Bw
rSgPrXbd1peUzKZHYanYXKTCkRyZZsBseBOpIUCzA0MldkGrd8BDDh/ZPLYHasxNy2EwFfm9YYsk
7a53RrwJ2ORWjw5XW2hfGdJEiETy3IAGm5acvnC43VhMTJWsSXJVuwI/mJcORiPlpIvntppZjFkg
+urk4FBhasjEhmU3ImY1wWXO3JJ9ItjkHad3X4GSyFD5JT4XrNo61IZy1JlILjhTh78CPq1gkp4c
qLfdilWrP8SLxIZ7Hq6yBXWl/JcoeeJE1UyZVFFPe5h1amR1GHKvFA7YWkVuyKE1IYgcoT0WWJqW
qwEO9OAUv/NX6l6r2aZuEokE52n+5sr5nm6camlt6N/sI9XpkJeXC1L4PNgptZ9eUTHVfckDfWgS
BemQRtkrKG3wBfv+gd4aQXjg/9GfgX/DyGgCB8MXNRjuxHmNpAGOHlwqcvWnZYi0Uk9bIOOFCCi5
EPzN9IfeoCQBJ+SV1alIr0smlg49zz6TA2PF+KQK74AhIcnK4K75kaYlCqKHqfTdpjM6S2za56gd
qTHGj60C/Q7D9XMCcm51aN4VOD24I9WvuXay8ID3vt3aHisjBIOoLOCXFucIvRM6xeEBA7ZJHjCm
TDYcnDZYl8AFofO/htDupjabenY4iVxTklSfT0D2bhxJQCfHNxpp04miy89Apr7JiDuTluxbm1X1
ova3Lcty8WVawb5MN/zjlSTnpTSov9wJpLMVVPq1Mht+aNzOvvcgrpVyA9lOqs+5NRB8aLpNJlrA
T8itk+XtfyTE3xdFFNaU/6gBbi02atzPtlxAcHeRHYKq2Oow04REYCEx62UAOPcuA2BY0qscPHRZ
5m7Q7a5gP5JlGypql8+1OWhv0YaHfupMFOfNpGNm2kzLMxQgr+T3qOlQG3MdYfb3BqUKfEdqO2Ck
VCa+GWjC0L7SBl2jFCJjDgkU7BXrfeH7IaU35MHwiPLx1XX+szT4jZwxWjgjAl1BGBUsrTNYRZDN
7hgaXJNRWfMmP6CikhoI610d6hohVbYxjcNrLjtVkrf94Oty5/fTeDOGqyAmmvwAx/qd8UGcS91d
iS/40hqaGMzvYr5REZTXtUs1jd2lB1MOVs+RLjtw0ooL+YLVpM54uUDB8jxlFtbqU6AgbTYIrOaT
OFScOnNQ/1lnsDqJK3yZUIT0M9AVyxaz74YTAoRLEv7Xov95tuAnhKwQuQS/6JiMZRnWug0BYtsJ
zh1SLzns5F2Fp2j8xhkBnGL5GQj+/eSY9uLEN+8BDKIWMSWxs9hB2Leilnud8j5MKHZdMxQzcdTv
KPSxa/2ruWamz5Z9txvzsEZGDc4nSVXYrvrdTJiO0R+9qFrS8y4qjwysob4jHxKDJ3Cogu0204nt
leMA6RDmsoToZDmRn1b1IpsgCKXXSd4okIE33r5GsmAgVe8h8hzDX/FUbXonDB24KYLRtSOp9emA
amIpe6y/NQG6dZ+vsp4bGVIn9BL9K/O3DEUg45AfJ0nae7z7pXYkH9xkgHxGOQjWlAaFVniYrD7w
ZRyJi+LHeMBGKoN/8RPqmNyzrA4I6lHMbs5HmOFFDVYKbVzTu7MDUwfT07FOtKa1XO2iBPqOFXws
UvVWYZBOctX0IF0NoXY21A/6IW1hC6emhg6dL0Sc35M+dyxbJMQwY0u9b48Klji+ew9aurNK6V+3
OO1kyqmjK1jNgt4NXBxOWWLdC2WCUasYyBJ6ECPkWAzElSF33QPT717I1j/oY2WaTc2EPtWG1gaf
o9KZ9GeucMvWC7NbCGu5uzK0Y/nFWuMTlyJGaBDLIiBxaBK8B9PW2bv9S05xhj+WxAzuSIjS3AaP
Q0Tnl+3ui2k8iPFv8EBztdsCAbmxyv2rQa8Og1w3yBE1xPk9seTRiFsbKaucdDZmTsxEKEi7DxY9
7ZwL4uCM4xDUYnWr8QiQ0xyFoGmwk9rGRH9WOB8P6FSAV9vg1mtm95RXERkXFIHIjroBScm1KsRo
jaU9s5YrEjedl+JhQl0kG45W33KR4kexgvj9IlV0Pn0fhrQ6CMEMZQ0wynBYNf2KBgeuDhqmJXud
4e8/9PHXJOkHecPwCKfVwvMeXAfWgbx6suUwqpWezYBJ5OiODBwVYhZUpYm6KncvitZMlrpByGb9
E+3VQhKGQ8CNn48fWEZScWxVf5LVZN+mhBRZ2zkvkuQpaQ0TeI2vEmUmQ9FROeMcmjbRSMvtyLoA
az4Hy43/fBAXUB+hsXjfkZ5RrtrnLP2pD9FYUTM/ZvQawjxMcV9U5x8GjvVlhhzhg4Wdlon29UhT
f6dpP7/zXJmaGzFR3qAOKlZ9DcfToaAoTgVeV2boviB9B0bvqYhFUAttklXTbszjeHPbCMdlDBDt
P2UzW5JM5eOmeaZelgZouuHCYGQ27a9xga5lWhkOzwQnFC5kgZs3VFprK6EyH0SKLs5Ohni4Q0m3
8x67LaF6Oo7t/4aO7ihxtMLfQ32SyD0U8k20QDjxn6ZYch2+RbxfOHeI5/ah+Zh9KOHLdfwKo+tH
ob69plYh7Rt1TGvN+Mt613fAJ+K284rNNrewonPIFOvv3JowLXQVvOyCJIeetb55VFwvtSUOgI80
D2ymOz8n/ncWA9NDfZhQm28XPJcw1L2IZ8PuTiUu4BtHd5l9/QCF/ecrhiHXKHfpkQIc4DO6prf/
4XyzsI9NeWHl3RRHqLDe6/AfNHQOExVaoAxCGpSOA5tykR+1s2ok2u2z0faqaWObeJ9ctXrK0xkW
+KmvvzAngYSlXW5dPgWg/yXdoFfrQnZHqdKaowlGmbIR1VnUkjxvEWLkxTt+dM7p1MJbJdQtnG/9
HWXZSfSH5kge/9NJJBV4SZKhZ2LrrtkgEOBIKuijrSWbuIjdSJNDrBTAucy43v2pGS0Nlk+ZlEMi
CTtXX5kb0Lq7W7IK+lR7AJZC/F/uV8F11iPexavPD6m9qU0Mrq2stfR5gb+KVaIooixM+EOQbUF7
VQdwLxfvca/rtRQxHnl2ByXO89cBTsuMYiTWUMH7GiqSTguSEKDSjTx4/lKcEInkpxYLOv7CbDin
V5ZtvivqtuqtE6yD+acPCwlVihFAQ6x72unE1MQksdx52VDJwzED5K1IoDva5HZgpdcuuLynj4bL
bIa3DZFkgck2Ol6PPIkfFwz1U7l7d8JDO8jd+cobqOtQyV4Ky9nbneH71TsmF2de2Agr/cIrsT5b
ReM8L33OSq+1Owoy+ASZelNjt8FXot+hoG5E/xH/qSu3iCcYuMYy9uqgiuMh5BBphyEyEaUC9eVO
IwmhMquvOPG2xOxkMqtgEFO3iw9EeJWOxQr7IgFfFjuNj7LDc6Ff90AA71WLiyMxuY3ehZzK0Jbu
SSJeNiCWxgii1BTXn/dcnt8lM8gYIJMI4jnfUmx+lXE/k21vYY3if3jmx6JbgjGvKwnCXwy7qdvL
JhFqlQzJyc4qw5ua0LyF1f2NVRqrRju/SiWAUWDUCwx/kZucYPmTEjMqFcpVurBkDzuMzn67kUT6
yKc5TSKwna/4wwHL1ro/64g/LpXbcRHKMwQ2l1OXtn/tQuiJ9f31SO/31zMKXGjxaAXzw0uNA63Q
9brrltmywApHbnZSOwa0W5Ncx1pFP0474TrMQTMfaPQej+c6z1x3ufJvryvRylSkNqY3OCt0FzOj
5Cp2m/0por/Ie52F3vzNFSvFXIeQsz1OjXEEn6SBw8pQCNuhO37Ua/YSIDQhZ9Bncy8LB5x/TGdH
4DUzwzTE/nMhmv1iikITo39ht+a/nPApeRggrrZ3ejvb06jI1YOgOEw9vHZ2tHEioecaDNQeul1X
qS05bGkCPF5lXGLYdBgX3vO/3S3srmjsbpGyuXw1DXW6DVkjr0YKcA095bdoIebPXqr9O9mf29J1
dlsgGc2FHV65SfLyFSyzJageVnojqmkMX7b6coZVLyhRXfXpGGOq28USKIV2WWmWTSDupF2/FMQS
cDyxZIEbxVZ2i5pTijt2KPTEjljSni2JLjI6fCu6Oo738L/gO6JBdX7rqfoMj/UNidThJtDC0GUu
4YSRS5ENgFh+ff3XFvrzFuR9jB/y+PeOIlceGnS2TVBAOiIfdMPHqIXHfXKyt7wXWcjUOqDmj4Vz
TmRFj4q5ajjZH3sO1gdPCZg8RumzuBo+4dKgXfSW9OOG5iaq65qkWH1rkNBtBJuJujy7Qaw4wcal
mCmZ75KsYVlzNx8JnBmz8PcsVcnPwu3obF67OMDFcxCbfPCIlXtyQCls/swdOI7guME/qvUg1sTe
QfLKtkrWl/iOCt+OJ2eWO4er3GRNTGC1Vo3OV8GJOl96wy/UZYFyJJc9XZ+2BqvN8rqfZAax5E0s
Q6tx49VjRG7igxnYVgt6Uo5EckyOIdSRjtsH516qDOs8Wi4ANuVmHIEQo3MqvneKMWkDqLSkY/3P
Hjgb3KNOEfjUWR9IyPDMBe38upnpDUJYjPjsJlTtDRvo9X9LEdjzLTFB8/PBQvRC03QkkffWaUul
J85A/6j+lh6zI5EasNUWIzR+x5KL6Mn6qT0aLG3be3sdhWyKE7Lo2tj7ZIzQRHomF3GiGIvjOKv/
B4BkWznxidRo+W9cSMwy7kwWei2MT4SrauUH4fP2NzyU7li/2P9qH4O01+4SqCwIaq00mLehM3wf
z1xKkVZVXKs9QN+jSdTXvQm+VK6o0ypbRR5qDzafeiQDQwseQJX/G4oog88o6IArMwdVMoTckHk3
BN493vAZlMy+qSPeFLDQ21R9vyiUaXV/OFxiWpGY/U+A7IrQH6ehyHzOWMJgreHf4L4Vzgz4jWKw
2iSI4ecLncM8U1crsfC3TMK6OvAZuPAyHh9f6brDJiLHJnn8Fu+3QmJO6GL85NddkgyOjNhQvCaV
CbPl6PJX9SOeKl++6Sy/QqEuhwXyt7q2t00fm6caedsKoT+zx0N368mcXtiSF1NKLsBPLr4R5vfQ
gNcgiR4AcaitSTNaMgACXBKjHqRWWoVYaJtL1oyRQL5qvVg3zoX/JefaJ+Z1ZwuqyYf6T6qhqBDa
vHr29PkcmVnD+f7RIVwuYp5YnWJLu5lEvFOhpVM0fFjYYG5ykz7iWCe0qNyFTjvLgLWV0WvlOzcz
KAm0TZ50FftUOS5glOEUYBoEqKsaaPxcSP7OzPCRRIvveVbeiARQgBpfKYZ49oVfU/ftkX6of/6R
5U6jt87rsY/Ad1mBm5xxsZIkPBt0sUapgUKpTs21WYUqsUeiJQ+U9MqSvKZl8qztB9rI/5a3ILPg
19kmFavTKfyHWq6u485KJMMSc+awIg30glUfNsiddBHEwayZLSVWdpT6/x4c0k+WGJf8zIe6lpz/
ojiDLMm1p7ulRb6Xhj+mVF6EZsg3N+QnXZJQHunhwhO4IryUfworLhnCl1P+N/cnqK2QtafNCT0C
Sa4dbfZ9hknVehzLmJ8VvavtovmliZ3/NoMJCxqztzZ4bVxl+pI8NHJxjuo8st4AI3GYV4MDnuDk
ucKCHFo+8XhuDpLmPYBJ8VsQT4zodI3px/wI8IwISh6YSZy8X23ACrfq/8DGoxYHwEsrCF8vUIeS
WVYzIaFFiVEFGzlYGE3Sbrx/BZZH8Efo3jfDeMyce5UXHyOF7OMVdK3O7PrCkvdPEPq+1HlPh5gr
LKmb7fZCJRaqZuY1WLsi8iykzhhoW4WXyiGYDIhmQwZAKcXGeQQuNgWWotZiTmn4pa74ZmXxqVv0
y3OY47zrKTmlDg0CRn2RyC4bBY96ZB6yRXFmECeq6GXDzqpCHeBEoAANCOinQ/jXlHpR2oXD40HH
IYQf46MEP9w29eJpFprpWATerv3NAhhiVm7JkxYfyKpl4HFCINMAu+8J8Qr1Iyy5IV66EZ1ou0rj
ewM6Jt5FYJ1nKSL5Jxsii0KGkbcvRSC186HKojAISvxhmtL5fx2PaJez76hrucS8ATh7/RuzTS2J
2Is1CZ3HQRAc9cN4lTkFJrmkA6iCGLSQ4DYVr7wXR8JUZ8zo0b/dsP6F0qF7KgrdQZNYHWRp1LPU
1QJOsZC5iNuR9ki0WASrP3I+dxDgZPQ24sjGFT5L9oOV1SyR4iGxJHZNhQQMSLUBzUNgRa6ZHb//
GbU2tAiXovh1e6/qenSqhORDlsl9wTQCaXf1z8sJ9/NR4y2st83Bh5I4iXCFlei9SHQSyCyxlXjK
0WfVF/iW4FWYnmUtt/GJ88Y49mNc1A5ajTN05yIq7ew2kNouOb/VugPxTmZdzpLRX2jOUBGbOHoE
mUkh6MBR6xNlZlpQTMTO8zNW2SUWSNb4As6cmVJ0rXkS6dML9JTzjcGiAhjiKQwi0p7ENbwCRLEU
/skoF/j82bpQCH8n3vrbXxC6aiJKB8DiTPAQneKSOe+2yvlE2F5nKA8BShTqITSRE4ozIY2QokRi
5jyAnpO5n93qejv4PHLaXmecJZLujaiJx2/wl5u5pEu7L6LN+aCKqaWslTMhzlxggO+nH0nGFwBH
DQ5S4152BQ74EXlfy/vcZf23catBU/W78i+/6gXpfkw562Azkfus/T+vNivRIhn0PgzAITY6t12v
XiK9uSWgOsGXy/9GqKfNR/SCIvZgiQPkyMARgHeQ2MIN6dOMKG6npVAc38jqoefc5fyGh+Jx0OcU
LbbkZsHRPviXEGP48gsaWwTnSgWZBtXn/80rtAyTtdssiUBk3BiE94egluC0xoGcuCukBx+ndU5e
SQ3ZDYs0HKyt3hmeVGO5eQoKp8oDH7QzkqWstcNFZdcVo/vLGXNrtmVRgJbuzp8zHJYsLIzB33Rd
HkNbfI8RLd8/zAtrM7GFfmQRnbKGwTJpTouTuIKzIau5hY/zl1S1X7624yyY8DRC91PaPRVmtEHB
Zaoo2Uakuamq+Kbz1+hdLq8o5bSfyp6uDehty8cac0YKcVdSyxgvOOgoaKhR1T0EsbWJEaBHXJpL
BQP96vI5dXub14dJqorwuKHqBJCCMdEE69Pf35z+HAEWOtlvY83XujOAJB7L+DCqbIifBxQc+ED8
duRd/UNfe6ssseAoAbZNfYlxOP9ZhbHZ8utOeQ9UkRu/UUl1XQPfkZ4vmWpdkyZCxFuxSYhic/pF
dRKwbujmavsjfeGEM9T5jMlA2l9pjCr6TNPJjLpWA+/I633Cx1yx3Y15GKSHlMw8Vdca9d4P4GYY
aEb9XeLcRG4dhbrBEIUylLfM592t1VypSL07N5d9bw8QxbjrZoMsiKYDWQjOsdF5vA7MVgcdeORc
06Oa0KIIyJrz0ruwrulcejYEe2yz0EOKSKJZ3p0qlHRpKsUjqS/yPs4+QtpdeYQViOvNrFg+AVXO
Iez8Rwi0S42iy7sfWmKBbp/W/LT4qnAdUFmWtrMxS+Kgs5oGee/vLMNTLhfQQRahEXiwtMUB7Rnn
7rqPQb0i47Ah6F/qLLKxL4LyOl7Lieb426nmob9gwA03KEYCiKt3klkPrvUGjJUXz9/OJLISiIS2
wAt1ujzlurbH0KNlbq9+T0ocrFqmrvnnv07czLLQDdDhhlK6VeSqf/D6lVcZ22vxj+ocJQ3bJlGg
bHTuTtlDYTqq2ip3GAOgnmbrZU2qT7YQnuz3gr+MQPBlEpmefKyUbuHkEOFQtgpVD7QjZ4W4JAHr
G6Khi/46XxUrjI7Vf01wbQLQDWicgpj4Nq9OWMhYbEjlbHISCp/v5QU7PT4DhSwwfwHUnug9mEoR
nax9s9Wr79pplgfnqqcDq14sBt4HfZeam8UNE47YQG7t96cGFLxHE3vioTaOAXWlX1F3hduDR5rx
NzyO4orTYwIx74ZEBXpKO06HvgMTc6BIA6WME18WB8RObQRWPl6K2sLNJLyWe9gv/LQTIqLeuKAL
8Cc1PsqYG/rGDCH+i28YpbWntQUcE0YWlQUAGOrQ4gKdDLGpTrmIrylmyj5sybgM8XNPCn87k8Is
OQ9xEelt57OngjgDO9bvmowPDs0HRABeis82ZptFz2sVq3KRi7QSbIh6A/q7VbOGZlI33e8AuIG+
K8y3ZKV32ypS7rFNHons2qdN9IjFZHSIKyExXUGLkvFuIJMCOOKtvU7rahDhAIoI4d77vY1ONGCo
lO4WudG0zxtXGuD4Rlm+wuPapkVCotZdo2DJBm/7h/FxmcfmkZfbmLn4vWlWd28WoaD8HnbJTM1x
X/lLHnZsQRbTbaDa+ujdGfPJOCY8Tv/AbUMM/IQfvWEWYGY7+rkgMlp2SUWfzyQwTEflCGl1zf8j
4cWLW2Ysc7toCh6J/I9El5hIF67R7h2tKuzjtWZ+0eKB4/kTw9X+D4QdlXl70RXv9k+LUxVT81rM
/OFB85Zba35E9HNeAqJnPW0yssn8qqA/pNdeUTYY7pbqlUBKb9uDRFVMP32BTjtOLjhmUIlgsxqW
C8LpEo7/E09JtLOYvsgtb4NHCiHbAbq8AEPIhmcvKOgqw5QQKkGdXGklBZGyRvi5QGkDCC9D2s+D
wEugO4qWkrUnG9awsS7jtpw4zhbGYWChYhjvx1X2ONCeJZIdysqPNnMpgATnsMXmNYbHUiY/Lqja
Ra2fKjW4wR6e3XEYT3nLw1j9vkhHZRaUIZ/sIvQMcPmX35yVRF7jwnY0Ho5jUwxXwiGrX8uhO//c
EBXWL/2HUruEwCKsZkUSbm8J6WkUkTabVkmDWIaSwFejEOu0m5K3n4e7ziJKQnhnqSuXtMbl8VJr
Y4WJij8mNQYbtu10MVBRFFwWinjwqbxYJ+f7UUFXiNWdofkdIwi/Sd43WSZf6AdjJIr6g21Sbo3W
OGAwzVu06T+kI9lfSVhezkGutGJhMiaTjX44pR8ZpZ95Sd8Aa6Bc6Cc77+IKFJktvGoQZhmenAUR
n4uTgMFvvd41zRJDJDIZPgJ98pJTLkHI8eCTpGf75rvBFKAZ7wFJie5bPG7Co/MPK0mn6AT523/M
KhEp218E8YZvzZnnjqZynhTnxau5bgn3AgDFIJILcIiQWMgmxz3Ks0ZSDXbbrgUdNbaiAmjF4r2P
GkIs0YlEg0/AZfllk3CmCZ4b6xtr1xp7mxW715yySKcpx1oppxngbRNhSAO7dvf0i4wuQtazKVwS
ANt5WpHLvcIiNdYfNquZi6caT2AC0s7XokHikcEkm3IvR0xmOeJtstdrdXdme+7XVsQ3fc5aDcmx
zfdhvEs7p9Yoiz+SwY1Kon7GS+XPadrjGzxPzYgU0iDTNgZAA3kpLjROvLiRRqcM/3eZ0lyUmXvA
erGEmJ+T9yUkGWWkBIbDTDwMqAKOG0U1zNGZ52QBgtRSmO9xFfyYna+SJikZ1Zr8A0cDAoWCfZw/
z6tUTVjBN2u3OQ2gkIK+eryvFa+f3t1oL/OL7pm338KvR8FGRd6qNr8cu0E7O8mz8KftqR9L4+z8
TqnuXBsQX8bYXecIC9E0t3OIz8jq8qMjVQysTT3CV0rX+ct+CRZG5zcLrivhXFfameiKxQXaf/nK
TC/+ZLJanwok9K5uf1cty2HrJreepqFhNlv/g0bp8oRK/ZEyUsAktXa6Qu55GO8phV7VzPQwnvp8
Z2grnZHS0AmLqTMAW2KY0hwzEcN1vQCb3QULFcsQiaN42jHDvRgfia5YzDMzfHrCIeIxXlzAoTUE
nStdn9i9CMGrQaqOi4ou5zcrYqnsq9NimsvnyX1j37T5OuFcclEhlxzzzmAxVtoW1cu90kEh43L1
Eky4k0Pb6ysGVCpwOs0OKVo4YblSXGAG1hoHFY5nEtjZ4ucVebalnFqcSXQ0lueTI1LN/PABnpm4
8IUENzErYu+kLvfRhf/wBRodLGtS8mrFYduNPKmFvJK6AiReV09HVxXhAcLkVPMhZeqCUtiBcBC1
/jwIldf2ihiVaUVNb5NIMsIsqwfa25ZhCy3HPDvnUkylsIRq78unv+pBFuvotc2cqlfGcNvSdYr7
nLVQdJwGTW+ui3Anvg3CGvgbBckOii/VqcBOtTFMYW6KoYtcsaix/dhPx4drAPOj+kjJglrCnDcm
6yGBM2DlItYRZEmqL1oMGStpuu84xHkULNDAvlZ4dyZVDro9MKsrfS/N3IvnktTXfyxkAL0FGCH8
jtChyeOqsGODKPpv8RVT+fWVg+s2aywlOBPnMWfgLjBLaK3hS0X4DlaKVv+QvPspFgB9DypyZqnt
H8f1zb6uHYD9CxUkwFl1+RqiGnzUhD6qarGBo+PThlxOBwn9z6zocLr6uIkyv3QNJB6OQH4XMH+M
mDpzphBztlYM62VJXZQVuCFRCpVYlPj+vR1fSaY+8EZbcYKXk0Qvh5r4JuYYCAdvWWmEI5P8fmzA
SQrX3Hp/hvy2FydzKH4GXkLdhSuvp7Z6m56+FEdw2W/gdUE7YJWCJ9VeWGqxj5PAbP65AORx3g3c
0sESUiN4HiKAWfPSiukQpo2VsiyCsPNm2Lx5rLNYkxyGTGY3LTiP7XY5a+UGgPFQOF2tke+xjwQV
C73Zyi9ixH3ytVHmtsuILiE40C3URHOADclbrjcuJJjWARcADUJeTKCb5BpnsLj9+1/WUo8I5Pi2
rb7uBjWm8veSKWDZa49/4A+AEKyScegg05j6mPr/prK6gDtsFNL8BimlKAVVdG1ievozu8CrFPg9
0V5sNo7UzYQ2UR3QYY3y1bVb4VO4I3v0NDH7EK5CjdWMKOXSG08zrIynPDcEZDc+ZYsjav0y40RV
LK9QXtWLgtHV1wICTxn3hxTJSueyzw6plOu/jzNI4v+ONmf42O6/i9PdhaET2PxemzwCiRgcLpls
ooeVgPaHGABRHpNZ2E/obfY5rTCUrMC/BMMj6n8PKx6R6V4Swvd/rB/C6NgkbMB5ozPgQUriH7fc
W8aNEz+M8ofVZW/smGTndX9E5qgszsWRU8dAzvN9Zsw/ucRMzEOuMLcz+tLT5FtdFL5jgGJgo+9f
XKKssctYviCZwrFxSRkz7NSqDZoQxRTpipu4fdjjsGehUEAThMxe1HffPz1F8z5oWwavuri6fZbs
D4Cb/AWiEsuZB60Ub7m/Ptwu77x+nK14l1+yH2fgfP8Y6nH8ndnmnlAMX44/AEuvfeEGkR9fbbvs
/FSmW1DYN4XwkoSfY4HGAtumE4YKCwPd3EyQbrKgnnJrk6tj9fwshboVHAruEPeJhAZ4a80QLq/J
mPkx7VTF2btARJ53jHlqSwAuIWSCM3xiK/sSHR3dIkM50nOd7UWV2tMDIMWZnrYdGxGuOxcLd52P
zxW7Zqr7U4ctPoZ4T+TDkLrW3eng7PFxcaDTaibpEz7PIpRBIAGL3XK9x8VNtAKjHnBrtLD+qFd6
ZBuK/kM1eWU7jOuMQaH0380EBaA7vx7y3ncrpaR/tumWKDtarXK+mSxEM7UvKHw9pxuTdBqpYScu
7wfr7WN1fd/mnNUvPRZcMAqDY8NPNWgS+2ySktEouV4pgaqb6/THnLvN84l8edjojL5StRMi7QC5
5Lk+h+9GNZ+zGFCN5C5MiWRHgAxdwYUNgNYMMmpOM9+5fsTGcQVpHjet/T6AxEvTvIxEPi5Z7qsL
EEeMK4HQnIY1X42EQnfIc6fJyw4DLmplItck0WzpnBDXmUavZDsYoK3LcAPx/bc+6bqOz/YM4gTy
DayIHF2kZOOFY4GIg+CRj5JoFNv2nzMDA8dO591eafENya/hUIfUfjjWNOiLchoiHhAoSHjYJ944
OnsBPZ52xUvhgO5YA2KBvs2eFlgojghRpeyxOTBIgZGKX/TH/5V+r8RsIRhWEVtt08gazGTaVXKC
mVTdHfPL9OaxuTsW0beOpktti046L0wYcqwYuhOlt2DsmPlZCX7krxGC0JpKxkXiTjiLub5SNKAg
7qtvY+4SEcOhfjEeQtxmuhbeWMG9oJR+B5hxgvdogdSZQsn5NaaUWW2hNYn/dVZYW5hQegRDEH9K
RLfMaDLtGwyVsTPz6SQYy5SWVeo6k2EPTgRA3yu0+Fvn4MiR63WvFaIWPuA8AN/NJRfQ3UO9Plf+
UkZjDDMBjEgDecNC7JcIdLn0M3LKSSpYir4RMhdnWFemuoOoP4MLhGM0thzBOEFTyMi9HASithX7
jAwZLtWvfyo+ix1uXRtXaUav2lXiv8f6WSfALmVT8j1qrL/iYtibRMXRRWP9xgWsudSg+zkV+ioY
EkeItdOEZ0EB22Zz/MOMFXX1j97JLTAn09HMB5XAKNB0RVuBrZwwO8ztqBWuqpjGXcR7KXegOH4d
EtV0Jr4M3iZmbeM81VULyVZ/WdTEugoFBW/0k9bYYpCn91bSaOYNR3LcKGUccQyJ5jg82HWwHz7P
JID49+fgpa4hSHN6kO2lSJiiZyJoe/0ygUnmAaO8KsDjXh9mJr5CN0c/jJ1AzJIQ+DD+p1BvBbBz
rOn2Zy9wplqZW9vadb1hvwytwrl/qZUL+sBjXE6tgrzMm2ldtW4a1sIvVDRPeBPKikpHVXZkdnBR
fFJ53n2wlumj3FKL2N9/lMR9W2+VK9okKocH5rfZt1cv6nW9+WkX2rTYkDv4I/WQcZhg8231Edjx
ca9Dd78bb39Z8LKcXEYl6DA0v80w1HGNuftTbYzMNR8UuUZuZvLA3iIkEfEYdUzlXV0WR5C9taPz
TpYf7t8HUKfa7l3iRgx44D4fwg4Lf0P2y0AasB22hBt/AtFSXO3obut1bXiDuRCgieDs8Tvf+Ebr
wZqJEBnhCjR5Sy1zPAgtWjUdMLnKVEoGbKhi5FBpLS+qK+E4N0HmoDzd3Q2maPIQkdUD7oHXRvyy
Vras1MymNkFsToEAPmwSLf0IhlJ3bL2MzaSYU3KOuzxmQ67IjXscJQF00SxQzvDTte03mZ5E/IRQ
JDxpQz7s7pAeW0fqrBNsORWXCo1Nx5RiVwRw1rTy4Dj8pg9Pxrfnxbzw1rvYqyPHarjPnBtYE+T1
5jHbDUcSxZsS6LWIYuyKWtxQo/rHYt83g7ks2Ua4UhfekzzIuFBON9Qsld6+OwZ3720EmlHddpo2
OednHF9pIHRrksibmiGDStyXs0H7Fv8YZWrFmq/BLpxhADYYkewaPDaaWq1TI77zvt1965fKZNAj
ZZ18YW5KkbpEDGadkyrL5xjB/i4suWkMH14hzGr+vHz0BOWRcZuJQ9pZ+KZv/aht05tLd9A0WJ/L
PQXrdMtiMZLUjWKe9uYfSdCOfQYVDB6F4KUik+zBETwPPwpRWi56u/76YV1ce2LELv87lttI3nkz
eM1kgyEbtg3ZXrM+o+4C78Ml7kAX0Op/Kkdbjghm/KPvulmy0P28zRLwXDcIdicxvLgZZWNKXWGb
u5T2231vVUKgkW0yQeGbERvYiOQ3cp/6qoldBYSAhcyVWsiP6+NC0ID3yBFCsFfT0+t6r4/o8Spz
dCVS7PmjlwuQB4WZtbBKB7eoRL9mFpreFoQg3DIp/ybiojG71b7rfVcFLWmT4s679ZbfCQXw2Ub2
LWohaLX/XO/skXMFVP2JcLySKJiVERw1RvOird7Nzugx2oQMlvFYVbOWM/u6VgcoqtZgokfPoD7Q
Z78NBUZxAJ3qf8RMAJximV6G62RKKo4USh2s0wjUZ4viSG01DqrfhkhZxeIf2tZtDh62xcDw0nml
bJZ0532WlQIrg62HCQiKfGWh147SO0SMVqXyizvl+kLU5Kf6eKxRbqaFoArJJg3mUjlMHdfFacsO
Leq6tptQRFUqoohoijuDrhsnGP/bV7GJJ8/yoRfEsu3FK2uhrNpR47iG7k1l2DotpTRr3ZQnco0f
MDRRLG4rpvsh4uB/2ClQpQ+GsChGeMDQOMfV3+uW4YbQ9GwTKsBzLYV5UTwk8cmPTgjDW5mXLWEm
8IHFmi6UYjE7BEyvMV3pJBI6BsBjDol9HYu42VDQIbi6enoFTBsseArtHhI5PjA2OwqkVLEHCWwU
/eoithElck4u1o3kNYYhGMlyPIxhqxW4nvKIvVMw8K+pP2B65Wo4YkTkAxVFY9RCHVw1I9s1SI0e
T2AhF6s/bjTzQDrQ4eMqWstN15p2B6rj0G8Oy9ZexFh61LRb6gXvvhqWMiPSVjDdh5LYUf9xpv9f
ecFCKa3J8AT35djJUdGATMmlMlxjmkYWwcfTsOrAWhDxB5lXrNZP3md6KcHbUgwKcCzs4kGCwyLE
33XLeec3aZdzlzQgrm9gOz18yDcoQB0KeDaaR8jjpPwtCjwwAVuaYs4+pQkph8ToUcqbOLrCUrZP
wbLXdE/QGgYy8Km+2opqxXsL8sX0JEBK07Tk5E+2iojTk1vqA7y6Ke258Z/IzXgowFvs4KtdY/XP
rwbtViUVO2xtpVHHX7Gv6fRlck+wMflmc/wuVrLZAWNjy409KCnS0LFX37mpus/99mT2NoXzIx4y
ic9DaII7VqYbR+W/8ytqSmtoCyMMoZ2DKA5XcSCwfuFLXyHhJwF60xsC0Hb+ifq/WiP5CknJ5KT5
30VtFo28GpkYN1nZYTiQnB+IgVerixRfFpATtpZZqzJvPzWZZE7pfrQyP0bjrakOAqIGHpqiPDUP
Gkk1gKz1IEl83Io7OPKLBGZudcNyj/Y22oOWD49eeR3YHebX1NQ1wzwEF1ZTmp2v3ZDX/qe4CxTG
B6UFDBIn2ypizbeMs1CTi6US+MP92iw5QRjXRt0lpHddC9zCqsnjMYpZ4G5y3YZz1D6+tsjpE8F8
Q1ZGuQUXOEhm+SR3pVL5WyEVi9s61x/SBFS4Y3SAVO6YTaWvxzPFvY8ZCE9wHWuzetq/wN0NhUjm
XzeIQ6M980sNuSf54SFTyxyh9MOjpp2LUcbzhOoEvIb3jYwAD8ny+JwkneT5VGUaA0IuI/2zwQlh
kr1auSIK1p6oqYS26goKXt3/XGtttAxthLrk2iZ6+alz6Iw2DjHaqTZXq0KfTx5J8gqGvRD/q8OW
nUh0QrubUL+BaFDcH31bf3bp2tB4bBHRRvtJMiDOePrkJ3iVyOnlT1Bgb/hdna+K+Basedt2wIZ4
FJGkkfGU6odgP7W+iKZ3bK/C4TInYDh9vSUPPW8QNQDjvGecWjNspewH48+tHRZgWVlNiriP/VfX
SprBCOHNE6Ruek/zHAttU29j6o+e7iOc+W7WHwYYYhYX0c5BXFD/l+VE6g8hAeRyRmlgt9R5AC11
GPIDiyFp9IFu/+zJwfyFJg7dtSIK2NgDQ1HlF9ur9/p9WIFbST44jVyYyvhGLX1CvbIjHWD43B8S
wD7wGOMbEHE/382pHvCczieDFzAf9GWEvukm9v03nqApC8H2ZVcb5MyxK+ockfDFsDL0Ob4JtDvV
pZQHGbvEOyQ2NB7iTpKo7PSNxtKyCdjJPbfCFy2TWUm9dU+Fe/BKOEuSXQlAfXljHyBzMz4dVzeZ
iQDNfWtpe+plXVxayC1SMJ0afMBVEe8QRYT7weROXs13fUOgGZevJATF6HS0nXVGDMml+uKnD8ER
SiqdQkJLETMbPrgxfHL7YtVCnpq62Qj73333H5YNrEvitHLCmI1qu+qg92fOPM2FLdKqsgI3ipSa
e2sAl7jkcui12S2qCKhDXUqw404wad63GS9wAncwMkmxpCfS/R2x1p10M0Hp7IRk3DLl5Q1INxWl
iJqbvxYvUKmmgAjTEEPRHUxcaEwWt1DUmYvoYp8CFZgXcJEdD91IPlL0GuXwbVXr5pA8/ITaAgA5
LQDiHPL1s2fXVyX/ctZt2kd/9hkf12C4oa2yfFXzAxgUaLm1ggaYRMy9p+6aFgJ4BpbdRClDvfGt
YKjHp7UU82ig/1cGxqrwtNIYzzdlcHtn1u0dPnFK9931sj0noTEmndoByzEPJD203KM8WA35Fam+
VMneC0y1OymObfIVX219UuNADo3UUUAkYRFuzZAOW0NXOO9luQSaOqxFREGHAfUKdrEtQBxXdbW5
Xy7g6wOjWV8/6uFXCeoVXqa9kKwHhxLN+fhGNFiKbYo4+T3mERbANFsoakuEL7hRHoInkhK/9PX1
VJVMUN6hrgUIr/fmEP5q0ah5S/jkxUZe6jNk8a825aLGdmqWYy5r9V9IUMo6dg16KET/MJnkc/76
Eh9vp4AxqZvE5nUueEpkIhNpHP23bL+UBfX3WbWmtsrzLHpA+XkWeBgwslQMU1ox7OXaB7+QSCX8
/lEbmRXLKNWLwXfYvh5S0IcRL4GBnIK8awNTwlM4ihZMu9esMYbz8QQ2BWnnmmtI/nW2csH3X1+i
/8Eif8OF7Ar0GMC8pb52jPw65FZewzWC4fDg/I93ruVcwgsFu5znaovUcmJg+5L4u3zuVoGnt/tb
duEJ2POFi32GnxL9POQPR/DOhFqjUOIMO1FmBz4h/I4f0GDGqaRUnhUe3SqVWI3pEhYZZUwM2b4m
ERmoCGsppaMo39nn993Wj/G7WQUZG0mr0iKG1xsHKtI7s8Uus2+k0iwaUJSDCP23n14lY1u9Jmfz
QmnnVFgiPDxjXaIbBVzF8SZbadLVrycxdZ3667KN8EB6m1Fw3uo2Ub+56oGX6mPEBUyDH+yqwoRc
Vz9d+GVU8ghl5KY7hHlLlpE8NrTmEky0XLHifzezC31hR+nJ2g58mvWYKiGzB5DP5uMSzenfU2xL
IpGmOU7Pu0k0j2ByB6nanmDxsWIeFWQXEOiU2oR6b0nHNRuXdGZFLqLEGJsVDQA30l5njijM4Asj
07koaeoPWqyTj38JluM8NAWpkKgrIBOMk1RN4+Ff57hrJAVtQgBZsTbWC8jSszDyrzapFnEku8Iq
zM6bukHkm92df/W+v3wfzTQQSrNsTbxIyS+sLFfj+pc9ZAC8pyEa584bE2hGF8qroHHJusbafH5n
8uvd1+/hv3RriT8j1WTEN9PAq+36snR4JrxoU6a0QawrgFO3nFXmDhuYYbKLFyvbDYv8pX3tenfj
6ll9Cjw4b4vSqcqnu8i70joIw/uKyVOPGWGUCh/thzHFdlael7tx2WaI0dt1gd9PM4hepKu8cGdJ
m3zrYyazn6Vccjx0YHnk9jYkSdHqKAqJGmnYB/Zs+QZQEdYBIAjC6MhCR6c9usBRgx6mfr7fMdqO
5KD/kaQlOz9PDRA5YY+liZRu7dB0pxC1o94tXQbIk+6R5WfWESEg82P2mch/l3q9ccTjSiKEgHop
wVS70GxDl/TRHltbO83Afdo1tj/cGgvPv3PR1ewn0MrxejlARU1+ZPbG2RDZVzndzgUWyQ6cino7
VHBXKHjAH7Q3p5yESyZyuDfK0Zg+nCexsCc4AMDFHj+mep5a36HQg09JsoZNhWPPngZ+Z4ny4dTc
8TO7e26dLLeGxEM79a+sY9yocMxEtYeEfLCkt/4DE2NcAgLuFC4eSrbaJfiT9jBk32eTR4mNL7MF
Nkz88glOOpElRIjTmb2+NrQj0ShJJT7EGxECRFeMKSjREP5GYR9u93z2xJfqRXGVk2tJhp1MAre9
19jrGxvkIe706jaC7WYdXyaPyhSWpePIrDp3pO44Z4EHNvRd+AgohYp+KPLN+Yid+vOTGf9FR9qE
5Kg1MrtyfLU32c2zqpNpIuH+Rw7MVxCv6Z/ocRqaxTTk0DZ/iAU9ZItiCLTqcuztvncRQwgyoxFg
I0m8l/X4RnhyxoFWzK93wMy5g+DCQc9uviMAMhRFedUBbs1AkveqR9JhbVnnFBOCe60e+o+J8QQm
qG9aHMQN8xDWSOS3rWWZsHv7EKOkkdD/gRgDMWaNmrb7XIfdvx4/h+ILzuflkZmHpOM4470SqeLL
ekVrj8sGUFPXWtR4W+S/cDLaOLAASh6HO1VQYO9o0MBAMp5BeUj7EvlgdPGW8vVZO+TL53NxFkc9
NIjPe0/ympe7thiGKVszvOSZb7L1lIQTebPQT2iQ64yoxd49H68zettvcSTPt7L44pv/V5no9qAI
rqXTotdcHf0evJbLaGU3Pr/rxYlc8b4W9gwi1Kb5g29DCapYVy5oyla+iKhjayeT5tjOPzu8qR9Y
aPfjBE97azuxIcZvpt5AJBMXiSNdmHegB9ZCO0lu6AH5Q52U8PwhAw8R8rGGL1QexU5ZsTy6FaQc
hVvmJRBz3Ijx8TAnNIpErGdP0oBn95JUPR++Rez93KNrMcvlUQTianGY3roASMWSFUQx7SaBmsNf
Cf+T6kBlC4NMFcJMcizl5axhGlcV9eJSKEsAmM/HqwsyWaMffZyMTi07x65g+mDS9ZB6fNk7ktie
cO5tDqdVeIqrrkde779XfF8lE6pEbbhR3793U+7ovsAGkck1U8qDpV5WWS2Y/p5fQ1UK9Pq7PO+4
z8qWbgowsWisM36l9O+sHkZXMa54mKol9dEWJiuGDiIl49TCSKrOJx8ickRq2NxVwxof7fnwEt/I
IH/nDpEDQHfxkrEzWGpS6CA89lGR00Ge6hlCcqzN4fOI8XgUuWvogFRohVoGk1xI+u30YL/VaVts
dqRFR5rwxkIAcpHpj4HRO6fzLR4VsJcpyLaiuyUaEI1dwJRQuURHtVyE8DpD3pI0mDk+84nY9D7R
LM/puJWv477X5VFJvuFXvlwwgoGWMBTQMHB4vnN9kvUTvc+9OY5Or5dRi+HLYmKXncKICs0Xg6+P
X0qAKzOQ5cDdkUY7W7S9g/1UNkE+7AnSxZc4rJxk4dUhChtV4c8fbII53rI57UrsR1ZZFOr0RZ9q
6Mrxf42rLcvxA5bnyjdra9zRyA3RdydjLxKHDedw9k0hhErhm0b33YRdmXo3BZWHjyh445sAfKDp
LNp8LYOOJAkaJxcNl+YWnDrGubsHNGmVBx/dq/opLB+8KuGRjtmFTOVxdlP4vI4gpbEvrOEZST8I
nj0R6yLuNMd1IwrBUYIukzbmlOrhzMx4MpKO0v4PJqpew/bFdU5e9+haVke31PQ2BqtxIX2YUU5H
MEvNwKj2dOU3F72rn+350+y6oiWdeHW8uzdiBVJGYPCAHiXhRJfokbjN39S4ggid+YZLYmS8cx0l
u615Rl5Wusn93DlQ0CSff6E+06lXp7pYPlxwgaFwG3ncCFm2lrewHYYKRqWWVeYiWBxHgSwUgZ++
//wXexhUiep79TAIdUHVgilCOC1V1ufYuPDE2hN/nSfqaqldPjgwgFGBuwSAwzphv3Su/4IVQNFg
vJqeyQAOcu/UvMX3joA8En3DEFRx83gsscjmNNiLyooucog2zf2EDLfoDY3ph8K5QjntmgEgUSgV
76x65tqUFQmPhOZin1ZlbhL0vZ33kEe4/ttFhZECWOPBAnXYCLL1u4XmgmjZAjMUzoKDoX1MvyMD
0dRrt18mEPBM+NSlMKKujAbKlbJ1MnRyfbaVpa5rMV84S+o2yEz6tPo/DfFRutcQ1NpIL2dsNPWM
KcOG9GKbNUIImt3hfYup0giJZLXRT1uQhkdtJUlte4Uv7ESIfG6RGLaVHyFRKK09CbzXDbG1uARm
ZLl6WrThJ+R6qjLe5quo5LDJ77s1ZRFvlmR+I1/uVHb1iJEGU4vae3ajKrRoDjxJTEnKzDY76FVC
BKoJKBigRKhfzhBWG4Cg9hgnOOOsOWH7hj/8k04omgh7cfao1Qmkj+xLUpjYEEG9cKHu8bw4VTEj
7AnjbNk84IVQXdDZ43rpwO5pPeryO1Ydxwm5Ej7gsAzpb6WgpwlAeezk4svdKCCG+rQ+ctloPDOy
k188heljfbcS5AaUcwZ5Y7dMm0npyi+bJDo7D5fZ5sgnet7o3Zv4OfE/shv96XiWsCQXaeioRFe9
2zpIK8VVt/SXfXULx/9TVt7YyD8M/DSsKXxpdUeGgbAYWrK+cQV4ikc1EMIICpcxx+cjKhg0ePhp
YiHdOmLwtsFsXIVCQr7SEBmNXd2dUUPVAdhDiIlcWxjRqE1VG2ZzzSJwOUeEacJV1C3/j1BJyakK
i/+4o+DNaXBlfB7C5PQsjN9Fr0njB73QK1ojtIuHWjjeOhJf927uVNfqb3EB89E9HUcKg0fA0Pfz
vRIsEfixp2V1Dvdfrt9VgE5GN4c87MyHDHhpuo2YhaiNaXauuTgwmh/zTKJg4Ha70XFWT69bhqDX
zc1VgcWcx2G7+pIAdzN0SL2CR+qcLqpIZam5kWFgCRBrLzbTOp6ph0gkZH49h83LScakkT/DesML
RKas0u7Auk6NxgDJ6UiZ8ahQrHsN6o0Buincvubc0liINCFC7veIJbJh3DXxq2Cvl9FX1AVIn42o
JTLOz5jyhw6Dna2uI3cDZJzdXtbSW7Kb1yPonegXDJVQCLa4iWvG/n+Q4lR+azutULLrvUWLXx/a
QzEpixmFR+HgzcftDHoh2GdR8k7qCn01T3kAeHSsqsP7ZETv3+6AuzFSZ1QdInfrZF7NaqNp37OH
xlWw1qrZle1o23CUW6b/blWjQi1gzSI69zmNUFPxQWEyuyY+Zg/Gxy2AkJIdxck+8dg1ckHG6NDy
v4DQ81vhHTbvj+W8kwukwo/rjqOf4CeiHteSMeudfFjeoLkXPZIHqctBMp5DeLggdzlV09+8OXBZ
V0XIylZQqj+hmLb8Y6sErEBhdey2b2bURdc5UACtpvNzbGnTZlJUvG3Wk38dbZ1W20qi6dKG+gii
nS6gjP3ZLCQ0cwq9BrRFe8V0UiK3KqdTJyGpKwc7m8plemky+s+T6sLZ6FDW+rbY37YCyMnD8Gf8
wr9u0S5/X3aHI1jpuoDyaVO2EueoAXDoQe2ihYg8EflbW8iuOtO8FN/k9NMSkkmH4QiD9v9QBX3J
2XPko2xMn3Gzo0y0AMHiGKlfsOF7m07A6c5+Rp60XqqpqIezBqvX/5tcVxtIJ1Q4LWtqfzI35MMx
HMTo5L+PI/IZ37dpKMAnqJCASTujeRNE5szD9qzf6eH5yl9S1yPT6lVGhWelUh0WMR2jwl7CbGRN
xyDRMV7mgMj29nAW4iZmB5Il6dOJrq08K48vu0FFm+Tz5EnznZ0dCZcW5/7kX+uOTsYwdBGXaT9G
3YcjveUFZN3rHyVZgu0xT+RuvrBTKFsR6cTKW+rIk1Izdp7dxOV4Bm57j2t4B14hAITt8F6tIHjO
U+S0oWpuuy6QmBppQfjJiyqTcRXTiKjmb820rC4/PyJ/fbBQsQik2Hh7x49SAPmKlQYnBJXZiU1I
U0VmEYxsR09o3gfpvmHHhFPJ5rg6cOUbQopJz97MBQJHlaisn/iTFnKvNAN5Pah2cM4RfCMDwJgP
CeTN1I86jmOfpNRWfPguFSP61f5QMZHnBqyo/tq7CSL0kf3U2De9R5niywi9NVdsQpBamYpllzmf
sBe6daoemVe9FvHUjzg1cVqrrvIdrUuFgDE5Cq3sCKwrFJ7yho5PrU4Y4M0Pb8aASAs8BRaIzmFv
hD8350s2ReOTxW6PcQd6US9LnaCeiV7FH+aMXWVqVYkpRvpWfPXZXbJWYsZA9hgVH1C0WiGfwwYm
i+6wDwNhoAseDUaCyorjUN+5MT5rpsG2SXlly7gLKhzOdXWaO830qGdOMpo4JCz4ZK3BhOKW24e9
OOJ6Zcq5EMkpbP3kXHtHoi6yi7nz9xyZMtcHWMK+y5AGtVSSat/P8gb0m6xuj6c8lv1qiZ1hzFTd
ow+bzrD5TMRjAkuY4DWk/FW029b/s7NevE+p3aAfrYWRBkP1zP/lHE6qZZQX+1wcPq5+wpVYf4EB
wUJdLwzqEHwB09hf4706CKVWX0f2cLsKRL/XyDCKiB7q9R441331ay7HUuNhHvONwJ+1fbxJ001Z
Ye0Gvgu6m6uJmakqIRdxKbP5CCfk+YXazs9hgRg7ZavbhsRL60z4o2vusOKsaxYCQoqRZxZNXoYo
J8lXWUbko+nhb8VljxEF1YC3Gukvx+nOSxw+JBWPv4Xix3D1uou/ZxjZLQeNifVQrBEpVdPiOBIj
b7kHovBtZBWnRxlYFqH3H94i01TkLFRjwv5cH8wqHh3sHHfdl8h0puaQprEK/2UXSoOuKQ2SV9Xk
UjpetXC8EP7aE4ewhIRWMwuZ7P7VZeDE1AWXnrTvp6I6yKRAswMUi7G9yBQhZjjby/Bz6TCdC5fe
+qblI0dzaUgtOzEwmAD7P3FVp0RaZ4+qnx78GTPAtR8IIDShRt3xjojaruK0kak55bLWcLIPXn6B
wbp454UjaW+BX+u6/DkIgAvhE0r4/H8h63HwzaFaZKxZq6E8+1cdTmUMhap3raTnzDkahbUx+QAk
3KJYB5HQYZ1Qagw6+89v6xhLPgcIGON+BBkhU7b0ISZkNv9Qh91kQx4N35dUXLqy3kN0fId+qdAU
w8FTSagm4fGE9futZcdX6vHBX6/dOdZAZ1zCFYCu13aqdnp7L1PgwKjBU9fkaVFMwsxSjUUy5Q/m
IAGRRm+GCJfiwkwBnjALanagB3B8E3FHrQSv8yj5vs3LfHVG9vvEVeBjWYDtP0IYv6u5B0iX47oM
T2U0lbxXjYY17xhAqAq3nU3O4XGYecFpVfB3iEDHqMYH1X2ZBAWdfIfXWSnU5/eKS/lMPnAp6wNW
WwRrcvzWPnDbH4ffK1vwl4voaykd/vivVzNxI1wy2o7NMhOmX7wBSzL/2KCmsaY3ZFhYUGVZYTGf
uwYghixAnrlQxO1Wa9FI41kzkukGSfMrU9FoQ95wWWyN5PVK/2sE+9DJWPFqUMMrB2qAF1aYYu46
8XpR8MlM3SmGW+Vy2NZL5cP2IYRylggOMpaONEYzEgR2kKi7Ujy81KPQoGRaeXw7DtesQM8oW2wq
pm5DKkCsXJBVOmWSGEoDpwVEXscbJR5lZrE96zQBFCg9soM3wEumVLWH0sFLYKNUSK9sydglbPDq
XwLcPf07qRyHi0G0k6vGQ/w51UGtSuIZJJIYyjKT3CBKq/uMsZbWo25WgMGOc4QdZW2eKWyih363
X9ly3YhdpSRvPzsoJnZty/P6vqJVQcHPH4wP6SgjepwYKiHptSz6UGqeKhDX1hhfseJEVNOm/D6R
/D1VKOriUTLr7GIrAbitd7XArrGPmjdjxsX4IkLjqAADtM/KpFKILv36jlpn9kom5ijl6ISLlvDQ
VSWTjii3+FydVN3PQ+3DRGT40HRW0Yt2vwGeakvx3O/rLtalQkA4QHKbT//BFu11keqvRP7uCoOK
XYYRZbSF1mvvdHW/XA0gmqfnhHBz0vRc1xaf82tdE4rrJqKv4TdgQwG++UOqhMn/TN5cEhNsnJxE
7jVgWPGq8imFuYWh9vRDXNhLpmOfm4ZYPDtpSfx3O3+kitvB+iMtlwtI0Te7KxTSTdaJWc5LMy/7
MZHLTOGEwA8UI2AFL3vCT6nsezhY3yrFUhajtHw/uR9NMtHjtyZebo6R46+YTtKIOJJnvIcPuDlo
xF6989VgG2IM4Zynr5XY4Ecn+NbQsFnV/mfcMmnQbTkQSoL29hBghwo591vS0t3YbLjt3tuTJOy9
trnWtAFMxOoLELvp3dYzn1gE1Yj11aPcRnLb7U+bN6jt4TV3KVRI3AthnrP8Rv0uFbZH4JD01gC+
10P0AamxGbKHlGHC7FaWZItlS2ObBJEbAyuQLu82TcUXCvJ1Mo86hvxJ2T334Qw5A7ZZwVq19lXp
1s2V9X5+qRGY9JHmNvi3cJgKmLK4tnlJ3Xp/gVCF4xgiBQw9o9/HoZV2a/DpM9gpxN8npFn4YquK
KEwh30l321mgeNwPzd5j+zuWLPpYHmEId4+SK+toFFE6ezwUqQFAYelrBdmrbNokAqDZvNUTtLMV
BFwzeEIuKmbqZmskTjgtxwzM/JPynBILInxQtPA0b7RgPQ4+SOjttTn5+tKmhlZaBJt23lGfChMs
wIM44tgsUBJZgVZZVe4Do9B5ALs1HgWSdQn5VuYSVCHviL9Ksi8ixLoME/8EIorebQN0oXcP4otK
bLoYpPXJAMW4QWmYbZkosxX2SO6ecpD10VVEiURNJmDVzvtvWD1VNek/ifrrK7lDhJi1Tylhoc/Y
X1EOfhACWZYeO+wS2xqHxfIYWBXBu4lvsG+MosKAkkgpqpPCm7fZ4jHPqGT/EgXD3x4I016jMUGA
6kRVXQQ8/st1r2QVkeShhz7Ho7qYVFOhcby3PrwmSaaJl8ysOs2yzMBkuYMgWAM3zQ3FaY/0F6r9
t3xioMIb1O5sqYFOUb+WlqxYZvaJwBKThyg9LOYgAp+Rb1Gl3DFZLuOp+m944tR8EcbweX/6M4et
4gozGO20FvkMbiz7F7JvrMGd1/98ruE/S4wkcSffwQELbo7iUALdCiDJMZe2yy0LG7wDjYkPxF8y
ms0Ss8jjQkw/bNXgfPM1cV819osKuN84YvHlWj2fGh42W11YH1wiJhxtS15iuR8P9cYKztBnSglr
zWmF2JMQnSFXaEWLueOXA7618I385Vz5j11YTCN63g5S+XfbAF60RcZwyHvkKixSLPzeZvGn+/DO
GPUwV0FC04zU2ibCgi/FrmINoK44lWXa6SuPfP3cbCij0yE1OsmKDUS/qrn4CEiukX5XOEQWknXJ
yw612Bigc1LBYYFNdNldFTwz8+iTd9+onTKQOEWHM6boYkFwQGcSi3cTEG5OAILbnknSTe+xVYxU
4hSGRdmFklfle8IZLVCRdVPltvU326+nXkhenSlHuTIQxfeKauJAvgMw/Ezh8UfQLek17tu8WMRj
DyV2LWycQSLRXKwUEg1reFUUpBVP5V1fcX2AyJ2pAwnYkPUNyvS00VqSKXoGNWPmduJbT/vTQVA6
xh7VomxPiMc7qZLsQoaS95LZHjVaEbvoCF/17+OS2Dc/q6x6NtnJjW/eBqai1pTqHSW8jDvxCGOG
S+z046gxevS9HMopuL/1FQ1rtmp57Ifnnq4W4cuI43W3yEpln1jLQoKqf+wrT8cHfDJTP4laf+zQ
MrkaJvu2QWyY5TaDHt46wjsGClpOLCxwkA1//rClNVY1RZacTW0fmelwlhEilcYXq3Nnvj9ttLtL
7rRiH6OF3UvCH3lWKYdPqzPlrhVqf6UJXikl5nu5HWreACL+h2FJXF4l65hmYov/mbuknxCGCm4o
0u0EvBaTgJ11D51SnkcZLME95mkEXfH6J06E8XUnyjFuVdHhy+35pgGRMLqfX4OfukswAy3IUDES
IIrdJtuAUVCIA7e5AEYRmzZu5k2tTPWanez9rO918NKz3gg/wOrPcDyEml8uud2v4dwXaytNtNmD
YKj3NilxN/q9v65GLLWBAqdyz7viBIueJKay6ao4REe5Hij0ywxPwv3Di2mB+TcPlPCw+rlTqXp0
zzLEmE0I5W1TeY1np0RuQljN7FUXYDuRE8hORWTVl6+rmTB1RqPnNWgiXivoenSjWe9A8sY1bM2S
x9iM+OQrPZ/PlVx1MwzCbnEmNfH5ec8JXgVTdNkzhOwmkjXA2WGA7LsoGg8+cxPE5slKwUS391D+
r0PVX9mwnrEn9277A/RGS3MXrRWt0I6Hyyc8C0I2ZmIbPj88ksD+jt+NqRjaRbaQCc96PXcBo1AA
ubGpFY2CJ03aN7xNnmvssuiP5h2M8s3YRdrVmW8PRsAgGEzxmxUk8sVgFJuqyQpHoUFgCxFrFBtq
PUs7hejuQIWrHEHxrEOz0/TlYqKKqTdsZRks32/4yee+hLJSjTy5SkebA/IRR5ESXVWBb0BaQolR
RRmEcRaktF9iA1r53SfzA8bDQYb9eO38R5w4eA7zzpCRsueydXin/+FFReoqKO0BLmdKlKdMBFmM
Kl7CoCluqoQNk39Jj3S3JT3FhoDJ2To8XYxR+fyxi4UFOQXlwv56dXRFlGMNrQ254C6yDpm247kd
ylmRq+aQUITB6xPwqaRCBEfOsK+MMqZzQELnAzWLQbT5jxagdA179249TAdp+c6y3nSpwhzITzwF
WP536skgwC0HITeIjHHBG01GXhPLz05zaFxgdU2F9CBDB8tqSd4mq+jvluKZ0qdUbyDtps2F3C3q
jY1IvLftjWoats/o/nUFSUQLXb7dpb2dyFsE7GF+6d8C6gujuDrWX+qmf7VdyMYxNbrSjjxckoSi
aK7PxDDyEdBNyFKKXjvEHUc/xK+iX7eL1FMK/BLZlBbcGZ/d+ksuJ4QJ3Wt6LQExwPZq+IN3BD0Z
hobUilEajXP0zYVARJ7FaGKDBEA01Ze1NHyu7rRSwXtrNHDWVPB2vx2FE/TJpFh/CaXXoTHClDHn
oVCDN7nzfJLBvqtbHRQ5XAt00lHKYUV6YgWb1WWedFjdcGTNKqGiH8FeQ0hP0yQvI7Gnay9ab/HE
snAjw1qvVPyTCxSESFAvyYKge9IEHml/UdcmnwG/Y5RZQZ+XxI0xjIFzMWqeM7S9w1ogKIl4nw6j
uhzkllL7Ww1Lcd44nq9TIIEZed+tctXt/f40qnw99OqfbLO8n0LQh4UV76wIsignesVLDULUEVF7
POtlOVawj+s6VWJbiDWxurpx4CH0xR5GATF5KkFWmacQWNtyAkrGnod9wifmK27z4ACqK2L6kR4K
kM9NDyfabFOCcKy9RLyb5Jkr81KDZKdqY0IFnicpRiZUtByuY9AJDcSKtDHlVL59AIC9iiB1b8kx
ZI4eQ6K6L+cR3ImxlV5iTU+dfVhtYwwYR2Yc3WEN7m500B7iYlhh7MwCTjWgjzhHKb+pBX5rxzAY
H2hDv4ZX92579yoXzpXzb8BMCnSl7XosD/uz1cj5Y5So7uS0tptJXEDfRLGNwrWvpF29z6o7nKiP
MpImewLzYMRSeQaccFYhShe73PeUcmQ6MQiJCXpAgyA7QukoqebtXZUR8+dWFoaQUIoVJzPy7+b+
H7GFBBCIISyNuleOkypQVX8/13kFb4yzFPzBJbM3HcyJxZ9wXKa4n1QU3mxdtJdJit3ZGt3p6ZMA
10ir1TgFDPq77q7K0nFzZxpMGO8/RoxRi0OP7lipO5G0oJgofvDd8tZIRB5tuP4kDZcBn7cT7EqQ
hbVIb6+czLvhLhKZY5YazpgngMPTMJ2fz1ydm3nYIG+gItj9ViRIBqFHL/pAeeiSsobBli5zklUW
aq4b6kX7GjaY+92OcDfGxWpPzTIh8RKC6ij9Hn9Rq1ZXfObWFArZtbxNOACMcHQT2KaADql8a99W
JRyH3qr41xbyyoUofR+Tr331vkljx2xgeY21rhnQ12ZFXAqvdWoYdp9VMETK+AUtim/J0nhuodpP
plCJbmakLstKgatFCiYnwUckvX5ljiBUmGrG0zBDGY0K4fZZ8INuzWq0MJpGjGeFEzuwVMBt9wkM
GNzk/LWmW6VUn2tjPP5IBtTnyp8kueOoN1+RrDFXS+1oTInWdiqk85JPneIv0yVrSRso788WgtDx
Y4sRTcwOYOm1Ol8uh7QZzPDoC2hJII5fZqSJU8soO2tAZZUk22S2yCVyae1jEXvYtuHM3WTwYdF4
WaUUcGVjfd1l8zt3UHhU+HXjRDyCQwrvai9uJG7y4KnkTPR4G2mbHLyTyeokZmRJw6iwuLAekvP1
ZM5KGjaIFsY+ur+c1zB21HGRqhZFIhiQWFruIAHDlifPk5fa24HGH2nFzhSfoKGsie+4hSuc0Q6V
XTF5tFaObe2rToEm7qJ5MSWHQdnSsOL43nqOk96Ixsr/9Xs9vu4Rr/6CI+/G+r2l+8yADht5Q20Z
NUrGGJhUPkZmT7/ZdLd+1liLbQkhSMHF8WMn2GII22Oeqvc+A79VFzSwLES3P/Xy1dYlAyULT+hc
VBZy9UMVfaN4Z/WfepdWFkwLyapiPRLPGBtfnmsErdxdMDj3rHkQU9cZWeGGMR+tddMufJGVe9pT
q+aLQnTfSCpVZh4gy3I0joxx/RyOhh4zPm8WlBQe7QmtIH4QNVmsrSyUuWi0uos4CuU38AX8dO1y
rdqxLn8HjNMX6lXAM4Z0/kELLAHBt1B4eHslbghsXsT8iXLS1VYdhmVG+h2/Gjq+Lb22qZadP7Yc
86Dy4Ac5VMETI1+9uDnQtjeUxUHRr7dumKU017jZ3MhBm4EBZmVp8HVFbTf/lW8heq37Fm/JVari
XPHoLsfs6U9WeqWpDzm42uupvA9QOFufOYvQBsp5gwgXP4LeA1xOTPren0rIF0q8g9jlnBB/U8p+
qvZLWOtawc93zInvm39F2j3z5XzWQrrzEnHtYBy5Roa6drrkwIWKkNZh8G/FSvzRwDPAgbqA0lYW
nb7unc43TMwOk6o42VL4btL8bM2WY0etTeVTJJJAHiVFb10ZelgImmsZd5IAIW/89hgRWLpxnaNZ
rYQa8tJUh6Uvnltmhvwq89e9Ik3B1KKD76n+f1evPrGNSR719MtySVpuKS6inpX9Gv9bGM7vCIpu
zWZe4AqbAt9/oczAECMW/+NEJ/OA7Qlx1p8RUtMm5JwvGWRc/+t6PJQ2KZ81j93Z2P9m4n9Th76V
jKdND6HchJkTGaiL/CiLfQ5but3kUT751n6jTPRalXXT4oNdSzvP6Fta2OJH1qTtc1Mkv+G/VgIY
81+f70EVMR67/fS8aZI6tLbaGwOZJ3t3xyUcdVDxucykQ3a/5/GJfo97Mm24xj01n0l3UNaH1kUh
3J14XMjQ6zaM7o/LEjk0ZyyVtFe4Ppeat4s5liBw9I0q5Odnd33lbftbHHVELrmnmCv741Iiwb5N
TWG8aUtl9NOaloMzwReFH0XIZgOTrg7I8Wo6QTGEL4U53mPHCdw7Yapsu8w+QCZWAGds77t7p8Bl
yF6MpO2X2VPbbo9MKGBb5ckaumVL6x9ePpZOS5B759Zlel00e2MZGeENnNSa2PTsCKQRCLpyaLoJ
BcmAGY6Ij2WFwAyLHhZjosRKAEG1eRaigaFo2aZ5DixJXEqsg8H+DDNxZRLjnfpL/99ybvumFGku
PU8trvXPabTlvERBUpUoNVeTj5C5Zh+IG85C7sCsXYN/zRwJUQKNK93Xt5aJ4onHqBuO2UIVR8yZ
6G5cmxMUc6hDufM1ODbnoVU/WZouHHctqrcGTQdfiz18hZunlt6tJlyphZNSbvfR3nvSA2xMKZnL
zIepzJk3t3U7/wtizsUuUUHg2309XN0LM+jAnSMfV2cnwP0T9Ay9fd6fCG5/XsNmNeCj0eYEcbEV
MklmF7/Uop2DbUQkwP5XE3MOMHW3MvAXAw65S648S4f1url8r/kp2F5SgGvtsBYb11EluyS4E/dw
bZkY9Bss18VoeyFL5hJDL5hAfLOnxD2tm1iaTN0F2gZtuq1qbFNkp8xCzyKe8I+yZlMJUniedfTJ
zTOXauJjd2jiOqMAGgCudT6TUzey/PHPZWShw7ASJjL2vNwegL7Yze56GKo8soJeSj9m8TNJTtnM
Egt6QZCwaDchUdS8hqqUui+2lUMdjTEvL1v41qP4wwM6uSRpItAw/IOcXf2hzZpebHWfKfJNMo40
W1+NhFnmoKY8XbUNqrEYASS+HRbn1fJO2q57bSubizNdihAjAVwL8DDWAiFPS5eJ8haEXlje6uDA
Vz0PIAxW7aNzAES8jOm3CXlCueMpGBLvMaWDVfW70ZzVwYghSpwiJhEP5mLkfb5HF0eJpW7TL+3o
kLoCXJsvLj6P8zuw4x1gI4eX7HEQTe9Bvm3Fjpupcyzf+WLjtu1D/CxIPtvxIM87+KBQQvRUgCKT
k66h6Ymosd4FXaed36HfRAWWEKyV+EkVGB0kfH91FC3u8JZkDv9LstYosHtAXmoNQmWuW+Lm4vLA
Ie3GdBxGpUlqIdpLlVtQ/Ootr8OYTVjaouqOOvUj+O2+TfEuhpCk3iEaXg7/z86a/csB8XZZ+T5a
Z5xXEKpNdh3j1BFNFAsqblTpI4zacnLKXuZVJqy4dBbvwUzqAQXfUf8HkhmNn8GA+lH8S5XaIawu
ojuAcds0o9mM9wujtq8R0NhnSo3itqb0VbVy85DnwMNszO57R4lcF488yDwoqhusxqB8tPJepWdq
CiOvj3L/327HodnxOjK1MbepFrJCK3gYfSKRpnZ4WO9II+bayywI4e2XqfhMAp5/go50yRW/oi+0
kUMxab2lC3XS1TwwqWs7ybp+ptJ9ZxXmbsQN1rZPA+vgarJPtgBipY4QEAVO+I7Cwz3gEnbQTCt+
c0vQJjWbhnJAAo26glr1CXuFdWcGqADkFV3FFSA+udgMS/9TKSGXBE/AqmWwBfZrJsR/0BXsE3zh
hDwaZCPHWLuyxnQVCFrtsi+ZwXOF1rUfDeiq4KFZ4zEzdzdPpespUqUqaGg97rDq727mAKqvKTdx
Mn+lhnb1y+0CqZRQUoOa7pPc+4/8CqZASifRcbz6wzYKlM4dMQSufiC9zqdq3iT8XuIgbttQTSYH
HWRt3Rf83j15d2JrqoWJAa4S/J77YUD8pUkI5UaQPPkvFFPRQoP+mUSIWe28mcdtK3nEnuC8yp/G
uZXlfEtoTC94i9YDD/sXQth5yioYvT2UkATkZGTEEX1ss6FkhtR5+q5wLjwdo0IYcGeH905rlqS4
cycMhQKZ4CBPajMoISs6pvrqBzMO3fKdxANxfRSbz5AHwfwJ+2RsvSaj2x1kgR7ro/3P4bqdVhEr
F4EodN2KztVV2KsbfAmJAPievoyocQdxgO17INYhF/WhP+vAbqnDg9c6daPWdOoDl/hMi16lexN2
oYrmtMgtr36YHPGFeJtwJrnMXL5Uju/bs2JdyBCdET4WaG1xOzopGtDHH25I3obWSyg8JUzjE+MM
c1yanvpse4x386OvBsfg+D/Z89uf3tOjnLDT+1omdboCu11Cg2MxoAt+Toq92EFNXtRBrG3v8wl4
RLoxcT3vk6DwEa8AnpcG/Yc4IIR+R0Rck7RoIKvs4hzIPm43C4xY/2J4pb8kVnKcauw/FmNDx+bk
dPRKt6dI2uqIjDM/lRvvSbYHfSAB7aYe/Bm3R0WOZF+9QzzSxjb3M4JaIB8x/IQH2+nk/ZLoAUbt
ZRsg6ru1z/RS7kJ7PZV86SnyRJ8THMdi5m1tSXA1Hd+ya1U5+uyzG74sc+SIRivqv3mR4BmEGXEX
I5tserxZYym7WfbXup2aVgDuAIvGL28swizcRUP7w603+7cuSAhQBGiannkCtlasOQpAcnxZYnEJ
VB4vK5/UQCMFRzuf+eogz3WZJMZ+wv/ylUrFJFLLGoRfaSDKHjFim19KjNCCq+FI+IYQ93Cm14yH
ccQltJbgqak8NocghmSMcRMD0kq2zclrvDLlFTkk3fq/jiCOv5/GwUUChjdYICBJDSZ9IwvXEWpl
o3E6oF7bXC8jcFjwcAvqqJqpLkIqSvP+3ZYpnnfnvGCFLwr+UQVJ2AfP8ksb5lZTGXNTGVTlshdL
G4rOw9xEPamwa33REtJZlK0mU/9UPBtRvokpGCmDRXNONj2tqL1ANA3r++YmON1zftBxH4lt5Jb+
MjvcG0sou5rb8UofGg67llP/qMANVsLTo45kBChx0Occ0ckZHFiWV7AOAa9Sp9Nrjm/AQZW2haYt
Gz3Zihh+HpeduT06CMmfyiV+6IbBDz316Bv4YLCDZ8mTxmnuoSZ7e9GysVRafuBBq178oIq2CfJ4
Zoq3g5qxo1LvNObMMtnlIWdYF4EKVKbNGXGQS3oFBWwEsDklFoEnoGudMKeBQsD2ihAbbxFw+ydB
tPEzpuTl6TNNZPRQIhTNTSwQpDvWyBrj1OVffSFkzxbGjyOeClvhdMbdNaqUsRbwhOfLZ/yznGhg
zwqxzKdSsqsMJdnn0LksexVDv5WJwyFL68aLqcnLcEmQ6TZveWbfYcp3CuhYwBr8DQ1/ak8Dozcw
xPcUcADc5pr52kdZA7i5KyVQ/QUSMYQwE1gTUrSeGyU+SsrnmaImy8KXwpi2SCsP54cEVbu2vlNb
GzcLj7ZzLXY2r3vu+NkxAhVA51JM0yW/+ovjnecdzBk9XY47xLe0OHRLtkUUIZu1U9cuHT6W8U4h
xmAc87Sm7IN62SCpxZzFMUMbHmahwIHH4YTOFHiUVolzdxW3PEdBkNnGGP5gNI0Abp0Gm4J4FgKb
wZmpJ4HQPOiWLCvTaLPu3wIRj+lBEl471nr1NRitp7kJPBcI5MWgNIaKWl2h0IfW9gK7gMM/uicC
R4uibNHFueBPhz14FwrGusZy6jiZW9GBynu5L/YafBj0uNwcgFRJrrWs9LI/v2pOPYR4hgS0EPAC
IVmCnPOhmVEf88wcU1HUTy7R/lOJFQubcHKF7FnLpmWZFgGfUpusSbbnQh61pcRIwxyVUMpnFIVV
Zv+mtX26DIGo4RBpCp0DJSNTmGKtCv9ULjUNiVN2llZeHmhwoXxIRyMfw4gV7C4h+gJfuZfjKFo/
RGbKqjNrHTi9o4bevaOGZn9wl0DlZt47/DqQ72yy6aEEOVyGKZBMpuiJVz7S795gqm9TRwTlAmaX
iooTJiR35hMm7h/ShIrH2CCQQ1u7y5DTcff5J28i9iZreeX3Apsbl5CgFiLR8846M5nBWnO62sA9
OWf8TKW5e2lwgXVh1h7dyT+1alIYQVUiqNQXlg9ZZbdpPGOvVnLqpz0jYK22bpVulr4pA99JkBrJ
1JodC7QQ5gJIlNocPAWvDqD5jSHqYGNDK8D1V2B2YuQ06tAAKRUj7RXd/WEuUAUychkLGRPdW1XE
ir4zdttGdksQ7ZnErzaq+qzoZkBwp1JueLXzyMG2bSbtaTOvQ2cwvjInCw34/AI+MN6X4YG9pnod
sT9xgXNX274GD/vevwKuV/gxjLnpH+NAOVc/tOwV42YkIpJdwCwrAz/0Q88buGOlchNSh8D7sH7n
79Lpo3UkL0XHjBSq+7ORu4y+nIhwmO1a15uLjOECTMUIRIsVyBGgKf8K2zF5DcHgJFOwCoM1nOqd
WLjMH24r7STVu342fD8YUPa3SwLVlpecbDiU4g3Fp36g2BABpq4cmKJdwsv7/KnxND5VAxliVnMI
HGuqnpR1lTjHQeBqv8B0+IpBaxCwXqmTo4ACNiMqATZORL7HJr2NheptmEuaLbMtGK2SwMlGaNam
8mdAmwuEp4kcDxJS3WfrtG4Ks53bWA+FUYxNolrH25+KTbAbn1jJ9RVYUP75Cnr0Q1NFvlvOOP4t
4/MnO4kP5BBOh4bvw0yUtTA5s2gLHlUNw2zAqDPyKnFNQCdwU3VmcugeGJxLezWfELVj21AIhTKz
Xur4UlpXr2oGNyK7hjPvHOvqO0coF7nuD5zAa5/F3Ybjy2RNK9h3FRyZa9eNqWwOEglz0GHl7ZjJ
FltLWpUZjlDZvpjHUSJ+u5qcNRsyOeO4LuEjVHXf6qgfDKUoogUWGvkFT2NZ/fmdIwD494XjWKL2
d7wYm2sVZC4fnB4SB+8YjdUrbAcPsGTbPXBkVR3ZbUt1DW8Xj63yNN5CjFiB4Oi4D+WIJtS0OgSw
2559x7PQIXPqOsFBl3KMhZZ9jatV50Ko10WEa/V0cx1MvGX3QsHXM3Y6xLIsh/A/1HwcLgfxMlWg
rRutxqtmJ4Qtd6J9HpYbaDvOu5sb3Az0g3wyeQ3skjOnR8LOfXoURWZtiDRTGV3c+Oorq5ssa5gl
WULElb8xY/VU8+EAjl2QkuG3IohCO2ezE5ps/x1veq/ioOBaMS0i/n61jYg0lzDLivisVIcE7sus
uJWaSVzgXpUhZ2blZnB+MAjpsq+FXOwKmgrhWpO0zP9o9zcF3TakBf3uOciEtTggzKHIWqVMFSS7
wFIs0XQ503XOH+Ynwjl5hiavUCJobfAyAgRzsJBlUxKjXeMN6kcx8lLFtyE43schmmalcM2ebSjP
Z0pxh2k6onE5k1+IsTT+PUmz8+TjJo38p7d+hQWoQJZxNnYnI8RjzKPC48/cUfhyRx2iP5QK3aYr
YUQGdj7yPZSfeW9GkAAsZIqsdr/fYmoMrBpo6BSayYJZNZut9aSOkMefx6LmZWv/5o76jvroxHBE
/AcuubXA4iFDAeGiEi5TgOnqfNmrb8xCI6NYdo3U3rTnqWKUG6wJ2vQKDURJTr3jmdAyqvDJrtUP
RmTDkFf8J5vWHDyRsFunhE/LEyELQSRjL9B0SCk3qggo7KRHBL3bA7FQjDCRKlv+dW4EWYBGCZYp
nEKpVRi8bIA5tsDPCZh75nv9+TefnXv24ghtOeGeRXO7dUUw8Qv+A9vCy3DjRPxcqz9vZZcFARwW
gLY1EY3LOkIZIHmOJFrbHkctOEiqO7U/g9uAT8hIj2ItOeYua4E8LCZyUN16VGFPXEVOburw6Mul
/1ySqTMFPufSW1RL552dj3vkrYIQUgaroZ9qNQEewu9iboyjMGkx3hlcPRKNJbXy72C6xwOFz9T3
p9EBkpYVeQRNsZ7hTSAcjXwvFtY2s7PXfaGrWaJvgGKv/zIqPzrl5yxmNBPNBrOfTmVEa8bWNqgc
u0ByS6lKxLW27nlhShrzCM7OqSk8U/SwG/O5ID5djOAzX6lehpvNVWH+B5lkmEh8VK8vLgbK2aQz
7DKzh+2GXW5w8RFs3l+rvixspABmZQvaluVYfzfCa0yIbdSQhaDV+I1rGnu3aVzBsk5SVGzo57iH
7mxsNbubI2eRl2C194hYEHB/FI100QlEKC6Rz+jbfz1/abZ3Nopmfe1NHCqKXYSsypGdw+AS8MGq
Ev/yzFu4K1sqqRx4EGI3o3egJFms+KxARmxLu8UpUrCaN31ikmNGmGxnXGV/sRPm386Ce0xTdj3c
iW5PISGfMej/omQAYaVzpTCzkqKrTfAbW0Mtfhg4MhpMZaCleUla8+lPTSr7O9P85+C8w2LPirmV
Rc+fzL7cj5xpk61is/FbFy86z5BMn3k2QCtTwb0hkDz1XFP/LoRPSbPdvYCtbAqrBnrsf8vWrR6U
3ofUOkOoTU4HQ057rFSTZZN3YW2YlDRKUhhL6ANp0gzpedCudQv/UC8U5q4cfvtc4lJMk2IHKTwS
Tup3yYvu7t0IFP+uD+KYHsNKE9cjglX5LMJWm/8FG5Zb0/Z+3kWufVn9C60nhe63z4zmdOMuo3FN
6J4TcXJK0ziwDPZuacAeJq5gDtZ6rrFStJM4oTfNDWwnolsti2Xm8Wkmb+tCuUuBZQPC/nYE72kk
2OawjrSunrAd0RYrlq1rLZuwx0hCstawVrTvGnNMwmjrn00UJGurhTPhh8uajz8at6A7DBQ/XJKr
cSSE3F4vZZwrhoBGO9rHcYCHovU9wma79UVbk0MYmF/g4tQxYAS2ZV08xx8xB4OgInx66ZiSyc7r
zUZXqu2cAUxu/cm/i3K6zgqSwe0sc/gexFIWLZngZh/JyyfZeNny4H1n1YcUCr5XwRUuxzBt+sdO
CekyVVyBsvgTvDmJXxaraxPLGU3SbbLZ2Wyjt6uqIssEQqFb2WCrBEvJUNZdx8k2mOsdsV7IRmLz
Ol1jr76/juORFObZ2xj7XXVKoc1ZcyYXhIcwEpfG9KrUR7b0EAMvCJ6AZ5cs9PufS2XeaESYwny/
dIkuGs8ufI7wG36U79il8nZXJBIxO3xyo+gxWfYRKEqBKbQ26WQMX8KMJ31t4TOYl9Xgjg34tLKb
v8HYuB8PbdRuElkBKcnjqNmQrzmoanlwIl3sxtw9C01eYxbhF2BC3aSU6/0Wx4ZDp8OX2MZlii7o
J2PPYoHnVsfrbaGfm1YESkx+91cL97iBgqDZMugPxUCLCppGeF1vmEu0NvLZSVFF2j1mM0hMONyI
9/XGFoWPRs5JXtNq3DOoz1zYEhlIFvP9UiZP5zx1i8XFmfrO3xuy+prlzdDKuhld0h5cGh9Vc1SP
sQEoLtQzZoVVlTYKaBWvHcoZWbKNmBu83hi51UjFQTp25OUXtS13DnebaE2lR0WtBYYBHPbcox0G
8bo785oY+6vuFWg7ktMp1i85MEtUZy5eOJHKOf3htGjrNDCgbtRyNXRkpsaB4GgcCDONiEpWDIJJ
1nI+xCCsKJUQJxZHSx9BVTtwlC0S7CQ1XgOYoN6aVLtNfBsZiCkoyhXOPCMaOdwMMS5ArHGeUTc4
fbWfsq9g1cPM66elZzlkCBXXX09p3OFg8okXyYt6SmjkvMCbbqyFxsQINDgiFgk657epguqk7nc/
Y/Wg2FxpE5xawOqcE/0VTo7yXjwwRrWiqEMMj9a781pRflyxkL3PJ68Dlhg4uzaRVN1Vso6q+h4C
sbwBtekb8jJJUqgg+1kH/+SYXv2Q1bd9Ek1ecudSQ0JO0bQu2U0z25wVLqOQ32ExOpQZZPV6OvEt
e23xQjCoNpmpK6LYEg5Fs6YEXU7pgl/BzQYXvtwGKT3xJ+Zkk1gDk3ni5mvjlf8UCt7aO/TDC4Lk
mxsDxLMR9QZzRxrBtIFm/tu76uah+/z8Y3R7CGUyXoFWcxiSFKAjKR78BvF5AiuwlMfxeKvk17HC
XwBCBSZ9GNwJe/QZx7Lu5pXbgHgz7DSaq2Elo0Xeaqan20L9KTU1mjijGk6uq3iu9yURgEpBWWbJ
U5+RJlHqkkHKfpdl/qmX63MvhisPgZDETiwKd18T4j67vO1JgsPF/S4vKH9zWFNk0nt1XqX6uHUt
Vw9Go2YzzMSm9+CYbrF9oFU8qokFmQXUTpLb5CT71IgHc0RbVqNbEE8otmOjgCndtlMTO9OvRCnf
fSdYx1iRRbGfRAoPP7nVT2sZI1FoZ+Lx6itFraMQUpssYDmq5W8bJ1zh5Byt63/3vqNXYvIAF3qN
DNWhtzA3677ORGce79fwcVD1Ms3xiCcz/rvNdI5Q9S6rHrvCmMWNft2Np4XfiGQUD+QQnmfgaJSo
F1NkFF3sN+gQOo5OMm+2uzbuzD037cvlA3Y937v6mPydb4WlsX1z5EYaewqpUWGeu2ShwriJamd0
z0OYe89B+BjwRlgDOxQZeRuOsvivIDbW6bSotP5PZCYeirdf/h7FwFfCB1L/f27aapTd48SinBN1
RQFjWzzgtYY4wnArZmqOc3uRYEQu/8yUlki3g3zbY9A8MXv6Xh00kSNv6tipkViM8O+8QTghHmvr
r9xx70FtARjYCofeLKY8HHA4GKKEcXoq0i3xkFu7baLIwVpglrYYSmZETwXnPceZcbO1HPSd8ERA
ZoJSWOH/SG0Ve6Ec9N3d2C8quOizyDiBkxE1mgHwjMmp6Lm23X89EXeWM39Z8x3p9saTKPvivDxy
3Nddheo1Xr4515YBpHhqcDG+yD4A6wVsNwM1m87HLl8kW2oj2fvTph1ik6TyzrRvGmmItG4wu8Pg
xTHvI8lYX7yWFXanZaoh9POqJsDoDhpdJu2cukuC1CfV8JEiczpsDXBx0T7pU0gWUm0pn99df763
su4bCiw3yt5jnd5mI+CpAGQlPMey+O8Aash5OIhhcfK+2t/ifiapx817s8ZT9SWyUBmUsiXz7sgE
BEg7CHjuEEu7x+fPDImy9t8r65r11UjmlbMXA3wAyiGoywZdJFR4PFzNvIbwO4/PMo8UmkIbifQb
KVXdSOvrh2gxBFnjpd8hbeLp3MV8eKJmx+mD3Cp7E5gfUgyBZw4BajSi38E4D/do+mkoe392VfRR
gR51/9mhVyQZC5lEDioISKwzqxwhskfCllm0CEeZFuI/ujv2nWWtnRgxb57acFtPB9AzHlO5AJHR
i+QJliNYNprFEYP/UPtgwvdEX2RcxES8RzIiiZBDyeyco9rHZEOBoXSc4qgyit3xGZ+MssQ9QLgf
hQiJCfCv5QIJlOsOHvy5rvozr/WSft5Frm4FbNr9W0tkHLeLIuVLKkIptVU/X/ILukgxCeS8G627
NjJoNUM2MUJlZeEiyZm8ovuGYNomUbjWd+9deUy+4+YeJXQDSDvxLUhqsup4XKVceVltW9tjTa+e
xLl9Cp+632R4exAZLTHQw8Ncyf4GwfbnL8GhAeFt50zvCQOa9+6Z1KZbk+njwbiL/1i504ktHbnx
y4GpfxCBTTwbcjeKXxQQawM7r6MPwlS6rsojkiBdAv1DCIr3FzpCxO31qas+WZZT1t9H2ZCiIz4i
h7IsLVT7akFKoPeOIUucMi3EnPGaMT6x09WTQefLFZswaP1W0zMEHa8BAfg6jRhEohC81g6cVu4m
o7eIFSjb97+MXyglxe22qf1xzEBON9pDrhMnBTkuh6dyi+j3CvbcqAawDe9s75KEz8ZayYItG2wX
kiFe6z7xy6PfaUzVxyoJFvDozuvyWQPPfoZ+8P43RNisMSmOySywDL93ClajlMMXALhp2Cl8b7h/
2PmwuSMQfInQrh1o4LZloZq9gk+L0Hp8apCzZfcWOqiYvv/8vXmLAOjGDBbnRTv/DwTZO4TXkKjT
EIrQXFn9VLmIo65zHWZlVHRALRh4fEHM6snClY4Ogfzj8touo++KQaZPzBFKjS2WxfM6MW/ak/tg
Fgkpoa9HmO/vZnUfhCAAP6nk3xHl1QspG4hR9TTwxfxYsXEUWiug4SJADUc4BbDu3j65eoV1yJRg
CC7Fs8v3hhD0QeSfW3JqNVs9jbUrlva4LISQc3m2I/bmux27A8FFg1RYs6zC6uy9SupBZuILM4pp
2D80LLjZoG5NKvBaw8Hv4ZXVG2ZWwCQA5mYJ6ZrgJc9Nqn6GnLgPX/OhngykUcqCg6ktSxtz/rtU
M7VCh2swF17uoIlVQ/dbY6l/5HYFzeJKlciUE3NAhhXV8pJBZdg6Oq5vyJm19JCCmApsSwQoGfxm
emrd5aQ57QBKzpdqCwIxK5W3/afVKKDFdaCDZJpyfNgKNc4iAA/gqSb1DudLfzHtzYcV72uROBIC
amLlq67XPp/0pkzrY+VQ3GXNbky5vxEsm0VCSLmpoov3Nsfxls1GpOsOB4EBZunIem6NN+Ymp27o
s24xPkXFz1jkdBOoQO06NxMqH2v7CaOH9yip0Aq/ebmZYeYgwSmwXXKmubbyy/ENb9dR8H56s+Jw
vDLhi5+2SnUZGvv7bHuuSZSnylGt0tf9BQ7Fk8kMQkeAKwUQtvO6UzVyJ2JRFWTLiHMudcFXwZmQ
jmVuMzwT1P31vsMSO5tdcoXFmMhK4vSMVt1O4rg6peQAz3mIS/vGjQH93SpAAhTCVxU2nFzvI1L5
BrBnj+aUnmSkv6G7tm0qrlfb7A6v7bXlgxnyjICzr2/2xz+JTHsjscCx0M6E918nkK3wf6YUMQ5G
2XJtJlTGp/e9f78wkrVMzSBJGivpoi1TW1mSTxV+jfhPG1gSedYA+0XTMwVGo5HM5uYvxz6Wm5fA
DkgtFHQKQXSOlO3C5sUkWLZaqwfj1m0X8p1V1TYsPoyqeAf7BjkWU2hpKmIorSVhqViN22PmVheP
Wua70SjYXftiouaK4f21671a6TlwSKVVym4CEu8lHk1HP45QroRwvTWQ+GEIUfUKhTp1BPWBuAoY
DvUC6+cnTVmbS7eioTnN37fRpfPivPaxa12LrIHG4d2ykANQOzvkS6/Ok6OGNSbvH6x0u5uIs5bx
pzDX3mxgqk4cP3Ytf7/SIvfDXpnM9/j7quKcD6VDxAEuNtwZehf7NtoM9nklv9y9zhp1CXKguRed
loGKzj8Bvukmk1qmyhd+sF823MAcc2y0y6JG+ZDIwlldawtDAPlRY33PEMQS2WQ50S93TllgG6tp
pUpt7/RjQqqCjmhfTt5OPvPCMXz3Gu5XY3cHWq4Wxy0n0e2EcLYI1/dFKV/FGgS7wqDvlU3h7Xcz
MyNNKUEe6in7DOs6SvoU5etWhKwvI/C9XMex4PZ/pWENF3noZ5ytiig1+kXyDHFxrwB4Xm8AhagU
s9tdb+SrvDgMB6TLCNb5ElgseMKiGCtcOxUpXoDEueBu1VBvt3g2nrx1AW6ZcKay9ibWRSLzGdeK
ICk2nbDR2PxNeLX4XX4MeqTWM54cPkaorF/Gff5zbm3ITcEQwqJTUmWZ7fWt2olkchJhkXD/2uy3
qezYvU2yoFvTlvia3c2xhpqU+4L6asjjBH8M07OBGL5LIQVlL4fts+K0IUW/A1hAkmRlhjG+CXIR
hC2Gf04/BF2Xq/TNq8AyXKngZmFsReVU7wKG++2o8UHdLeNLUdk5Tb7pmcDi3f+Df4rpFfV1eeVt
CE0U0PXFcyuWaXc/Hq8VJ6BGbRniQYN57BIHulpWoOx7uVhQlv6B6LfeB1Cs7S+UjkQ51lz/vX1E
jzuYISJrVpUpOH0qAnqLEBR/q7mYbQLKHG2oNN/9eSDJ4onyLDh1oSnfS1Voihb2JKqMRaa2UvdN
sAmidRA4JvIJqrx/0p6bo6rr7GZUof9e4/CePyyfQjAIo0H7G4GZG/h1DcvjSl3EodJrpfiTbG2a
ds/8gjXfgWzM8MbtI/HbTPU9L67HOgG6LqxeXnlM4aAsctwfvgAHayemGygV0zFjlXgAB2hvI/B+
gbzElnzOVMPoI3NL8g1fCVLGIJ+29R8HpqWip3T34KU5AnEzXU7DWl/2wtVP+YtmleOH+qVbjCBJ
uaFsD/AyZELjSogCloegjChlwO9/cMnHSJg3uRaJL8JLxpJqNK2EfXOp0ey47DM4R1ShoC6S0PyR
t+dMSbJhVkO0+gYGF1jHYTMnAxRX2mQNz/00dqMiwgzutrODRZFbPxc5K6v0OBmiMsej2NhyAgp2
/7wYxHDxhMgieKSjjxGrjHkhNhskMGUgxuNJ0J3dzBug7ZndITBSbgCezl6OcDOUaktENNjhjdeN
jZxoK7+V56GFnOQS1PDh8oHOgE4BiRQTzCgIrEO7sD7YxN2S8q1LikvUOJeqZ60jlYjZf5u5rSw3
F9SHrN/gmI36ZIeeVq+vvty9FRw2Y+3ElINS0/LfMvnsdns+EwVfJftNO2Sq0QCseEW1tau3yfvb
y1d/aO7hi0Zxd5NUrQlWvyFIAEQxKUiJEgHN4nnYbQsuAsOkBp7LBx0ZzRXjYEN2us1XyDXFBarw
rMGi07HFTCAeXyAe1sjKe98vFz/gBlQmbZptTUyfY/WXBAj/Y3OU49ZZdyXAixn5hLAo98oFmNM+
Z+uDdPInkWYm0AaXHj7ZEN6fR+ijGjsO1vM8P4JN1C5rXyZreI3gcpw+7+P8w1utRALFtCyUhrgH
r6mcoJbbrBqKRP/eI6gRMDWR+0SGrRHonuz4R51Q7klPASzJsp6ndoRt5u2LKgHesLhLkY2j4TwT
ZEaWxZVFs+2uH+NUvwRBhOdtN3+liZmYaWXlHZ9ZZXXb274a5jvOEZbpJSEPqXnzB76Zz5qvPWXM
7EzEM2yON2mXGPcxxINh/LrfgaWUrWnjVaieyJmETRG5FWquxaWsTNdoHK9XUVE1dXS6TJYDEDo7
7McMAm3oS+xuUj7QOTTBXpxe2AYXCDNN3f4UQ+Ovav2VbzPqAADactxD3lF8jGaI3e+bywhL3+u+
a45x4gbxkHFgnjyxK59g4r7mviiFeLkURy2OhWGkXdgqyS3XK9Mj7BGSR5eUzKaOCW7mQrTKPFcs
MLYWLowjubnkDHv1R0zKmDkj32S8T37GwkT1ECFvWNggulHuMTYpp+/fsyM0/12CGzTZPMIvC+cs
E919kxT3216HvFgCk2eLpsbo+z9gykRDR+DIrS+SJzXbxyKS2OrDkYSvf405/FSoLtii+xO1GFpQ
xMMNDxfDwxpsShTcivdC0r0BXUP0jVfKHjtHa1KfyH+sgjWafnvs7QcU5RIPRkG4wvbr0WSrYW03
Dd7GwRfK9+H8O1A4FE7eXywFoPkuliQnpWuT9VquN1pkr8o9yDGsxPrGuNq2Bjs4B35ZpPBrVOhL
A6KPe9ASbTG/ka6rMEutcfuzegqCQKIGap3ZgnPeAeTurHhZmRuw9RhRygSnF+ghKcm+QI/LqglS
Zu1067UQ0APIuxwpEgtvZsjvzYlwjelKf7d4Y6BWJb6tlJQZZGNfs4ktnr4C2enBjtDFCP16SqrH
4gbG4otuRQhZfkBA43YO4KM+5VBOZ7YJyhXX0UlQfKqjbfAlhiuAanB/nAnvoCoO5u7IDvKocovm
MlVfIk9vIWPMmdQt/imM+GTqUjctNC1YtI00E/cDD90/y5K6GAMyMzXbi3ypxkfCgKY3lNID9RqU
k1G4K4PCiMAIkA2XfdwfQeP7RHM0aTnSrKbLo11U++giYWNH8+SCpu8j639FCQH6wfgzMASXAzhy
lMAPrcvBtH0ahj99E6I41cXHu11dprEDSH/TT531LQcvJoe1t6vLRtTUDv00jiNadjW94xv3kreY
UHsP+wTPDJLmY1G02EnTIoKxuaSoIOH9gK0Mneyc74IXf06WBE6tnfjAtxNCnzWmeWDljX655Bj3
jeHuqm+s4PGzzIL9ad7xII/mBjVr5HssZfuxFgRKZQ3jnqn0FAtawj9yUXm5G2cFsu3xp3B5cCp1
81tUj2Z2SVPn00beDYG6Q/KixoYdDjqzi9fLATD68htbRu9ak6y/RkH1qbudM1HCB6trpVKIVfUA
hHajdo2nVkR+EsfJ2dLY3zYZDki2pX0Hqhkv1FWfIQ3AO6VLxprz8YiDvJ+MhRlBIeCkUGWNzm5J
nHhEjm/gd4QeDalJf3pJWUhWedhLKs2tLTwkOltDwo+Xsfm7/ogQdq6RSmh9wW96Kg6q1CLuXj39
quLmi79tAhOmUS5wlbcGzV7zIewdgcpqhZTmmgMmXI1OY9mxLeDotHbquPGYVXLhWgGUDKPQD1D3
VeXEuuDy2At+AUcdiHPhOLnpFDpKSxkZ/sXWjeISTccVLhJ9v8JlLN0VQBSfTv+TdgbP+JjIJ1zV
NaYOUPJYP1ZGBOFBn4ChY+NIyGfinTAEZPsatRpb2vKZCd1sfQcscooIprqTOcPewpzGEjLxRhE9
dB1dtHP2izVLHmvXAWNGxTAT6ivCY865obnhb29ybp/ds8xwWtBc3iCJWe9B4EQPs9nP6LBCrbur
SUtrLD26WOF/6wam+IHDSt0rx78L6q3EHOAOYfJRKyCPbZRrAbFfJ94PbIKpTx4LlBHNjvWbL0Xf
69EmQ1fpe+Gbivh8JmU3I7kH0jly/0cds77ur4MwasV2GyKh5AUKbSYZEWukUyvtD5q7DyR79A71
HmBh+YJifgoRIWDGN9hCf/rlwzJmAymM6SSOBYlzbAU3+Ojfy3vvZshFhHTPMDzeXtrF3oi5lpGm
9TIA/dfFWjHVCwnp4abk1ffxLuAqXDw+c+Ix57er/ujLIsBgUcOAlpoOWkfrVC6WAZ0Lftj7GFCh
r6ee47JenSMWK38Ky81AbjdASgxGpc/84nhmN+BqZ8Tu+hTfe7MnUB9O1awhqheceNCsWV0dKbty
4RSum0YNr2nQ14/vHKTAEj2wkEKqxxyb9qmAI8bROPmqZPFpRLA9+L5wU+EtLufGTucSnORkyLUA
Ir88KjZfh5R4AWdIUhAD9D7cLz0HKcF2wB8m+R4SniaW7X6/luqPBDtgVASPb8XZOigID0x1PJTC
WgzIuugtgodQkQT3608j8pywi6dS2LHImngkk3atQ/azzaO55yagidF16JKPYBmb77qP4ReD9PfD
l7sMMUWWrJQAUog6OWjJuEyoZLmM0DDgxchwKUAsW1mMyYiTYidtYtBzfWGW2nQUTTJjUSaccrEc
HJBzT5xH/CQcGAM2PNkU2dDA+kr/qNXMSmSD2bB3iiMWz1+UwUslYccy2vmRQvhpkGf+mq1yqRzN
WmUk1vccoiSpKvC0/sESSc5paukI2RL3vGKW+Husm08XCfrpE02EVLF7W+/aLyP5YflNLRtNDLCk
cg4wzAr7vIR/CA9uNZ8Ir1d98EDK7K/LFjo8pIeBLAtGI6pFio9S6MW2ykE1TRDh0ej+K1c4chlU
HzgfflrYgLaDHfcXjoBDE0OQbtxdRPs5j/Dr7zVD73fkVq21iuHNMCzewiEZ2pkxc/GOcl2erWU1
vQ+Q2pJJuDuU/sWSvExPRkgE2oTP7Id7IUIvgYBgzvE6NLbk/2l14Slpyje8erozHrFzulGCBeQr
OJULH7kAS5ZjCLrHrbHZE0c4epB3f3A/eTsZuKUK/FqllBxaJcoQ92OCu2BuK6KUykeIMg6Q48EA
nEWZjoarSvlg20aPvKdxkToban369fgSXM/cOEyhozeifkGeEt0LdU8i0m61A0de8ulhQEjIHVVa
bpF/02bhJCZmCmFTylqVR3aIMiqiTiLkiFqM1cxZQPZTClKTG4utsjenieYQVOecvvaX3leEB+Ny
AslmnOC5yC0yCGQ6L8f1RF9NxG8vk1hpqfQfBcLrIqJjPi8yRMRZZJCYSJwuCXdA5kAYOgvO1CeD
GzNQzytt/CVhqJerNMVasoM0MTlDyMhuqLv7AexZJbOynXcS3vJXueJdCliNOZUMYZiA33KBK7iQ
dozSJH9ZochQZQ9vLQnR6A1kH96I5wYUNoq+ULLkZxwjaR8t9vrL0QRhzweriW+iGO4iXWpxnwaP
TZAmiDlLhn/et+e75EBrJHs1q2xUYekHKN6lvVpzFQmZO0VoN51KpgCuKKvD7t74qewiibwBgHD8
ydvmKsrpRE4p311jldH2kzidyCHwA3pkLmlC472mvCTJJblxgV/96/Z9pSP34oK7rMamlMODvku1
hRxHFVefPvACQ0T+Ao7tIWrGogHB4xlWTRDNHbHI4wBhaG+pDfeTTwC7kSjIpjW6kQFAWwTSc8Pl
/xQakI2LOX6FitpGUx2v3J0gUx0NUFTiIuI/n79qiKv8LP6CtZl/d3jNbTUqaWj7HuorXMSCo34D
qea2PMFNjHvW3/tkyjzVV4EhNKAEeb/ORHIwQXZlJESFQCv8WzR+y9ZOR7M/GV2C9wJLP3LBVslV
vhQgcYxWlnuTtnD/0UmL2KJfmyrfm0tHQxEntvezPi/2uHGG2JK/F8VMs4D2wVmcFpNQMy81g/h+
Coh+riyk3z5ns/WZzon7q3tdr+46J/CROtzIDWlrXy9Vsr+UuERC87jZ59LMHf9TBzU/Zi6FX8Lk
mJQqpl/VMPEO8GNERakF+oM3Tp5AtJFlOn8hzIa5mOVF21o4oIK41qhzBAlcmIiI0H/nxpAZ7i+b
xiSMuP9TXPh8xN8K1MoB+2kA0/YRV+fSHYAkd6S/le1z2BXvGT8TiuuMeq1HTm43tok2rj44WFEY
osOA0BlCM+urWHONF/Plz/I8AUcrokqsPTrZYBEs0SDgLTxblSWZ1CjBqIl4mBm/7ag6uz1T3C00
ApRIlsFvhWfezKI3C19LmEhjSC+FbKdE+uQZ67ZYGVwMl1WVf9O2KkJ9a02ELZe52TrcaqCqLfqZ
6op8tiq1QeFg3jrbGWV9oR4i/2ksbuC9VWkjNOS7xf1BHNXAuzhmbJ9S66jarVlRybzfKKwcAdHF
2eLvL44Bk5jQLe0/6rZscMUhFVrqLjjjvf/66+JAxzFrdT2SSiypyYbdQFY/MmqMhKuxceCT4pUy
nPsRQq4WUkLxKkr7DAdPRGDFBnqvKbCPzbTfloMTtJSUkvCer+zm1qziqL1RSQoGt+e2pwaRwb/3
4rk+f2LEfHoEIJW0Ku/2Boh4nCXhUgJCVeC1fSK9SCeZaZOohEuKiYvKFnXTe7BdSDHq7q4rJMH+
mHOiBa3ZF0CNxBfksuTPTWpGizuLtoZA6qh+d6g5Grr2aHMUO/OlLETKWrnwoPB9v6F57KbREPYw
4jN7ZDuRQyTiHSO0aon5PdOIpVr5obTgrrh9ZmxVG2VpNFeSGYuOCLdlX4EMO0HOQe4uNGiAsAFF
jizDvwcSXRhf5GibwiMYnqOyt2fvecFm4nGX724pggQNRsWCypadpYBdGYdQmZRibhGPAGSWHMve
Ak+HVjIEM50VNM1J9UG2s3Smm24A2w+Aq2tcF4PcIaozn7YGQ2Vpaye2d12+F5FMAr2pRJP2Eu4w
b80M9u8RxABd/mIYRlh7MPxBZppi43+GWKW2iMPyN38QsTylY+8qg0Pq8JEc1qfro2x1cMH65cTo
UM0TWZiCWiDnV2auaBBwNMR1mVEHpRlQgw39mhtXYq6K98Ms9Ah4Ui1lFB64F6kAOp9VMK5Kojhx
dyKhZoq2Rb3CWg0mtwh5h4GdnwpFfSx9yUeQWWt1B2SvWFUfoV1AwCAmSrT1Pg/dY0qSh+fbNEp4
2UvrHEhsTPyBCk542f/ma9x69puHPvdXltU1UZoldLIPPhiQ311Cg3z0vgfyP1KG+J12LCWwSI8u
ZO6I5kfXuw0bcFixvAxDSxCZ9zFtfw4+/MAEE4luFPB202ScXOhtgP2WJBXSgvlatVsKlPhMjiKU
6+PBCipUD+jjkwU7vworRBEBzmiTz+uAMoqBXP9cDR6EzEnimLIZLpQI+n7q43bGuBQcjvHKVUlQ
Qm0lOc44vfMRYvIQTaYSRK0RUzH0Ab/45qtb0mKJ7uaLQvp5NMTeWtCnJoF3byJnBu3gjE/Ke+0U
Ns6BM7xw0OHBvUy+AiRq2Qr7alakxZWxNS8oF0zRTVgYdO2dQpP1F/aoZA96pk97wyBhuupB8VDn
XVek2sKdSFf+fPgI2QP2cZY/EllEuysvXcrfvKgB6KtE45Jn59XfOkk8CupzHlR4OPDuqNpuTMeK
gFVAB/vPgq+aLGIaJ5WDLjfKJl61Dbm0G24kXHxoFGgj5BwpRK//qkmrQTjb7k/u/LEPwCeDfCPz
3JneSSDE0LrnfXrhOg0zEvZ7A0kUqtLj6qq6u+Lbs6l/iNKj8O51Q5L02gnApvwniNuGnEwrqwqS
13+BKeSOBnzIGHirNeDMrMNgjjpR/c3z9k+dZgAdhrZKaKV6iWnp0NPx9Utg2PPWGsQ8NT81+g17
A+avwPYIC6c92bdERRja8VIM2Jf2n3NKiKe0ElvqlM+BJXiKvvaIr1PxvnCM4SGhqYDSNY2Pb8V+
HsNam08W/P3gEEw+pKwyB479Ev6TxyAtCeMbSDNygRy8jkHtjQR5FmO4Mfo4PIELPDmEfqKNyUDD
FXMZZCPs/EecwOLu3qHLnUP/ap9kzCYcU6Khoys0gBMHGh4Jyab8x9VHtFaEvtcrp0gw4K+vJF1g
lglls1dAhTyZOJv1KHIJLjyaL+vOogvUOqTe+GSR+8nfw+eYJPuohYWasyfgjLPRcOWb2SAYLA9I
KXKDTkNZEg2/ZWbuGnGjWw3gcurUgnw4cPDKrGy76iL7GANV1r20cejpn/jGlv7TtsJ+tNlTUuPR
/oXRzuXsY9uVLOzYSmW2wELkLBoAVhEVPl24F1JfLB9jW6JDN3Sw6oXZu61KglyWzzq1MQ7uBOrJ
FcWzP/Wbu5blxQ9owUhcvctx3sYJN2Q/UWasrAg2AjROuGzQTW0P7+eFfROSv6CiPf60tyyiFc65
8btGuuese/ueMdc/w+V5CVRP5oo7VocU5lYSDmGBan9YQA99JvWhft0gDROCvUojxrSVhLWXNy0B
dn0r4DO3581plCYMwj9/v+AZJ84F0sA7oQ7L0cyLFbBltCO2tvl1d4+yp7H/KVu+tGvaQ/LE4dZu
aGZlevEQbPVRtQVF+NbgdAZkbnw4l9IhKfBW5flhAlUDDUDJUQI6ewZAbWSBn/aNdocpK3KGTTM4
slJ1OlUWr8Dorsk6LJqEtDP8uI1gaemr3gaMyvLMWR1xH6GhbZv+1w6OtoUC0cg8AnXqWsyz7JCA
rPikbrnKdHNSMupjY+ys5iDpIowHc8ps16Clv59L3camD4bLPO0enFYG0PuHyZrm8nMZHz2cDn/D
NEw+w3P0X1yVOX8HP8y6LPNrSEcRygIqTRfQCtR4CmQnl4uG1DByYpzvfptBX2RqOM9ZNp0GNKOZ
gxEDNjF2mcZHlAFSjnj5yCfUOBlqucMVTOC4e5/nnqP9ssZjBX6d9tbVYohsaMqw/EBL05NEujF3
APxriPQepDIMpUWJ1ynwlnB4ZpulWVPILR3yp4hJs+Ns4OiDTUfcMc1sV0eQCFJG4hU+FoS1Znk0
2qOY4d1YyPoxliZfHIRzuuXBPbx6rYLeKGaq6Qkea6+MnCYsWGYnMC+t5okItVTZc1sFlG+uoRXw
aP7PB3o3KdZZnMYW2ptJEAZJjfuxiyg6nAu3YLd4+sFtzg0jo7QkviTHM0xgcRF85Nkp0mm4rELi
cEusnXC7bNm844AOGeeUeQABzW5f0W6EeL/gURuorfVQyeX0dpgh3JBxlakGR9MsWA1oElG6n7LZ
FJZagfs83liLgs2NTaCAkV99ndtCks8/ZQC1gVhoVMlSTUDvATaYMYnVlnPpXPiq5zFn6LjqOiMa
ZFFUGPo61+gmQisexnSeNO42QxRzG1onQ07f6Tx57Nma/CwqifaQI+lrfw/ktQFLmJDhaEx2ZUF/
Lpx3cb9uONLZAai4Zdt09/4urEl8nEMijaevFCBMuQWNWt71EL5Y4K2E8jGPxSpyV6am95BU5361
2sd0ZZpkbNb+9TMlVZ1QPbLvycVG2uj5q73d774PRIjAB/v1kVIMSTu11qee9GN6JucRYwX1lwHo
ft8iOG2BXuWKRuSUauzIYsgnhRudiBp6/Jy5kx9AL31OgWu1GqHWJfJqoXpQOMzohUNH0YiwSjjw
yH6Reqb9hVBS87dT+daEG6N9Dj5KWyuheNDJbKed3LeqwM8GStLNpa4eRSO2xYPROjKqtRv074y7
9zRuHLX5ZxztPzld/iAoEbcaqjVN92Fgmqj+H2wrLgB/B9chelcMPgsJBVzd9H1FnBHRuCt9ojJZ
9txqIkxY+g8EcB9CHdnrK7Icsg7RktRfuJ3Bv9vpwUPOO2lpsEAzOgouE2DL7gPtWfL2gWmGaO4S
VLMUvx4LgDv1OmUGZfTjF0NbywtDmS7m4euhQu3O+/5/ShXMchkfCVFQufFURl/MRh0XxFCVsGu8
d/gZJiAi7M8UmRh7Wa2uCGTtIEwLHKSMTmRfoN9JPZxLFmpZdE11GbZFpn7zEDdG/qaTUKXM/+Qa
f4FwROKfHEzZAiCzri3577cLPoZwwPhpC2uHO5Z4m4XvNq9KOBmUx28+E9FCdYla8CI9Jxyi0qM0
qurdelo9Fe8OCzx5YsEhekqVDc96/jqXPKEd0295REvEViz7LZHR8yOQuibtfTkV8HxTRl4dxKz2
x3sA7TtfrS7fdHwDLNU00katmZxg4CUof39e7I5krQXDnFOzpi20EqQ6hDbzVZOdn9eAaMbpaY6y
SsoPtEz3jkpZ8ppexZQubAIcorg486+vRqWFJhfLq7eISUEBVPFKm1KH+5dGFadHLmjbwZjeBCg3
DYBrDIiynYhTMXxH5e1c/2HXb48CaGYZNboZsfamZi80aVVnayQBPkH3XT6dmMEAWrLP1Yde7HBG
PwyNVJhVMf7LFdytht7esFyN1p4lhUX4GPrWYcsUGZj1brjzNO8inoWhMwFFMG8G0sfW2iAinjdD
DReMmfCQ+UxWxokJcwnFgd6gDFXvCtgYaubhmq3c193yi7PTlZDOxMzjtygBeLa7XLBcrxFnIJEe
d4jOVS3yZdUVDb648RfAZKM5MJd14r0kx5AzwVuYzzNtSyEP76HaSbJwKiR0gTfZxGfXjxoTirTT
LsE1Cyad0tAYf5pjK2RIwjdm/Da9/7zX+IfNZGTduOB/Ze7QQUJEzBU7W6r+GIsxR2sSZFvBNPk9
egHG7lmW/NxLUU9KS40F0XScIHVhZOf6X7TMLUv9d5sh2DBffF08E7zLw57qDB/OLt4M//26gFc8
sTE37YAidOHcWmJ6PuE4UzCHm22EIevvzVouxFCNbxduGXExH2+ALFWz44NrAoI12yt6dUlK6/Il
V/qw8MFgj1sAb55bK/D7+ULYULEcVRMWw2lp/BS332aLsRjzbqbbEMscqRuIYWId6PgxKf8oRIhi
cifCk0QirnhUfaPzy4Ajaj9kxfgs7toVBrxyceI+B1Uk+5ql9YKAbhuQGctOhmClD6hz0+2U//I5
uzRBO7xX+VneQ2kCxKZpbJUQcaKGd9cyh46ayCupYpe5MhrqNQ1lE+XHRDGpll1ehjUfhrhC0M6Y
94dxNnxGQiMOrRucMuz2J7ChtVF45lZjq9flFaNwJ0P/3zsbiBgNRpEqQ58JdPVOtr3B1h5+AZcI
cADOAzVaBidTHwsTy8s/PiRN5KJoNAXzsGlEnAueGbC2Tmp9mYurb0za41VzZyStH/0rtvGt9xKf
yU2FulIeFP0NFinZM3qteNLhbrGqBmYc43Nb4Zvg9mi6BbLuqRW/t8klV9pQZim+WP+MLUz9EcAR
uTx/95B9+mrwWe5frl2vIxaPJL/3gz4/nvmhbf3yi9OVKPsX/BBLXzHebz+wdJRBVlpBWOaYaq3V
cy/G3byQ7bQth6pXj4WUHgu7Knsy2B9h0DZajZLwAgPN83ZDUtv/adc+mkJ/hvzEc+aLJcVLI3Vl
R2+Ty2LGuutNFujsiyqOEGT7c1ZExUdwTZjoGrdkRo4hMS4EbMURbGojP6SIgfn+n3RTmJrJg1oe
gWz2KZxXf9LG7nBXfb9Hg1yKNxgF34KXWCjNx9Rj9TUnaGgx3/v77xTnbIfmpcNIkqvGnuyb4v/i
K2+i/DOamY+83/ER3+podDaxHrvT5aWN/4wWhPlMs6QMtboAIxftwRhofP5YH4/6fQeblxO59EbC
0CuYBUqm36k+E34RKl7cMM3dCYoLXOARTQE487byAeEKpk38RPTSvOLzyd8flpGfJciWgQHWOGFP
P+/TRdz8uIwjOv88P9XyhrMQEyklExiws0OgKL4sAMrN9+X+65punq3GzuaBLh2eT7X6lZHX6wQJ
EMBtnSV3OaLoIO7p9LoBg4TmmZbGsl/ClgxRHkOA++DztDj863aIVXU3vWgdF/WfoIqxpY2KRhZu
/FC2zRSzvRuwtPt+1Ze7wT6D12Smb0v5IiGLaHf9F/ijzXpEQSbMbzl8J5CV/WokXF3D7sjpMf54
pkV5sTRtHwqX5z3fSUXWxUOKvBcZPcX2ZI2V4DC4fYUF0SQHlBiN7esjls3eFHudp339KlSIBPgx
giuLi4/7GLVQhJveOz66QRW8dA6SoXd7NkWx/iIiBYpte0DSTUAB5MH5RMvvZFfdXTgdmG+MDQKk
ISEwyyl1K0avIWZM+HbSp77qngYkWT/T0W466exL9Sv2E7S2sbl/8R+HtbGnBNp7wXMbY8z2G7K4
G/NwdApPRsgnzyxCj/H2GDtzRO7dhRkv0Be4Vj+WXxNVZueaeOYk9ZZgcFoJmIwrWyZOTOZ2NmaU
oUMQY0NbQsY/V4gRGSzdImBk4vpAQxEDBkr/LW/ChL2cTB/PZQY2SlrC4ivillfQ/Eo4YAbyA1g2
8bpYdcJarVFSX52ggONKaIG3KqYC9sLdqxH82uIyKp1LqJI9V5ajsPHCWf6gHaKJhUumIjnJET/q
urIOtJofF1MQpkM1cKC1yNLLVlC9CM2FaCGsaPz7l1O6faGUrVtaxtbnrhizKrG1C2AWIKFcSt3w
Sorew7i6vAfJH78XEcSl2DWfu5BIvyNdz6zNdPTLXHODMhewvxWPXMavS+QW813jupvMKOT6U7F9
n91ofNQl84RDpLv/M+j08zRwvk5Lp183XfsfHnHycN4CJAzr9ASTyWqS0XWW/USfHMrFQXyLSV3I
uCNFI20vBuSOefkXqz32eCKVHm1IkX2afN3YqCS3xCYlQ0Mdv9Hunbj7JF8g3bmRFys3iVRunkE5
cPnXs9IpD6xLm9ab3yk7aPz+xprGNve1g/kEFzxvEFPzp28gpyJcbBE9PRzv1S0dEk6LHc0y14qm
0GhQ0qZ53NKZSDgoxL+HIpvoWVdkZapy5im1IsGW8pYwfSnZOhZml+Kj4rHwAtqXzJsz00lx4wQ7
cJM48hObwm+CUuw1byCfmYPx+5U0nrqsn8S79gNUByFW8to4EqtQ1EdIczZY8NeU3xyNgVDJsRx+
5Bo5HKBf6rH9t06YWoN9/V2rLNVrnzlzo6EKOGPNddCpTfOURyFj32b8mK6/ghko+bBlzBR8b82+
5/IE9+/hM3DZHPG1I69zzndGYRIV8GfKk7kl3FdKeJ0TBEsZVgQGLZg1Cyjh/CeelX/CrVywN7np
xe2kNQJDdr5yot9g9TkvQ2KQcUmFojc9HYu8vbnKHbhTtKngS+TVox/vB1mldxpgx4CkffbdX7uL
nj8fsB63vO8TfqEFy0LpXVteOoV0WgGDIdV0Sd2KsgTnEASXhe0Z8Jary16nwhxqnAOPM+lMki6j
65N5X2qq8vGwsCgvNh29+r8plyX81zUc1EFxlMih/cvzD0hmXhbLT3mc7AVRhbROOEArENRy/4H6
tDktbrTm4X5Q8sd4H0+2R+wBfBfzPZQtSmQe7jT7gXIHA99NpFGpKQDjH7WhTvAI1erl8iJBeINs
pcO9JQpjcrModdqYVm0ekNUQEHIWr9QQIQ0yCcuMOwAdPbOtfLWiOnBOgFDDWKP2x18sTwqX+D3F
1EDO6Dl/t7ea+9zkT8qE5fYS/pTqMo445PRPMUBpXN7goWMVIaYEjoR2FdW/O1sNPZbDvPuQj9lb
Xpw0pYhd++VkdwYTBsm3SX1/yDR0n5uO8PArNlDlwr70+u+BKmaL9xLO/J4C8UeqjKSdmXKncmat
w04JdzGoKFbWkVZQiEQSOJTKKEa7smZsz46Tr96hiDKmpxAMaJJ8i88uY5FrlowYhlHKOlioO31K
Acu1tGjkWP1hzdH1l+UlEsiN31Qo9yxtxDb7Y4wKzZmFeg7/n5e1jptuaorE0SIp9RAWwVFVnZvX
NTEL2pWzuRkAi37f/WDh1JnZ6bloL6ptqtxOZYdzGtHJaenifH2BGYE98U+p+8oD765X+oq/hGJW
/YfBzLDz1WX8Bl35kwcuia/lfn9jW8+Oho7wrHkNWdNDKidyEjGO4dspsjKc2uEZDA1+En860lfy
utpMLTA/ogbqEnR/0yhxoh+cGXccA/NAXS14XpMc9SrviUcmGyRLXWJt9hVy3LZ9ovkxZUwGv9hi
BsQiHc7WQBF+1Wl4sPBJKAgA3hvGzQCKFRDiyiJyERO3aLXV0iA8qcMUyFftoT12l3ngb6lOr6PK
Rm5bjhDUsS2tKMVnzy62wI1EiswP9YHToHejQFRHg6plhSwYTk6IMa221AMyDlKqJQPNQNGte9js
btFOmHhFRrRzveafcSUP4Puv9F20ND03NP4CAZtSnGni328pA4krbSzdlWLhV3yMM/ZRrwmtFbDb
u80dsZA4/+yQPvf2zPB0h6MV0dvB0b+6LHy6xRKgllCpELADb0QDc79CkphBR/as/LZwyiRuzpEK
qB8fAdmTHL1SYODzpHxTwO6LFP7HbO8EPj1vuXJjFRTAbWo7EMVWNPnnJ+k+BzirG2Lj+0Dkbb1y
zwIPA85Wxuphf5A2DML505Q/mFRggypYtTIIWG5kgy/HO4VsZVZ+7tem9jTlVab+Y+WoPy7j8Qkp
B4rTKB8zNBOXEPtN44A8aS8SY5LSJdAydWXlduVO9apgHEbvyeezrx/GP2J24bYaE07/252fA228
cHKPjy/Rp625984nmKM42tglCJ7dZ5ChzgaNudPCDgeuUnJKNkxNUMwLGvAq4tVgqnBL24O4LiQn
BtD6eIRFjMXp6CSDXzJzE2Eg18M8dvPJLriaxrZETxajyYBh0v8uh9geTHrT793DJyU42HF5zcT5
QoI+XtxyKHggaLsdHQVEbSBLix869VXnamq2AL1pKeXMGSfPkE/TMQKvFpYJpSq73xZncym/WUT1
utM1oiaXjN1iNaQoHrCXSqfV03tf3k30U2F0bIW1vFoexsPyPv+4C4M3M1f88azwNT0B8YmQikGe
9G3oPEpEIsZHZuksuqTgyrs2QoGZXQwLWl3zB6p7fRktWajRdw1TgZy26Sq8cGfGA4A8wgctjr1I
FBtT+V7Y1Rw2XVKUZ5KghdW16o7xU43xYbk22EqhwQCYgTaxB55H7d5h34/NJzCX6wReM9dt2L3c
pK44ucYtHOnMYRiZsA6n0LCuLOratjYWh3l56Uj8rhcjvkaXbJrFrArAdKEzSJGnFUEpQOKUQt6a
c0h8qdddB9oRWoxTskutWP0eGDXKmNmFZs3OP3C89sCRZVEhSRP2JUNnWcYXvbEM0BgRSn9RhhRM
loVqEyWbVvGcqWsnjXfubGEzSmqW9wPoB0Z/bg2wkBjtRwY5hLyZIXQOc2c+UJXn95ifigUaZsHF
s+xPUCCwvuLcd/MMKHK1+F9iO3wZA49GvvjbCV9GbDz+TJUhlApVNJdDKK7bTYT26j32++fohZPj
98pVtRcoNXow0lQUkBFAjGq9w1dSDKo0zt3QKTWguc3m+bjIR6HCQw90++8MUxSaSqpiQLay8loH
64Wr1rdkpsbOHosYkW7fQRpx8W409F87LQudMkS3DQyi3IgwnjGKF/oCZskLyCx/MOFug2arjHhO
aygWZqie84oiTdHX4t3R14BAZn6iI1yMmmPsF+OkU0UyKsPbWwuP8aKvtq8wM23O0RNMw/JG9yw7
LSXcjJd++h3zibpKXWUE30AzJMXKzVMtSxhbKD6uoV0HpP0BpHXYcIJehl/9no0eGtXsrSKIsPpO
fKThCPSWlHQwuJVoKiW03ruQeGDLKDBAON2JhkgOsD6+nnwGIQFFUYCISqyIxciBR4xKre/OCL2/
HTTvAZukJWpktHTBXYn+xM0ZE7+4HdlAG0s7Wz+OmZLXDum5Kk5Z5RCQOjzUXnR35kBuEl8ADJTU
HBKciak0Ii7CgvZy2iHr8zOgY1zfyV7Bqe8iZWL7cheZKchiIJQ7nkF6voHb5SLfKNyF1jcHainy
fghiqiSzDp69I3qAzwhlWpM1DOYJ6eCfm5PF9KJ3GaMoL9Z1DzH1mkcT48MfT05fHfJ5pr72m9Si
GRUuSWND1LAieHewAYzuUNmBcEo3lOgBRS2LN/obOYptqDcudqo+TRcKJN4NIInmko2QYZ//80Yu
wPBhNnGh4OFLVsPy9FxDC80O2lOGv0ggC3PXD1tI/46hp5/2W8/wVj4OJzDPBrIYFb/Tm/faSa9v
MkWxz4Qd8E26dYsUZjLA3or/gCSWqJRP03SxB70u5ZTYAEe2HKLS84Cpw2SFlHJVLyOOopF4oOh+
a9rDUN2ZH8gv8B81GluUVwVYllNrixeFZiW3WY1uur7qdPRQF61MUAaOGdi3WR1tJT9JtT+3g6tD
5Y2u/7ueifmx/gbZ8G4u+A72f2DQoB9kkrbRpgULXmR+WfVeMYsybqhEF58Szdrv5ZSvdeREBpuS
qT2OvXIrmlXhQ/VM1sStrQKjGdEF4AdGDJMF9XhmejCIGITrbcXnzIyLaX70425kpX9dB81i8Za5
QoEf53Lhk0slLW5ctiyvnihlvK9PKcX0sntqWu3z5Y000+LOA0uc0QslIs6NHFcW5ltDsRP3Xp7S
v7icPEkHuCU0IGqcXFiJVt9WzSL0bJtrxSUGMX1CMMp7KkzHeoqzz+/596tzRl2Os8NIwXCmxsto
UCf2cw8n9l+vRBtLO46mbRJx/jecKFxpJPblYMddPiOnrcvS59r+HHp4n3fxkC63Zm1M0i8Vhb0v
gG5hrjpsWMfVlrQYjdEdeKk6nQqCqeTtxuJB8XC2VWEvW1GnL1I6Ecps3U0Y/FrvMswhdO2+UJNe
b36Ky0zqddyeDUTGnIpxNKnRNIuaeU4bimtYBTfPFy5cXF9tnCQhGay6zQYArOiB/N/8zpgsx+Dc
u6Iaz8Rexen0cUWG7ABhQDMU7ZZ8cXhoC6+68yrJ0kjzMqpyM9RtClCKdRXhytQSHi4hT+an3aqt
ZvO5bje9uWxQlf4natv94KMpMgL+8IjCQCdc0YMfbMpKpFd7cJNhgB9CEjLEwxJsd41LTtKeyxBY
nng0mx5NI5LvUqQuGJ971Ps702PTcog9vdkMbLpdHG/NURN+IzhVD2G9ouJ7AZkD7MHRUCmYuc6V
OFGwVs3+bQX9vc9OrisM+ZV/AftG5AJcb8yLXbG62tAxq6+k3wBs3OPPN5EkHYaJhpcgQTFdHisZ
Qk7+lDI+SY2ORQkzKMNZvQmtAffKU5YDZ5IRIwPrAXO230Z5xzLTKRSUiO740i2d2VGBSgcMaNNX
M8Eok1RRcxoiom/qI5KiH5eMWiuZ+xPHUn93ySIlQMNoVtkZL7LooFfEUtAzzrbJhXQJzXHY6TAu
RVl/vdzFm/340f7P8eUbgbsScyWbke5unzHnOb5KkJ5R73kjtQFDAPhOgfkpPk6FX7Z6UwY521Jf
s9dO68qPL/D5bWnu3yMgQFDt8rKSIQEJnmIlzav/InRPJYru5iHC9n+uR2O9w5ZhpSgkwU1BSe5J
jTkU3Z0cNx0b9yeECtBXri7fiC7vnL4W2V3ZUF8hj1rH5R0qCY81mxQjptqDk3xCkhaT+wan7wUF
9dhZBy2Ij52lv2ZK9Zw3SvKpMOJDSx3Lxxu6lDPZETdloAswJXcljvdKs97jl6MawGgNnbS1V5kj
7oYRFnAsjBauANQKGxUQWMYgtBV2cq/NlVASd0QYp5OkB6flhAtrlBXjv7CNDcIOn+g8Q92xba4o
OQSEKftCtq7qnBliwrQu5YXie+QQKvIXqZC0iYjaFmqh1/SgCRR26tvYmitNsrkOPGsrq1MwnNcb
IYaK9lb6bCDA9RSSu/sKsI5mjlrnFio4yI4aM2bP2ARfpkRi6VgE9ipFv2ImFL5dAVM2PrTImtPP
VlYdDkEbXYJB59XPS4JifQjWbV8meLhpRjhxL1ncL7xtjwn9oOulYYcqWtCY7t3QgwqSRbFhEg7n
QZT69kAFjUysPflTlfVkeJrdxB3yF402nngBfJXOX8TD3Qnoyq18h5Na51opK9TGSBa2ZdXQGBH1
Ur13HqsxhRJnMglP/1flXKmFn4phRBzi1dlbQNSrJQwrlfbO34XC/e+iBFhYx13EPADPY3OOz4w4
eaMZfMTo6id5dBHY+0zA5QEvZPSm+BwSqIRhTaLsx8Us8kKLM5lsU4YCpTrhZlLe8jKik5nwTzXO
4DAmyqq3oGpKaAkEjveEdVvxR/BBjIdXSZC7RWc64SgjZB8jCYRwslXJ6oB99c5iV9hKRkJ37eSq
Q99gzIzZJgbMo4+ZAHuf31FcxfrJwKWssVpSa8Fz7quKVTBHlSwmNncF/0uAPiIOsvBOFTOycOOV
DNyz+Zl/TBDXv3JVjkPI9N9srgK0DZSEwzpHQv0kqlRQoBt9JRAsLs0YSeStJhp39yCqRHZSOaZh
Gcp/HYFfBNupQfpargqetUEDuepLuZ8f918mT6zGOtwxYJrPN3G0eIP8twxJ2S1IRcHxhb3YEbAE
5JLW1WpBdQ/IjNBdK6H6tRIXDx4Q3g0XlAonZI+tDPJJ6PGJAb4/hu8zVzKmkVq8JBB/uFSXAq5R
wvlEl31ye9xOka801QT/2mov/bmHv5bFWnfSx67so2pH+dBXM+zA2TPlfheZ/eTSQRUtq7q4t8Mz
pOMGE2i/3FL70pnb/1nuXf2l0txmQ1R//+5e9oYczESfS0fpH8gtBpeOBuaCDkwysAvtwwjoklND
A/3UA7szKp0gBPoAldl2Ej8geAKdywsocTZe/1HpuLNAbvGPfJT4aKgigpIjdYBnTdzEze9ucEPV
5htaIu1apuZdlKCWYqv7X1UhqesThq1nkxFFqinvS85PGoeJqp5+bEIg8pXkgwAg44g3laaXXR+C
Nm7JAiQDDLVyeE7nnMwlhza1q1x4YSLWhWX7mlLs/4JDyUeG+sIbE7YuomvKtUdIcGv4ctqYMqYw
WfumevXdBAUNSpLuk3DWIhV0PhTX35h5D6deyUmVKPlhSg0Imzjj+v9LdfOjlq720SUe4ENrTq5K
dZ0YRGiTjVGval0ZKE4buV05NDiHFmnUoJpWPo1odJfOyeXj3G8EFJGR/t7lbDkHXUbtmuwMJJ63
LFb0OmAibryl+/DlQVOXTie9MaEmNDLN9beQ4sQUR0+IeBw5uLErfVlxwXMLkJrzxdAKKR+lWz4I
q6eBbE9MAagBvSev3tGUK0Fyie/9ce++mXrNq4t3KSLfFck/05FIo57QzWCN6dnno3lOQs3h+a1Z
0j65bzBCwop9RUs6mGRI0yHIvzlY0n8zbpIOQH+xidnCsKzPjvH7kpOvJPWIKZ8KIJd4yckjRWU2
hAMJ/Y7+QwdGmuflzvx6uljtHg8GdfKlvMto5O+tYQYpo0//45WyfZCDq6UkJSJyCIrg849MMsLf
DKjM3eVGJ9Ar8ZALG+K40UrTNOjFUMlXZUn3Cd4ihwiX1ODuHjdDV8OMy2BBV43W+zBlufo5App2
vhkip3mMgwQH/lT5HxNizqr8uZ4T7ICJB0Cz0l6BbKFAH2a+PcCjnD4g1ovFVnQVvqfkZaqNWiV+
ZGNQWZkPogGTz4yLs9jACVVK/3NoEMzO6DbdI38dXHIyA24I9dIA4lYPDaOhHZ+Ug0fd0DsjrLRz
oRt7mf99oqQSzTO6Qc/Kjkmavw1k6kdejUgXyAW8iodMxUFGyTkigmUCGuCQrCZ1dys/iQZLNyhS
Is5FleAckT+/plQROPdH3CQBN69CzvM6nlaPzd7llh4IoUu9xD1fEU1MW3lQu/oNzj2XwpZ6cpCl
a8CtvbTRy0oyWykNHMVSszktPe7YCXRhMrnj339g9+JGrHZfOrRI8tTnyp2+2ihLlqR0DVRJUdyu
dzljblA6lGKpAi9FqIK81tJyQuVp8eMtAD7aA7xlQobZq0fINV2hGI1HYzodcc6gLZiOewqFGPcN
5LW8RndzvT0jH7ZDDPELbEqeBVoYldfYO87Id/7TAakSzwS9/46kqu3FDL1C3MH921lorrRnJlG7
d2FGrEPGY27WUBfKlja+F/sw13X0DqKHZENwsqWEfnV194Bebm/xXF8jRxx3lM2IZfD8aQIhG2Pg
DaUpiO1Oj3wsKxVz5PdErNu0tAOc9/74CvlrLqG+XMiA7I97xYBUakx6rp7KIbYFtf90pgVjSOQ3
MYbV4UnfbaQK5AQGiSiXXa3QPFP48f36mP+AvF43qKGHBR9cwsz6O1SQ1zOvNgsIhHthsMWp7Bhs
DXinTIwaHJKbiHoVtj6lBVLyjuebMC/xYXYqt0HtbLaVz6ZYBFFt+hCdqjm27Cishkxdq9uoLdUL
rXMYusGwL86JqNVa3tnwhfL0TXhy352Eu1tkUzEy7Og0+jzy13x0wjM+dfgkFWU1rMwTsZ2Doq58
MsKJFmoH+XlwOewqmfgZmZDH3ZAgbkkYpWBTV/5MdEwfq/p/PJmsyIg2NKGl5/TPfKgkHn93sux0
bkWKPcJek9cLBL67T62zGfFPSkmvLHpd7nmG2bXJK624FGUQPzXW3baOip0XxmqCmMwwPjSxp5w9
bmJ+AhhduX5RIwRPeTnY1Orqr90yjxqBylMo2WGJ/oxPEU3WXJq6qBsh9OY1uljlwkIx8jPg9z+U
+1OH21K5RM8AiRD4JYsiEG2MjNQjFTOffZQFNTFzNwk9SxAvhPhRbOxwCbY//fwtANImsRCuEf3l
H3+SH7Mdbh65xR1m8lfAdMgpKCqnBZoH9wdp3Se4EemWrM5Lhl8LhLK0yHODr8O/lfRne4u1ksM+
HNTQ/qn1mjlWnjkN4vXfmwrTjNfSwUlO20RMlSmj6SGijqxS5Rng+8Fs4iSQ5c6sNcNQGLz/sZil
rPsr/cZx8eD+cTiU4Xa1HZktkI12davpaS6b7YW7+28yT+bK96Z2Oj713p1MapvJ4SaolrmiZz6r
El/nmng987xz9m98lGUkevTzHhJUinMaK4PzjR6CE+PrmIlcD/SbwDO7acBHzEdrwrI2wypikX3d
Sr2pVhoojHw8zM/pmv7YZ2WJ5yaOrYCeqqArpxXdMTsKs/y8pMrOqTnIBIpRRi74kBS0P0H17+aB
5sLEOIx1BY2ESagccwzZ2N5GudTkNaXRnOKBjXB/IJKFxtzTqMnzRq+i1zpG6Z1lObgFcdpAdjlC
fDqJhbQmVq5hsQOelgTapMlm7YlcxxpgQuUT6B7c5x4F+2TyLgctUg/xVevjrBd4LqLRNSlR+gDv
Oe0+h1vc8HpAUPyZXbUmSsBLQB2GNZY6nBs6LKmtVT6vcfIDIiRRUMZzpx5LGGhf2EAjR+ncdIMV
ipd4kCJZPk127Vs3cDod0Bfs3wsz9ZivS1VLMhsv9EFe8wO5+c9Iy4YqG1efruCA8QauZWi+v3d9
SyLvwK+DDGlxIJ6frhXWtrmpXhf/HyLHvUV6oTnUFwV2wZuv90B4vre0jTxYd+9Du0/sOiAOK2Oa
x4AFM+OD1IOxPXTeip3e6EPdM5GS1ZhX8Uro+pQBp+Y6l4Ug7k4Z5jmueq3YuJic6lXjn8JGryXF
B4o5Z8N1l3oXrAs4rfZ9lQEghBTERA7vetYf/U1gUYyXPZsLcLhnTceOv0pc+gNkl4i4XTYSYIA2
T1/3fpkmLjVDpZg0w2jdFz5pRVDoUE/epav1lbiQDcW/nDAvFEtrU7m8HsBn+NUud1njGelhhIZw
i9P/J2Ry+OdfAHoklAVZqMx006nRzqOW+St8c7QGMdrx1eQmMZ9OpmICHYlNl1y78G4vpNGF20sY
02KIkTAPAAV3J0FFtaX1VMb/nveMJ12ItYMKxGtMpJt4lJ+1lDuHZ5khcsOn4jl3MbCXDAnEHxiL
u4Uj0HvvN/zQz9nl6xIpdZ0IC4gDiOp9OgBLRCoqqC1/xW2HdarOEnnGRvPFPQiE8ei1gZETuehA
uu8zg0Ap3uLANvsuhzGPy+WGY5ncRkDHG9uX81CiftvKnonO3PY5CjEI/k0Uwno/bl27SWwxyAcn
f9GzUJxz7ZuTLFWr2Jfsehq8Tr3kgvilcedL1P86qzJm27vZeP6LYs/uMgSLRv07sRMFJB8bEUFW
26oY6A2jzgy1JUTSAqpRZbo/eHNAnTcr3vac3m/4jq9ZCMrt8ojZ+Mocb5SMGhPyYoaEQnD123hf
OealFgvcp+AIexdl/5j5TVbc5EuBArCm/qlTykv1LcvGxk0Fwc79oJUjgBkvuabDsbfyaY9x/NJj
tgm8VZPnlYrwQO9kcu9da+u36p54opJXgjV/bXh1sg/J3I6NQJtpNNmIdhsu7CgR+cCdR+cSVnga
hqEUTcMNEml1n2ecqL5EoaEEJ6HxiLi+Z6YcKGsayRBBUDchRbW7ay0yb4i116Wu0TjMuPO1WJPB
Njwh/8bw0gu4ZoH2lBK1hmC4NekUlTfRI9ylPZDnAPq2JJOMOoeVWjseLu2QEwNjLYDibrdJHAOO
bo9d8ZHusaWRsA2OveF5frFKqE+s3QcwEjynqWhGV9E9Sw4p/nm+UJVV7pQxJKmN5XJhACKyfgPd
c7yMlauGaeT94fqZqHokuFazYnLQpuuM355zKVVeXscIzbdfb+NYw5eZfYZd1dGLhmko3mQi/Gl0
dg6CtgeoFPwMpmEXqcbh2UhUBfIQoUY3ZDi274CHYAii53ua3lWfHy1TDsG2DLYuNpniaXmObfKw
wDGqWq4YMkZy4klMcrC9BuwduDAXRhTEhrPPM0mc04ms0nfCUYKFLqSTqElK9nxVt0YA0yFJPSRT
hPgKLx4nPWy0v6EN4B1zlZ2p4X6u4gV9QFpBlhrbJe0oBmD+fg1XDMg5x5RWL9iCuDalmdaV5VhR
pbyJcGIcARKXu0M/A0Qq/M6zxpQr/G5E8pJbCKJgt5CuKqnowl+LsKzZYB1RpA1LCw/kUKrPMRxq
QGHe71vFIxDZR5LbJA0KhIIktFlpFo/Sf/an4Nu1KaXqMUz/hzDc9fyQAILzOcfo+h6finmvvNQ8
wfbnmdz0qcssC6vzCjzl0x3YiJktDJfxRuJGRED70i0Nau/edoHUXVkzS/C5YR5ewZeyTInJPwY7
0lAE9e8/IUl7dRx8gknWAWst+LcIsyOI7MFZGxkyNApAfE3NvdEFO7ob9IJ30c0sCdoN9dzUgnOn
Cys6MNurGhMYP54N18tXiGE0QkffY2jGpDm+agQvJLGRKphjp0wRY79wD/J/GaPW1h4ioJnriFwi
M61VvtQWMPxILUglt0sCrRiEvmA+X2uvgBH0vyZmyNGfF1LeAvkR3Jio4AJFg5Ym8weGjjEZNxGi
EnpB3gbSEzv2W46hLKcLNckILehe1Ic8QBtuxHfYRvqcUgH4cuCACjYAHTPURudVs9dbnY5oq25E
GXMclOFUVkXQyOJ6LkCpraR4awIHbroyFA+OXPxCTvTjDDzbQLv6lzDadPcl8KpKyKJqVOU6loeE
RxdCXsQ3gQY24iWYoeFqykwBkfSg9Z3GQG9oAusRplfxYXLULLjeouyIxXkI9PB4wFkbSSgJaakT
+rlrIYsvdmvAfOAFCoC8p29ac47RAkg1Qy28Omqr47yOURXN6qovsdkxrVTjsiPFlN4xYYkOpn6O
lOsUJYoBLRA6lpiTI2pCm7t5uRjoGqNNWEGA66BtqnJeCR0bV78cVsql9Cj+1k35vq1uBjYOGara
LENhmzD4At2MlY5CJO1a++holtrLRUMTGZckZWHkD0O224pkx44wiBY7G0PFB4DFQjL144wTQyuS
0aTK/Truq8qPFygvaDQ2tcCDY4+QGBBTdkKmIX26PdZW7t5BFUklAlwO/i3DKXBNYBSk0fpzT6EK
9QMrYypujDZmm6UqzElMj+4w2sANsUTmvx0mRK8naMbqTOW/RBnJYNkjCtzHW9aRwLgYEpXwW8ii
ctG53eZkTlV5ImdfjuEgVXDP4B3MvcyUbhsAvT5kTKiKEcduimhpJ35+TrTGLt+P5lc1Fhi7yDa2
oTNi6jxq0uXkg+dh/u9Yhl6MfeZxWF2W/50XhcnqMsVJ1A2IPj5tyWF6G6qxciTNj54s4Lk0LYAm
V4HVf5JHsc8cLdfwmxEe36n9v4RBA9FtAh+g+rNVR8JnILXbBXw/3cpcSmDV+dN3xI0GWVQ2xn91
g0yCxsDiP93Hqois3oJPHNIcMX3AgEAZWKXapcXA4vKDK7jLCi0yD3zAMw1YefueoUbNYjDw4uP8
3JjRaADf4RGFozWbb+i2A+E9DwAszccFnanLVks1grKxRcXWifLmrOMdnULJMGWf5PYeNiQ39Fwe
R/iJST35FRaJffg89MeRIUTabYABYZI++OY2qncVV8Ts65NDmBqD34/DumxhDMVI6vSGSegbNVQt
j/eIyKdLWZZ61Aj8fLJelf0QzJOC90xWspQ1oCraXkX2cExXpzT+3G80pgKSrORC8gvcAIjb1iax
B7dNCKDBoxb9xaHPpcPAH+yStK+0m0lN5xTMFb/jB11hL6eTscHRiIX5Y+Su6GEGxfM2SxKcsNAK
SjzXllcPhWecO5ZieTBvWgZNwvinfms2l2doKgb+5kiw0URmD4w7uAP+EvhKidmxiIcvSr8Gohr5
J+LNPydGV7xh1ezm/lOMZF08erG2iE7xGYL15wqT3+c9HjHtpp5ONpdIm/IGCfYfqRt7WOQlVy50
z3fLRAH9OK8ji8QZv9Va1nXVIqVvgcboIG2hOTCe/itEAmAkE5d0kb1K1ENQ0HfFT+bzMDWHpjx7
0lsSDuuOVlU6D1810nHtXhXMpl/sgdOgvCgS5HysICrWncCR/sC7poFTcRpKCzxvQLkwPfiXwU+a
Vou6abVM1FUMliRaKvN8RWCTczS9P4z8HVJKugK4Q4Tkv18sMnqTe0TrSuiEP8n5Lcp7WuEWZvge
6ksgIRETNcDI0l7tFvV0HsMmM1sbgLDZ2qW89gqQtHWMsLRLyCuSCpqwvwRdoCbuMj5hb/1d4nPV
cDy8u1zOMoAf3TxmLa/7g1838k/lcbkII5QnDmSA4IHJjNeY9UrIuunH8HQyftIq0H0Y05n+JXtK
2Hxi6URc9ApVK5QdSvMWcI9UxMO8hdgHVMcL/W6zYYBVPfwVa7W5q12LHl8n+rsRfSN10mXgdTek
1bZXqMefNZxSkyReKAcupRlF7wSgauqInH0NfTRHFZ0Ffbw31yWIllED0vNGpKemlU0EwZ9f0+Vw
24exQ3EozsBSYjd/X3nO+mw+mN/lobV/G6bqdlSeCMZYB4rFIIAGUjrKvIiUwhfdsfFzAKU3bJ1/
qHHpyH019dAnx+sV5Zja6dPf2DuM0bvr14Z7HbB2o5nHJ7yRwwhdYg4NwXGZ4/eUmRI/5xW2qTt5
b3dRNUD459vDks09AKOClrmU2A7g2t24tnyodhegmB/UHiKH8GRYMHA9Kazsoorox42WrDD1DOQc
xgzWJonMb07iv4V3YkHWhttSmuuEC3tBVgt1bVbn7/iOk0wbN1t+aT3L9RG9ebagxr4ProvmOGl3
1K8EPZDFA/6DQJQ5r9wkrSUBMANCok0UIjJkB0svlVpWfPibcxfHWPPB4tvFXE4y9MnDknlNZYGB
8KvVKOAhrVvPhZ0cWY18Zs0kfgtBZq+uvKnTuG1dePysNMeKxFSdI3Zf4E2+14QRKAc2CtLYVcRs
u4gtYbq5FawzhTdBeg/2vhreUBrvt3p7C7UiZ/3FGEwibJLPzWAMwWKIYV0UISNX06Ct7WL1lsww
l4Pvkr6mrRamb5OXQ0U4HM50XwVyaGtwa7AfhZK+UkJHteHgAERMyFTwF3iHJsswGXNEgA6pIZNS
ugKpA18p4xsinhdtBllb/M7tHYj2otEBpTPBo0aFMBbIZyFj55GiUxZ9F/9jfcgCfzXay25jDHjp
Ufer4+MZTZb+SFkhCD9200rTJ1JNVwovcYbIKIkNvIMeU2JcofZ3b1pL7vLk8rXfR5uDOhjK5vb8
AeVjFqnkoismQgHYf095Ek1bYiC+QocFvV5FIT3aWkffbDJ4F2Lj41U+99zwJuZyxCHPNhBM/QBF
t0IuW7YqktoKhbUKEQsmEynhP7nWxQKwo15FAOpCLzClQCUnMPyLxFgMZG5YyPeMbPDfbAXkbiQl
eRMBXgF3P7kem75Oi7Y9kuxUcymt2eFdLx6StZx+hvVLiArOTOlfHVZVyqP+0B/2saFCes7DmgvN
tiLkoy2PKcrk3cPnQ16jGc3DZjTlx7xMAJG6mYjmJGY9MajCHrTQpJ41XG4N9c/XdTKMiwm4129t
EG+2JeFvmxuFi/ULBwhDuImJIyvpFoy/qONEVxITW3EiXZY4L0pZrq3rGAaBjwCFTV5Vd2Vt7Pci
kXnmuQdCdl0k/y3bF5qiI7JRn6ap26XsfyCFIp1l6relyLIGnkYMQJs6S0x8s9KWTKbeFEQ3pgHN
S8YL2jIr0SzrO0Jh3pM8DhIm1neT7KMZ+GqzI18H+NJWoug58q+kLYOOprWimeQdMucSICXGPavR
4lHKvlvN0ZMMzwALtT9yd9EDtB7O6uXoiqtmpAa6UJ4hhZA1QqEBmDttrSgvqKkb+K5eeuIQvgFP
VjEq8vfweQQlYC0fIJvu59nHtmhd3krqD5Y19DfxEOAUA8YPpW7SaY2gPqNVFdTbWlp19V5gXG3r
4Qve675MZa5gAf6aWFQwqMD4QE1oQlYn3Xla9T76SJ/hIEdDQPsvJHy7X13KNxB76ZNOF9wCrU0g
l6hbNwIVEfJpyiZ7RkuOREwsA03YeluTj19zNeXx0e9nNg4+a/x0bZMx+ii33G0N8FyFgECtIeD/
Q9BZh8dUV0OKBEW4ASfCB0tX5exYfwrpKwk4CNOk4UZJx9nXi2nY50HNSe4R83mV9+34pOMyToNI
5g1kfI12KMrm2/VAS2dxEy+sC7aRyQvMPG2Hi0vnpBcY20rqULF6UmdAYDorX9QwZc1SIGqcjflT
m0HNIPQY63cBZv7m3ikZ7gABBSZZtNVZMx6+Nkl8/45hucV36wqetkr5mMv2ugaCUcEZ1BV3TMb4
61m4Bs5iLs7htmvdPwNG6L6KTA56KQoHf+LWG6X7sS9hMEhsidIjvtDYqy5PC8OYPwVE6wpuylkq
cNGk7lx4aPEOKfA4cAtiL7Fqh+hk6AzQbWef8s9kg/IjOvn3SuO+IDywWE+AxZps15AtGpGHxMcI
NFYCAXl04VoH05RdMoKQcE3UYxylqo4JNeWt5lcySnGyF6Uezjt1sxn4srrSglJDOVtQZigeDwrl
iw/b2MgLpPk1KL72hQVHJtgv383AchuViYOR9RWvuFY0Iq09sYmewc3HE774G8AI3ran4BiWwqoh
KJA8iYg3IsSqT72ug5zjgFIKpa/pt/eR8I6oEdEtLkCb5nbs7gRsepHjGdfOOOVH78WEX4k0XeaX
js2xz22cvxIn+n2glZoYtnj2+FJs7Jt3fMgNvE6hN3s6P7OhVIgBBl09QwtHZdLZ5U2HZUHf3uLf
XAqBdBr5lICNn9kNji13fnMZ0fBbKZ0OPzzwM63XLTdjUC9qgonu5+K+rIzyAm9gSEjAlB/o+gOn
xM3OcqsoFMf1aprq8bTwaMjmgxLM/oIEqFca79FRiebLgeNCOo0hf+hs69lVp63LzJAcGh/JJxoI
jWm8kCoNY9RR90rSoRQ/80iTfChcXOW8Cl7vqV0Rb/i5MqSuUcZVNXajkPgw/9xf+jlAD8itJQbJ
oZcMGv6ulL6h+RTLI17asDYYoyytw4h2kEz1Jq7UpeN2qzZsmYw7w+tN9LVwK8lWFO1XvygOEKH3
SZI4GeX4Cj4R+0lgq8UxGHV7WbpPeUvXpQUH4JDAZA7MPQz2QwDHnGX9156Pcj0piDrYqGiobth5
KyC3gPQZYomysHzMtMIUn6pQ18lY7+j4ABYp01R49mUcFyCtmuk7jqmQ64udBuwjD9Vr5pMzJCt+
MqwxL++c7Mot9upXlv6C9tYli+0gjS0GUf1LGQSaZ5ntCdj2vP/J1t9TWXRAzBHlDgs70mfKcpbm
PXkNhLIWEgkLxUc4tH+qxMpAnqcPrPx2qRVQa3q3b6bWFegMew6MIEC9tDNnJoN57XZ1OwlHo5Oq
6KVqE6JQoFP3T2b+P+YmA21hWAoIZLsCFfIrpI3790zmsJIe/5AXj5mYihDCfedqz7g29dV5I7bf
vWHksswHfVb6yWQFHNuMAjjgzWf+tHTBQLvQC+DV3RRh00v95ffobPy0FT6buiraf1J/DdpSw5mK
32NCYSGdB6HsVW3/jUtizyhG1mxDumxlxeIeQ6kZZAOMWxO5dvEIVZMKJQR3y9wnDLq/TCyMygHO
QA1HHx6b5p1g/uJ+PaIkx3Wmj4wzILhuoyKnGrYxRccGGaXnLugMWxHGUZkWoLDoRqIccrJs1Fdd
YYv/cS8+sGKRGXk+id0HmS6TN2gMy96lAT9C1RBirGcG6vFInEnICukH9Na1kW3iRLb+mhFo84BX
M4G3kkN2jJykZGe8CKwxblnUiQ1aajN6sPI+HvgdT1mXYkmEm+ur9b7zobHOHYnl6KtHu/ZZ5Eta
1EKm1GsYMOiDGd2lzE8GLxs041+pyiDjOWoh/paMUtUACq7jcHnpbgKBUUi+21oA384zhTtuzdYa
O1X15GtiaIp28gp94GOfTeLf3s4eUcyAGmCYw/a7x47mWkwOr9UyJ99Rfv1lJpvye0VpS6LiBBlT
t91Q3JYjSHVH85ymaXRjXLoV6VFrtY+NWnRu3TO6bGnbnM34HMMWTDKoO+kd+Pe7eREy0HnFw6bk
PN88xVZNNn3bIHBBnTJ2C/doJQUSI7G9cmqpWfjPi26qlEcMfe0VhC6auH9fHNeVpIo/InAsst1v
a9LKKuda4dONYXodFPbhzqj7G9t8jHOWj49YnS13EykuaeRvdx0vpG21z4sNb9yadajYbNRSsRF1
TIpUoE+IsVfer1yN4gvRTLko0bGi7m8fj3+GKDnlwOk7XWjEjvJ0ZzC4dKZUwGNP0BUKVEq3H49o
NaTeOOCDNwKSCFmprAIdKtdV7ls/m11vJDH9VQT+Th7srCZWpqL4VFYJm4f+RhsC60tShMd0GZva
PYwA+DW5GgXrF53UMNFbX8QB0AlwdBtUAk41yDVpjcUIRNqN2/bWi5bjNI3NA1S3g8DmPuo3pkwh
QHWLaqOc0XMrICE4Pc9hJq7p3qsG5wvbuftVjpj5aaCmFHtdhrs1BxsovOCeMHAkjHmuqhGzT6VB
tCCgPSU+BIXqGElaQGEHSjHJdp4scHJtYHFkRXbsNrXn31xU5tROMSYUZWl4cU7teLSXo2r4WdxD
EuE7TkIGLo1bQ/pDr0b+RPE06g9ZklrxH/l454HDNZKIOF1NQJhOA+b4/fYaObeST05WqWKlkxmX
/+J3xLmdLzp3X1QBpR6W452sDNo5bgi+5HXpZttsJnDcnRhSjp6i7lP6R+olh0VuLL6QjqQ7rhMG
l859B+5TJLwmwcj5sheV2tg6eZI8tpzmPF00ndv1EfAMruXfjnm23sYTIFQn/BxadITq8NwnSjFv
VTHzRM3dZ1/+++FkqQBBpxBPzpk8SD41sYA7ARvX7fEa5HUpbynROd5i2XD2MOUtsyBYX1n0wrgU
BpbiPEBho5B83PEreOQGUMn3KWGuAyggzsM+JIB+eLZoJZID8ohGXdzgpAAf48h/Q1GLCDmrC9jA
QcKqJOCVFRiw/1L/KyqtlQUq7XsFbjO/m7zpMd/VfpTGulIF6xYMt60ewdL9pn/rcv5kudZYnOgX
Jm3FQ/g5gXkkdAIgx7kdElHXXAhkyPMqoqxtcV7caoQMt2cTM9185MWYFD58AyFTCWSx5SWSoGnh
efPIwsmAXgb7B9X0mgez2Tl5pKcPhzyCdEwKRQwmouHG1DqxZkV7jCFhymWDu3vA46r90MIpSnN/
oB+koJLK9XyGMzgqMhlXXyzHNBGRsjAf312sam4bq1jblh7e0j9eaS+EF12c6hZiwDl/Si/hIZTg
RripqXXcIhq16IkoG/p7XKZGQpoDbp8ceWEuzf3NFxNO1RqfRDKt1JWD6YOPglECGmgILzEbmq4+
J66lyOxpHvR7t96XubUz9A0K2GRl8IKKH3nTW6XELXnv9fL6iDQaFwX74c4LECNJ+OQDpwO/9hT6
jlgd+GzQdBo1UoffH4CKqoGqP0mtH82cIMB63ipoazLeSNpTeCfPXHhELpfRIRtcmdALHx1hZeBS
+xz1h4M7PK0Pv3gKHJMbaZHPuibLGFDU3wzPayhCvh7aEdm0eF4okPA5ZWvqaVKTNCoUi/Snl5KI
LfnjiOvppwYQ8CivGfY+gwiVE5q32hieCbiHC9BfJFvG7XK7Pj2h4ao0sM03usshuhv6tP27LTvy
8OR2D8fr1UAvqyRD2GObJw5FDuuRsofxoWjmBH+b35RFa2enNO1YAPWhdbfk11NUtDoCB2Ib35/q
mab0lL6sPKw+bIKOMoKBkx804AHb6neGobeBvu1DteBWw/ocay1bI5nhhXmX/yCKJtvKYHiegThw
Kb7DrFKHANSHh6mpfsVeYzBFaZLU2lvF5J19BIGsQihfN6JsyXBoGv1lRA9rFRNpSfrUBg8TLJU9
D7Y/p2VlvYIbRXLcFhHkkctq0GJowBnfaTwU0H8gj49o9s/rcbl7WceGs2ZO2cG/k1KhoNQGjJOl
e0RogqC6ygWQJHCnBYK2/TRgV1s9rVl8h1OhNhQxHt48DyPOa3ODWCiNcQbMQq4UW2dqhCVpgWis
vDzVliOwyAIadUbdC8tiQfAvLAtfMtcd1QhcyQOCvchaDUQrh1oBTbpQL7O5NBJObMpuMIMwbs/K
JXsxG8Bpl7omTV1jF9c/nzfUYrRkKRSbNG5Uzv73MaAbJOttJj8zeNywRpAsvx2GRwrfE1nnS6Rj
KMMASOPjkxzrneg1B9gUWvKCA5kn8yYJr9Ms+emOmHskNWf+QYDbpJGzSFuYYyK1Gp2flMpzKch+
LIEj3LArnQSZ6QugWYOqyGCJivoMxk5x1f2tKgzgXCFbLTq/dA2TJYm3BxKrEXKyw6nngE3esGUU
a4OSWyBKsuD7vTtg2jc8nZ4Nce9EF7qNSieZn8mz1evmYQHoJmqErImf5uQpOj9x3eHcN2PU1aqH
B9Kx5i9+K/auyASvHOxrq4+2piFMh3igdhvDQSEHjAlIUSjgwHY1isaRcwRISe1boGK++f4njI1f
u9RQMkn5kadeVGzkbcXxLtbmX/Ti8gNbt7OZEV8jgFXxRBfLhuZ81JJdxwwElAVEmFSNhb4fKuIf
fwFiDAXh1n0leu3Lc2+1TDs3tOH0C12KHGHex0tjL2/ZkO69Gxow8A19rtbC4GNwXiNI8v/cXoW8
oH0evhd2TZY/oZyDN2Ue3TSTUzgLvYWyy7hgDLjYsaVmKVLapun14jlt8C1OM+THhRsIzfcUoixm
idtOnfroQJD30A+dDee1+SzTlTrihS6d91N69NF6pkLlBfv1gzYUI6sdcFa+Myj5gbfTYEkhuI1/
PmOdBL33DTBqThQALDpgTNYd6vF0ZSHU75YfWPUpNiKbxIj2IsZHDfxbEdFSegxbEgQkm3WqNyMP
ESSz3SPfQ8O677ThsqMfzlKigPj4mcINeFcOYyjbgL20bcJWROKLfXYHHW47r3HwHJ20O4hiQvhS
ZjvT1S8ESwvyl7t/RZgxnMLFZ0JZGmneqW4QJDXk3+pQ6IlqIQbR+zydL5AqQ+I4OCU7KehZxqFf
LxhWxJBP4LuveP1nq7Xeftu+5XdroHlAeAV89HsaMb19puJnDf1qOasUgb4UlY9mBPxuzgjl68cD
oOSQLqu9RCU5kVit1rYEykd8CzVHoDvubTSmkA7AO2bwMduk98Shr9Uh+cLMI/qrm1SKsBiSyK6y
b1bFCKQniKpjr70z5LB2UfWThMl7fiOTwg+P3aj6jtaHR+Vlk/ki2jya1uSFZCRNkgDms0KdbZX3
/wI0LkWcMi3Klt1QluqPCLDDXmt/iZXBWdp1KMa2/SVybUFeh5gQen3CiNkTVK+394mytruM475v
BoDbfLWBpNprgt1/5I2wrUysFLeKGq5as2oPOJTmXQ4Ca4T2mHjxaPzhfOVgNfmA0F6JtUVrc6Ko
e9YFCkAWcASRhEvKcy4XLxRBVCAd6pLDMFQhlzPHwx7AmdIzyzEJexVm6Puen7U9PNLaeBd1MFGR
MUl4BF3fN3E5tOt6k9bwX/ruSPQnx4VRYtonFFQSigcP2+EEd74eIuezIhx0ZBzB3tjVtFkG89Jw
zLc4iwDokroY9wphvM19SOfNGhxvkzB8w4UN5LooEyRMd29x9bSSZYXTUpFcQnfeVfL+FIqrPiYT
YtwaOdi7dLiYdnB1MlEw7mfV6l3cofeurzTyC/bcy0BX9Msbg85qeUBtmgFYLgMh6NEoDrdg4+N5
aav/K+LMNVII+rCmh11vTSHP9J7UoQeAm7AWsveAoeTeR3wbb68EMeCiqEs25O/hb2agMIUxL829
3YGSknNcHJU8SATOhjAvHLEt1yYiV+xRE5E+ztNo7AcxJk4IAJFOX5LYnO498+UQ9EGdAVxQnj7t
3WBHPzMc2vgzNJkDcJiaxIZaGrA/o+yKd5Xog1MaXdaVtB1rS+kGpiMHc0YTAfbSBOCilmu8Rchb
tOpfPW3AH9CzyElBNeG6wfQyI2TKAlhAeu6xEn2mp6aBbh+Jdq+G30JkR8Fx2MhcD5b7Uf+OkRyj
xcQmIwmBP6Ez9h89q/gqvR+CkCojqCXHzgy8yxltN2q9TaDK0mPT4IJqm79uxeKmFb0/r/fjhyLQ
RcHWwS4apLfalCsdtuHCGWpM18ISLKy0qVA1FJKM58uzKQJGU95EfJnGCgS3N8CP5lg1S6u0Q4FH
YK3muNPcY4GOVWFCx1wT+uzCyfMq1yX32jMk5YerbC/x7Bg//VJToCkka5lwhiHgUa4JPrtShd+T
GIfh3KUDBQh2O7EFKCL0kQjiE4avXfcegXzukj+VXPk42GklOHV8jAU/u69TfWmw13TMWYP/nru8
tVw+rb+J8oOBlKq4jQD4L8Os3ufNC340MSoYsFA0BqEAS8TSEtRO0DADZVmXuD18UfnSA+8SQhQV
ZvAuVRgKyRlayY86Z2sHD6i0VQ/M7fGIwh84fl+6WzETt2CdiB/N3czU57bJaqvSUvL0n2Zgw9a1
OW4VRXpi56o7+F3CDHuyheALrr7Hly7AwzsqZwjTp228AptCpIWAFg5+ccV6cV5WfU8sPHfo/cLT
PlYRYwf106EFBR8KpQd+UStESEg5Yi5WpUuv5+bi/Qc4WIJUpROsMOHs4dPqHC2JSzfKezhh6V1C
y7mKF3BiWnoHYDNP+Hkscr1oPnQMjK5AetmDA2qyUDEpjua058dsCxrtVg38rhOs9XT1DhsqnNJ5
02+xQ35WBj87908aUov4xRnk19DD/fcTSZsrymqBN14+JkCuHXOsKnUWZ8OqlavzyuJ0EDLzdvtc
1KxprYgumID9k+DDKgimPqfujOr5JHSyh4OPFmD0VkvIPBQJK3VKak7jir+BHSnaG2XEpoKT759R
KSTXr5D8gOQnj3l73FrP31CB5mFd8GColuo1qLY9HpRG8MIqnoRaahyooJy1gIm0ypVEjLS5Us9n
Riiu15MMwHpl23XUQwCL9UHvwLWdfUiDq68aViosDaY3uVMvOAR26IPTLffa8Fd8hbrN0c+5BQSG
S5/f+K7EZkawZCZl0ym5SmEb4P1uF7mEeVuNvkULifjVpz4585lqWVe5M818jdBtWoSMH6SaFHON
v2lIlC5y9LwXSwHiS5qwDW1SAY+F9l8Bjb7FGZRqgIS28qfjMsUwEzq/N9PpCtGWfBEHfBIoE2ok
lJYgVfR252kpJiMyUFixCtmxvX11f9FZ+62HlcofkT7KQJ8lo4h9NRH+Q4l3w649yc76zGrF1uo3
kdlUiRw0Szo2Dwa6iE5jkaWbBE8btXTewJuDY+qNhgL/Kw7rVzx8SW0vnfY9kM8/NouGNvQFbTAw
ASZxWkiuJtlAMAKGMjXQoFfZ7pnybnzOY3qkWXYBQVQ/NTvwwyE2VqzSsIpZPZkDODOkbg/op1Aq
cegEBFUaY/8gSpQ/z1fDR72MMtKzffTxE1SYVrYjN+YVuJ3gANk199/vde2abBdyCLFTX2lL9KKx
Z9+3DxFvdnN+6WWG+2/fG01N27Y9nZGCguHdcZYXbmWSqQwiANtMQ2NQMREjm09WBi8aQVATbvq1
f9TufDJkW+ONpV1nBuEWTQBwgtsXpKhjd5kl2kUzV1ys9wm+jQHzv5A/bDjaPSMUEFTP+K9wXO6j
TeqgXU//9/dDmIpSqqyoEWL28W/NmKEfDMhBQFqmykIksumD6egYQr8dbBj5RdpZ+b0I0FAE3K6w
PvOojMlUUTNMLF6DF0uOQRv9/cOvYMjMcsOcOYQaxIRtdCNwIpr4d7Ni1QvTweysUlaeWVYeiBYq
UvIAn1DdPweupTFxWBd1mliOOdEOaf1k7ZHe2K7O/8K6VrcPajXVzYOIk04m1NRqEToDUMiizaBz
/Y6OjGEQyDCzhFoElh9ZLKA7lYHmN2ijYIZkTcQxlHktPT7bEScC3cXJNdWVSZBTvPlpjwTgRZZ6
gTYJNOiG3ZFlZfAmBHFLzghGDyktkm73XYRKob042LbTCOE9NkNwuELSEwu5S/YZMgIjKZEGYiTk
fTGQ55IPJthZzsWp2BjZwJA8azicamPY8LoIv+OjFihW1pQ5wXEUpE9cbfV+5YCPfi4BjtkFjk/l
1vo6rtMsrDzH5c/2hQiFUympXAppq6a6Ebaj90OuevKuhqRXD+80ym0TSykxxfKd7thFWVw4fAss
L2oH8ibNbtwu6Ofz4KelHuxVCUcKrxwpDq4dYwRGcltK8HTRu9oz3lcZ+d3U5QQwW/orwCxt7bUl
H4QAt/1BWdnXYLDN1ltpRCTNGEiEtQkih77k6AV6AIO0q5lsqwR+wbC223xl+IVu6KQ8f116VGni
gW5gCeOURG8XbDE8yS1WBKuDVUQL7d3X1p6yg0Lll3u6nuuAAJzAHxUX+YfNPDp2xuGkXrVGhUM8
Ik3jbVBdMJOIK21ToV02+IuWGETdgULAgX863G1z61JZvCDvhk8yeFFjs6Mas6aj9gmdeNLstpI3
oOPEnQxhm92zIztEoQd6oIjip1svD1aGYU6aBx+W3Ten8a6lRIqhpBCwMA+fc4pvybi1MWlMiBge
Rlmgi0/O23guDD2KMolaLpcx3v+hAunLLsrVPFpCq1CBNpM/2w069NeBb0y+2mtlL0A40CYauo6+
J6lHknWWkWLblhVu35iDpJgjZDj8TeGUkUEGHhlR/LIeDk5tNjj2oCN9X5rbti+k1iDFeK9zHHXZ
Z95aiiD/LmEnCV+Uq+aM7YaNGX4POPo+gr9gfDQebXnYdDqnsTGA3VtwYtFnOI7AbyhMDGgb4fdh
8U2VFhkTgjCCSaq09Q1fx3QR0NfTjBXF6UoD02ZgYM5mLRnngae3NmQ3PrU4cc23Xmj/m248G8pj
0yUIOSgri5OyiAAPiAWQ4H11wSHyozKghyzYeP8UNMzyCf2ERnWdaJy7XE4UiJ0c0CeV0txUeY8W
vLO3GMSP6IU6SRkMejxnVZOVin+8Xm6rwWurUxsxEcOO6TXnLOQJgl3i/RBmo0ex1Ur8OHjVLUq6
JMaiI8GgNrpeP5IzCYzMXwEW1k6geQkAYmAqGlIjOFSeQ0m1BE0UWajkxhj5gc2Ta7mu+P84qXOt
CrA8h1jtrEJHBMmE0KC1G37Uo0dNfw+P2JeMk2dOJtmgBJdBI0QX5U60c8I3rCu4ZhNcClMp4qYg
mshk0S7ZcaZbb6j+NwceRdpPXvQ486svh32kkDhByoDyDkuvxwYKrJNJU8DwTIrDdDAaL0qGlaPb
COW7oM9FBZ9cNEZzjabd7J6sTlmhksMryamc+PbxCsvMlXUd24XOLXqiBbDJKOk5WIJnMUQ9obAW
5TSnFSSBpR5pUOepMEb7FRUAV4BQCpUb0bialE8B8yKDRxklTN3bTamNRLOCTvBCdFYkJOJjRFLF
Pz6zG8Ed7D8w/5K5Oq0Brph/YzdS/qakA/A9P/Al7nAhZLFrvjqn8pViafMdxsqPLWM8OHe8Rp0G
Gn//+kNvhbc79kWKrxVttksD9uBgBEPngqvTNCBumjRbqZJ8V9r6oWqPmLW78P4RvlqKq9OqhWxJ
c9xH8s7UMW4Ctdajru//xYlRtQWSDtCFF2fu4QC8TMUpRQ0i2Apdrp1uV0pFrJly0jRakJml0EzK
cPfg3ATuzxfSpbS0OEGqJ7WFvmxqQHpT38Z5nckbjQlAyN3jE8TZLwBNbrzR+EVrLhCCAnEsTM/u
PuJcuYgaboVqAz4xPmybMyJYaCbt9/Ht76Y3U7/VNUnn2XUE1UDPySBaG444f8rLUcsLwtprjPfR
BNUFl07TY+TGllGKNmPtGv5Wnjixwrh87ewlwnahcLMJdoBJ5FbSFjOqEUs5YgmDk8yb8FYabbfb
C0tHf/DeWHGKPJEPJlaXNRhi9zVpyq7M31ImSxkR7JuoWkVUXb0suif+6xbimRFXOS7xcyWddtw9
scvf7V6yEFrnVYVdPGFUw+bbAdt9SSrvW1YKBorO6fG/vIl1nHIyr0yUlO0JwQ8whRwksEzrUGZO
9hKUM3tO5aS3MPQ3CwLDkdRjtjRv/7jNo+2ub7Jk/cx94tD92wf/YazLoDCgerW+9y5B11rtUjhj
DRjBdg4QAnk86p9kZyFdP3RyoT/jWDjxRtK4mz5rQOz0dpO4UrAtNkiNouTcwoJyNFe3Kh4wP+DG
XtVpagOWpUDxHx+68v6z9oNylqIMpqObIQ3I32fp71GTXZ0M+v7No+ckBCHJRcIEfVq406ROVwyc
DpkMsBSnI/5DIYI/H0Kypb1MqzjXRTyTz+TJRrCDfzPyeAt8XJ0eNdLdsn+7OJq7gbJ0oWYUqaQV
B4c5yF9dgoNpLdk9yGQ4USboXJYZulAPlYIIdIWONKUC0hIVk25Jx3VjZpb0XYfllCJXmbzcasS4
/XAYTk2aciqkEkAJnt3yZBwqEpaYhJA7Ze8cAP7YkIRPky3WKFfeXTpmHD2XRB7MHlgDs95dL9jh
19/alSpxq6uf5GNJZNZK1Pwzf8hfcWzuHg5k33Qe24yGXUjSiFSwnleimkrRownGhpuq1RP3TQ3D
iuezB7DLfBPqdPLAfz2Asl1X/lD6rD+VBrAeqkOlg5MZjl1sRiS0FbfCmISleiwfoKSHC/NmAcAy
IsGK2eZ0yHFiie0m0ivNeKu3vk57nmBXlzKz7KyhutSMOneJ3yOWB1qb4pljcM9S2d/YYEm1z0yW
WSv1opwQMHrhSTa+OVVMOwMCfgwcseAbGuGBDZhxcyWs23hLV8oHWgt61Tnbt79BREtmplXZx4wn
nWTM9TwZg12yGL8JFCXatOZ1o/AKA6g6ckQKsomh24DlWWkxkGf3VH/pRCUH/v1dMc2VDc8Vh4ZN
58bOds6EmmHDOKNp9lq0dv0HQhsmF27VsG7R3VzdAwSPlxn72j4LsdHIDBQ7dZ/sQL3yi+W+1Vzc
aY4dxEmNW0XKMdymebLcQcqTKCMJlvfUZJDwzKBXRQBClvMVDZypFZtXIxI8LCzONl9H7OriRqT1
GWKVrHMVyZ9vStmYxmKVobBRgeIENjhT1AqY4c8nUEnH1or3/kEmX8zxfeSYzPibT4Z+39rgxM/R
I1KqE9oDh1mfOD6ESE0Ufny6HQJysnNBmo3lEpJnEY0O1yCmY2EVRYFHLuqLc/ugPZRvhK8uoxz0
rxdPRATV/uONLXQbHuRj58Yq30zUZI7YPRDPU6mBnC812uisVn0s1qdMfofFsObjAwOx9M3yINrk
Ad5ldjPLqgH+5iPrLXL++OHU7voMBFrBLDiqcqgTigmy2S5V7EC7DJSQ7IaFTBdpBrKxLwh52b6X
JsHCEiysZzB7fsQw724V5j1c+NQlBJhmeUuB4x6TYEpWIvOvagtT02Oi9X3ygXq8LLeH1P8X/asV
hqqaMDYx0Y6EwN9oRghIWQmsgtQQL1rVZBN/RJplNi1ZhuA9KYKWKKM8hIL8mfokI5Et1OzJeAjF
pFy/jUPg/0dLlBI3T4ar1yaY8Qm8PTSzfMhUjYQVYizIFPHkxCX2O3nAYKU3B42QBTcdgnx9RWUD
GFwhHD5oPk/pUVLkcjgRnLmKOgnRjcl9DEC8e76JaavICpUpw1DoXBFkIHH+lkhwKX154L0IR9pp
ft2/iKPw8OkWZmjEPeq4GUsahmr2ShZDBSUYcXyMOjkJ6N/ZU9TSso4QxApr3L27iccGooM4oaH3
r3DAHdxRQB85Uelh95zviNpksCLFzt09tTlzxtJsNXPeWIzxV+PKs8/t97h5x1XZdlJ8ECvJrUub
kHzIDiapeBkku4w+M+QMX2m0ZzaRDrN29Nrc2+Vf1RJ/Tq9e+K51L54foPgizjO1w8RMqn20Y4gg
d+j8cPFXocQ2oMulc7Ofum1/j+SqvYu/JW3PHtaaOhLKZ7SFDZ7kdy0SWt0d+hKgYfeXweXizSXt
UH2VLSG895X0RXEmU2h9txBgKGUb9tNGD5doS5wAz4z4GDuDlYPWYMF5H8kiHLTneYXEckcpmhcD
IhqVIgEMvpoxXQ0Y+VIMLw6FO3mcRlS3sSeMrk23PGEnon+5O5Ra1BkXf6oeE3Q82TeklH5UTUJf
jgVYX1m0mUKD031bv58YuZ2n9MOF1mE77clgWX6WfEbEgSrEsNq15YqzzpuKF0w43ITZvwFctkJx
VZnfGHg7PGxtm+V59p3R2mqahxYd/MnWEayHoL4BCi+EEEzqHhIIVNH/OhT5zlALXPLgpz6X1UBg
f7meVXTXqY2NLrRJw8a8+Wp/CMnvaZcfUb+YgQuDMjiQyWluXfYDcAtX4DZYJpYYRqhb37Bu89K9
oazToRg/D6NiD1ZS6MfV/63+b/lfNaRuwXkNVPCFAw2qU+r+rN93UVhxmu56lTtZ/QZUc33KcyP8
mWSzr/S04L1cM72byYWZiF6Nl30YSHaOoJO1ffWFyjRr9SZjPIRft46UWyvSfMpYtQZlkrZSAaUC
gSwUVn/BXlY7spEzj20c03z9qX2GNw8GKlWS4T+RSqcMEMkbnZKTT4t72Po6Tvn7VTEcjg4DfIxl
5iXx30YbP/afcopj58pGMoZcIR+rAIAbXhOOx6HrimLtb6vx3wSA38Zq+McxYVXJ2GpnFMlzkNvL
B5g+xY8I7LY+N7X69grLRIv+Qct9RRrrabXsCpCvcg/T7Vc1PASz1MYLoSUkkPcxr/fEr0pS+BCd
LGaWSkqZ3Q2oydT8ZvRpS5YtQJEtNQADhOTMcAvnd2gHqsTFiEP0S4M/XUKdhJwH0rhoenTQ9ZAB
TrvErXA8YSUoYnWTaYhNzyI9SEwjnmOjiWMMrqZIXaJ5Pt8SRvX4UGPESogGtUcjNDNiV1VZPudl
mTateF8VIcfb/myWO0aWIk77p7os0Pjp0mMRGdrSEZLvY9qgzKZ/RPn8m1zbaZ/3jGvkWHDwhF8j
cTjuDA+3LEpry4al91fudjX8NfZ7T20HOtsLqo+2dd6yyjXOeURgsz3LWi8eqYB8LFkovLjwjogs
4B3ZoMJAXZYLejRHFSkk9qUtU+eF4wZRbK4DGNj8GSRMs7GxtXsapqe9AsUgwP0XdqGbdE5G+qgr
X18dUeQYsdB7M3mDxTAtmuKQH4IfHcmY95JQ1QCsMSHTdK06qe1ks51BEdgVWs06JA/rLmr9GptP
mwos7W/WOthxjmRtWe4Gkj54LoDmOtVyxien5XotNbnTi596brmbqak2vqrK0Ok4+iiGUygyWlhH
QtOgpapMtMFmPH+6WZbinHprLXP3W/hS25oNvkDufeeHaatHu7t9dh39hGMy/EKOrIVwcLTfM9Gw
yU0s7At0xWPzf6U9JXMkSZWXQOrCBhGGHMrBa6F0+2jOIdhfkXKjI+R7wpzlacYnG3Kk41xcJHmA
ILNulOobpkK0V2OT+QsnV96Cg9ebJT3rDT+USoR/LllBaVY9EYamVLm+rCKtX7iitG/6ctX4BXn+
aL1FDXWEFHabZjuhRYq89w2unmjxfzcRj/1+UA+vBmnIvwQVv+D68Pso+Xk3+PsYr29tx50usf/I
T+qiyWoXUNKL75zDsM+fQK0jBSBp4/jTjOXmZmnsyHvxFrp4kcABs76wpE0qDrAhWLSeq/kF8Qvd
M6VIF4v0sIuyBLOCKSU2TR1FSlXD0j4Zf1D+hkYBEpP2qjYI926HBE1VMqorF1ngCOd+O2g+iY0W
L2JK3UVBNSB582GNxCpJbmSVs23XMRw6TG0U2faCYWBqL3YK4t5wIzL068z09ROLc73Xansm8WG7
6ZsixLnzwYExED7o6McKIc2uAQyaAIPqqG7LdOYJp7vslnCJuca0d9qLpj4qRWuaUyEHw4YcazTQ
RbCTvxzTeNZrezxBfzxvYbD9cMjQtY2qH7PtQkO3QfD0Kqk2wmcpjtGMVcxFn/Z3gD7P+jV/q6lp
UBEuR5jf0MZI3KTHkM8jDsZ93jxHfjETpEc/Vyu8+5rwJ5RMVeGVDfEexFYIEnpEw16SAWqB+/Tg
10f/DcHedsChTReTYvntAyvKIh/aywGiZpYGuYiJFsjkTTFnH72/dwD41uKy4emHXExfiVfqkoMT
FRcAT9/DVBCKF7LFLIpA364Uz7pHjRbtg9myDy+eJYt9yWkaqJndu8To36DJIhTyMLwKPgQhviwH
dLVNi1OL8SC0TdaJaBkjFWZB7HyU3VZgZl6AGt3ihWUPbPSdXhhmcSV+7ghD+ULo8k5iRBVfLiui
CJ0tM8/l9RDWhzpYHGP20AYEGcNhIBHlKIWnP3t/vRFHQz5J83aKEjBG/ubAdo3GihYN3O0/hWbe
xuRFukL1siUxj0M5o8JRqKA6y0R3ojToXUz3Qx1K7Ae4kpXjS2zTdBLntNwULuIHtN3pDPlwLMQZ
eZ6TTwjtU/T1NwJkpXH+DTQRtwQkSMzSz7ECFu/Mt4VStNYLR/EAWb5ag83UELzTaSSSNmuRE+CM
3CrzBEL4ZvrZwUh4sednBGodU8Z8LxMXep2lB5mVl9tj8mDcXTYKTIX8kIJtKqgePtwVgAk5fUe3
6Wko6HAKAE4QJlg+Ewctowvm439gcwQileJxCBnuVInHhJiuxYC4t5XppVn8DcAzNYA1Qp5bOptt
wSq6SMLWoz+VZiUwjwTsDh9SfFQhXq6TfxJZcBywhjb3t9kx8AUWF4YGOiuc2mchEbz5YxDTJK+P
DconVDjR3AeG5dD6JuEgxG6THK+/DSozq/6hgmaLUM1stOskvS8KmPdl0d6ULtBjAUQDtmxuDbU8
gzWmid+5Iq1TfW1NGJ1s2JUw/+c9tyv/AnsBOEFjBw68sh98mU3WFTDWt5sTxulQ+ZIaA5BvhmZf
HN2CioNOBIHqqFXDle1Lg+t3xDAR3+E1hlopInhoMOmxtzg2YYRyynaYPIlbX7X47fg0ddQ0llUQ
T3rwWLRwl5z7rx4ibDSmUhYJXeOdbJIiXHFOOqENPf7nkTmVuv937ZgGyzBDNYd+nsFJadR6oCpp
80hY+Fka5iaQ8rdamAkfe1dRceE4LybDT7oY/gAxyaFB2tAMz96AUOJC8vP5AIBYbpYR+uVI0zig
Un+MST+PAmRSTL8tceCUkcEXEpJrH2KqaJ2G3Ww8FW3vW6rjd5j/TbBr1xxoM2DRDElWbuCyOFpy
E30jP9sIhFrhUKy2yyTFvjcisvDmdZDo7mfmOnuj9QGX7j6zBruOj/qckOnL2wR5Uj969ICJP89N
dXCs1xFW03Aee5njsuqo1sc+dFjgkvr6bmUGeDinzRR594FUmH4vIKM8glmMZMnGzio0eVeVzOZ1
MReoY8RK0j++Gb2N3qvjqGnhnpXoXUovpqhRhwg2tvbvKOoP5G5/E23rj7xwzofJZK2db+KlLXkt
CjOIryX8OZkte+iq/nJuP82Y4xt5kz0Uy1tp2S0t6Yk33D618raALTtxOnVml7ZlthfpyHeySroa
OvfY9Xmyt4z5YtIU7yBSVUSxjbciR0g+CJ8ZCkW1N+W/yzHyaoFKBoRdJmsTsKOXVCk69ez2+eoE
o/e/zPjHC7yRcz6VfgQyyIy2stiLzdEMZD3LWh9U4AZ3KBIi4y/ROeHN4UKKq3NOeAP8v2hBVxQX
N3A/b3tsdme4RI+rRx2LdlPfUAuOVKq7NtbANkgEF8yaSSF7yvrI+wa9ajn9KprJaVVvetjMBeTZ
ydX7EY/4nlPaOuk1a6F7wawjbzvOQx9HXLkBTUq5cUL8rhWreL+wQcOCt7Kpgx7AeMqrinDLkMcc
OjGVs3jXyiEDM6JRI4qQeilh2QSQxVJg9VL5yQrnwiazZLaAXTIMteye/GIUtfSWYKLHp5ruizuf
9VmtVM8lh+evnjtks3zH5wq82kbHm46cFnSV9iEDSqkR8/mNB6YBPw2Aqz1TcBPT5qkjsjYnUJKu
SkUf3o91bLco41z1GJ6JD2zrUOuZ5COEZaFwCRNz0w5/VBkMJnuWQiADXhHrF9FKI4yIqqDeONtC
lQTgYlhuaSWUqfGiRYK2m2tofFLbhVpNe+sksStPlcZvhQMOkI6sG9k4zsGWJbz9k+tXhQW8oboo
7vamXsmXBxg2tUlcgvNEsCFwkjs6pMNTqaSRDEwaIFIrNzEn9I/LjGGuhVxl1Ws5RjLIfykhhX9X
7FDkQF34jQw230ZJuRei4De2BWgHegbv8JAnemyPRGR/cGxj9dO4L95sdljVw1+k2dN1N/faQXP2
3J8SIWMYpqAYaJg4NGBqGLrliSqczjkHNQZtTJc4WwX6T2mtbLEmjZghnEqLuLL6oEwJxNkNVe8/
OrneHdRLfncdnIZKMpyfDV9R8JDyTtgEC6kL8M88evkaBuF3yPp5mQ2FS6FJ2t+e30fCWMQUVZb5
M29FZXIdqMfnPgsPDjFjRnuast2NDsWtl0chuIL/eG0VtQl1DdGfvjA9gjVdf/PnUlkLlLHU6Oxo
13STRp3JAQA1sUWWRWvzpcArfRO8LRVqc2TtRnlSIQ+kwBqpoXfFvdvYBKcmVWeqmoCRFBxdz+fG
ykN60j38KqK5RlHL4Zu7pWVKyGR9UuLyvFtwwNu25Lx1n6EHY17u4hQ+9DfsijkmxF4wZryNRm3R
14AKK/0pAJ5mw004grqMLqBkFoCSYuDLL9VBv1AFQ257E9aSQeMvcbX1+qmVlbcHV4h9H16lknGQ
rDvQ6W9dqWkKnBUog+pvtyUUVNxasImYQBlGgsjfcAq7e3WSft6YGZkrrvF3lDfSc+w1+MPv87ca
w6UavGTkb5MAtjEh3nVBo2L90GKx+Y2QqkeYKNPX/D13NCIsdGmtJcbwZX56ggvq0WHyje5ibMGb
VEgAbl6MmcVt4c5YrM9PkK0te5x9HovXqJFpsp1tCTzke2ZiPaGYB90QnECFX0dYh7H4QxizgaLV
gm0wzDNPZTzlOTpOwEFQnYJA1Hqk1dbVEjaZ6fz/pcsFFZD0PygDaFJAaL1IEZiCPl568jty2bXy
fWGNqVmYjolBOMBDxXIgZJNjBZqGVgQz4K+C7clTaRkCvZxbLHSFF1TQRgwlCTSKVIN8eApAPI6x
wjyJrAu+1m4kSgoacQxvANC/H3pdB6UoFUzk8mo49UszbX6eK79sqp60O7uQ4TbP6tL0B0e4kNdV
LNtRlxTbvR3I3Y+gErC+bc21/Z6H6CIajddSf2el9XF0VxotQ8/dlagyU6XPPKMxJU9dHBiN/knk
75VuO6RGvkBkeMdy7qdbmQm2imrAa2ZJwgHHI+CYLZwcLqluKS2L7Jj3A/dU6FKBAzESYEXuXXtE
vEqXbFwXYS7rPiPaCEtIgZaU50UQ2XVQmvWn8wiAzPLG6hOa4f2tFkXzp7VEESD19JH96gyD9p+X
6vrACRdZOm39qsqixJbI2KO15KEyKGqprztOj8qlguUbuZe6cukURhE+Ds5M4rdn8UK9sQwFPs+t
UOIMWZgPhfgtIfw3aXiCaXSoE3p0bgCcU+Irou3XWwjZxJemw25ZuGulE03wSlQzcHJ+TEEwmDD+
Sm36HROmMeSz2YcsuUqO5rGWTLd/OS7wWt9sGic2AZtSuLLBOFP4VVJyBFoh/Y+b+NixORDmTCoh
DtLO6kiCphq9wW/mdf6c+liuBmHFpJDSOSr6tXq2/R3oE99AQYDPczLhnXIEbwf468nw27h7Y9Id
+grDhrcwmS2KhNnr/3mdRgj3ZDe9xIimKaaCfQvA1vBMDsIFsbh113eloexz/+wDLLTeS+VKNgYP
PPkxpueKyuDlxlZORk8GL2NnsH6MtGddI4hPzfru1LuYgHfiWmKZf4rtzJxslVrlBLwMq5AbJNkA
srwAMu9np2Q1P9PamdVa5qohHb9+uvjp5TLnMaDZcSecGxX8cKjnv7j5avPfLHzHA02GbJW8QvYY
fywSzaPSpuXLZKyfByjo9dL5nN9a/ByH0HTrYIiNoXae+khbd9ZPQVbf+CmUSwK49OBR20UeE9gK
uDTWT4bWgZdCuSEo4ehgCe4p9TxjUvgl8eL/Y46kPydgjWqipodtPsM14bzgB/qPq2TKIyhwpEUK
5fWgT+Pla51lGcI6H2l/PU14z//E73wqQlK/tZM1uCoHSv/dAqFIK+WByf2QAzSCbcW7aQBP4FjW
vDSFvZCdE0ikBD1BrZywRkclg1CfwUdPdNVrlQePhazfc0TN5oWXHm766svrLolPhj7ehIxnmZjm
ArVSWBrE/tHoOG3b9k+GZ9xoM/hosJG2fqc8dPx1Hu+Ac9769u9fhY+WlZyYnuKx7ZtVr83Trcxm
MauHFuCZSwMcwrFdw7p1ZuQvHjd4DYcty0Jkd/+VtTtYBIPkiGQhfZb3ui8H6NdJ6a17m+6u6zjb
5M81Chm2oNGsqh8Ua9MCgaqNPcqfvwY71wwQ9EkFho6Iz6cM59UDLkwsvt8DuQzKq+WOcB3Nzfrg
ighjtguv9lv2oqAmwyNVO+yQeqt69LZX5hbXpbSxo4G0YQ8Ay5S5SkgxlpTZgLdvGPaON9elKiVY
aqCdVKKC4digFUF5X+vERAFiQuxpwpUCRAYlDxQDYCXrm84tIxf3nNat0l9ih12b83o5NA6oGrer
sQYIDFTfzlKe60wphsZt4qOiUMkHcwUATyj4Pm+BfbhSPc01+VMNcYXMjKG9euPx4LvMwcBKzgod
tlqxYLTfdxZ/YwNVEXxHeJZH7/h/EAXzHWN0Cv+DFJ0n2I9ZGwy3wkPjo04IEb7wtWSJtoeMCF+N
/zLbnFJF7pUUBqYoz8Hvv4Slhz/ZEuQAoXW+Q8xCuDWdcio0p8htz2TTOtqA4sv7vNHCf3s1HlM/
sbFJSBhi5QOh5CdhSFLzbMoQcSSlUKla9pIzj50TQ4k03R278BkIVvIzbuV3skuZ1gw6dlJt3STd
56Md34/w7DNerjmgGtkvfm+lXSWi24VtILi+FYWVL3KaCD3UBChK4HBLPCY2lA/1t6vnr4DZPBh4
c3CFalxxL2k9pRZ5U+BxgxBnTnsMswRakOkDmdd7rKmY0DjNiziv6Zu4K/DfmQmX1To0zGL3ysWR
SdAt1LH0ipIbkY9/EEyJUcbPMgbuXSgMMpvQhDkjVJ7mvliSy7xLY+roTa225dw5NXLTjvhdKdsJ
cls4n39R1qrl7hL6/rwEAML8yvdPCk9ZjTzS5kaqWXu5Q041nPeKe09en2pnsM9IgIPiQt44vZxp
13Lpu31w3XNpU4+ETWPK74hYGHyWdEfB4f5A62FbnHImO6FXXZ4qiYMCYGGLm0dKuY3j4eg0qNJk
lc8raaVbqhMWQzY55nmbNl7iZoZYKQiYtwC2+pyFFyJBtbmyljoKAaaCoqtGWBSbWMfrdOXiL0g5
aoP4tTcHTinymQ4pX6LetqFldtsdZJ1BBipNHDyJYujtfg/4G/XZSqKxybuPoHkMPwqw/VqsDPBE
O79yM0za2n4JfLAQeli+SpvEaZY1yv/9fuyitXNVAPDpCZmjAmnB3l5MQexPACghD35J/xKd+7LW
r7bqVD1FY15BBzHlg8VbOg0GssSCqfH9kcT9yCJ6wQXlDPn8v1Kjh6yXA3r8dHK2Snt4uyhZYxjF
o9oI/zAx8UgcclbnmpdQNexfFo/ltAK8SdpV9RQyX1XpoTeHShjiogTrK8vH2uVGRkbY8707SrHr
qXYXnPWmzL2vUYptSk9glbgxfbtbDMvIVEJRLxKaku/G4S6O8P1Xd+KL35MsJ1IyeUfJYNoEHNsi
1mmG5zSJrvi2sX5K68s6lAPifO/LdqjQqqa/NaK6gNR/kLO0WlyRe7+cSl4VwEDl2rDOJtbNP4WD
NdwZlCsnw/MTopLVE3aPlwxvOcQSRUQDpSQruD70SieBV7n5BEya74VLTnXJKe+CE9P9eLNw3Rtp
F/LgzUBXVsr+Fj2uWYdK6MW+Gc5X58rstQI4auuRi+P1bJ3F7PizKQTbgE1RBgegvnm/BPIO24oY
/tc81tzcfy+vSEdO0Nvp7lgUqshpzg9RJ/FYZNTe2vy7gYH5uyv8K7fh4UjfBJcyOPlTm79gJien
AmhcmVeaNSvhRd5AQM8Il6gCAUr2zgvHtFSYmRoBhp/2bntOLuUr6yNGZHqbEcR/w3yM3C79eoQp
2pN+oTkQ/ajMtOdL4KOlFQV7qDvtgEuLJrtF4rKi3BGH7LogeQxg60z/alMcrdbfDAp03QdL1FRR
lOTd22uy+n9MMSR1vFStFPM6dTxzv7c0CkXHuLmjV7u0363IDxuiKgfDaVIRCa79Rlo/961qz6LP
OM0T0mzNSS5krxuOpBv1V0hIvYOunMEbUrcNQscPVifjL0gbaDBKViCgRt5N+0b6sERTN7+GXwjM
rgcQm1BNjgr7DiNPaDZO50LMZP14bS2t+1M0YU7PVp4i7R2CiBNBhXW0YM/6+cXxCwSI5f2qW3rN
VV80EwejkWpuvtkdJfEOMcy8/L55btpKPZAs4C5gULJoxTVva4Cr3tgy2B4PJIH0T/+E5xbOJJEi
kcIvrS64vNqQqv4OOb4UZLMmZT54TBRXgzbViOvzHdFPejfex4X0GBBU6EOJYckLLw3ebJ4Vmh/f
gVATFYwaq3l3Q0VciJdJbZEliPnH/w/Vxe6O6mfTI0/kNKZsq8rjidbU/cfbiMAgkQHeZDP/o6Zj
G2BNkLN3UUUiLzmArzDuSH8dgEeXGWhSPLxH46opn9dYdXG3+yvw1k/1kAyY6qzORo4giRgTeTW9
2nNSBUeqqnqlD/dCWNnkNa+3Uy64dqfv2g0pnM4TxSpr7BZIJbthrObuSIFshUAzuK+xTdaXanEj
Wj7pIoFAAGxJCX+vD6BQpQmLEHaPKURDiEqUluBBNlCvfbUpsWn88sCPDVarKNK37jyIhGya5pFX
HuoMTwuXcxO1RLsyuCN3tty1ZcrA60Mc+gqC1SOyULGkDwxB3xV6IAM1SAdreOXZc6/gDYZKzvVq
Qi1uHAT/bZ9C71GWh2EIqCsyj/2bRNMZgs7BmEURym+cbSGHUM6rEIJkJjN7yjahxJJEKt0h40cL
jzPV5fyp+aTraswD4WJetuVGTLMgwXerGIusuAoYpp9T9Tw9P18918PdWt4CtekFJQkgMB86ANrT
e0hb5k6i9n+SlpN6u0qZdvZUH2fw8iTqRixNfUxjxQ9MbSkMpS6b1eFcUKwkasUrWNX8P7FqJxwX
juNDE1dJmcJsOXYjjSCLK4RTWN3PZNqNsjPFl6QPlem0ln8siCoYryDzTmJdnujsqAaKYRfSf3UC
wQAzK7tzADZqz7HpgbOXpX1PggJNtQVE+EkqL9xOHwWXBf6ELlgbTWo85z2rt6IHkFabbwMM7zet
azqAlM/tbO8tbwNcsclHfYw9BZZ1Q11lH2bXW7fxo8FiNDm1GOP/22GAxvWzOdwscxO/EhpPNau3
HlsbI7kLpvI2cJp6vFxU8fqbHDV/SI+SQEd7rys0A056V6OjTY962PilCAtxcdezgAeZ31EYBfrD
mte60RtHP6KkPWvRK9zfXLOdQDrWdBettS48/P6GazUIOF/Qb/SMu138l9e1TT1x9XiqlB3jqQoL
1enSu4ErHMvRv/pvfNlTMr3azu0cC9grcnOFsK1EFEEiZQxEbrcLwM+lksgFBOwq2X5syH5MiaCi
bM0hM487A730WYwlvvGwgTUvUV+oTE8famr+QIQbIGoNQzN9WW4rMduF5hwSkv4RQ1SIdQFJoHfZ
nMqHsrIBF42Dl6axOu0TqcAFrJFoM8vOkwszdCBaLGl06QGKQ/8dwUSWe1+oUQq1kpHESEK0NHFr
+RUgihp8TzvWp06tI4yHk/mODrIMA3RxV4yV3HU+UD7ueuUHTrBqt+rwSvcTEepVrT0kUsztF6UG
osoXQ824rN0CN69Zy2uzhdwYiiD+lxt9R55eVCksL0MJ1P0vf9U2+l/8qbF9lTawN1vOC7x+0pRv
rAEZSeKx3KYodyZV61iF5n8KpxUqhgPHUdURGddCzGaIMT1gug/OFpx0NVKLAE4952HexTLo0ACd
2d3wJsquhhYw58kGINJ9BgknH+lfV/IKHsufhYZz9zDBsl0/C+lMjVGhHADc/Gfr5NJO9I6C57kj
3ll5FhGNBHS0wsiCCpARf0WD97Vh1Z/bySSyI63wGuAUdeoeGZi81ewhaGuTTFy4gqtSaNTvxc0w
OKHGpgAr1Ghcq0KtXFozxvy0ZjIq3MGDgKtx+g6e6U++1EwOEu/zaHq7uU8PIi06bPpSVqoDjpNX
2hR0hkfTWFBndtF09EayYhL7TXBV59zn5b+mDOj8GCRDcRsUFCo9/C62mIDVHfMppnJv2UNYgo+G
D1ghxC1DROq6lInkvyH02va123YbLk/vGyJuDFz+RWLVSyZmOKFObqi5Yvea9RpVUwTI6XpP6GQl
ePhW1Ata2iSA8jjej1oldOXjRH3dO5+dyN4iIKiMtmNlx9OeaBqP0vdXNZmlGFgz08Xu13E8I4B0
fUb504zvgMrnTjleadaFPkK4q0fP3L6YVYf+kDtAvh7/VMlO2I7ut4nYjRT3c096F0q+f2GcKsWf
X8T5Qq8ZU+0eOZ7r08x4Dp2RkkFiv6JS8Kn6Qu7JCLV44trifwOsdE3n5kv1jJ/iHTRd5SmzjwdN
SfE6phUYOiu+NdVe1CGUveQ2waLOHMBxESoFn/rzbOvfBNqCHXrgh/kPoN7CR5aun8X2Ufs02BQe
RuKaWD9s8ilSIVSnmgptXyqY0ygw7/Hm0Ucscvby81pq+arHTi+vG4X5AqITRQhPDKYbh3/rhDiU
2nqI8M4sr9+64WLZqjtzw/vybrHcaBhwQfZEhAPuL52BF13zHmd5zTHxNILPNUhTe59wfmsZONrt
Wcxk2far5S13Pwpn9AX2PUhJr54csJJpTll2Ioh6M+MAi4uT5Wa2hES1OLaPN+dld9oEN7NEnt4C
8+QzYE895gNUpPCuXAtPAxgqH+xccVxyWf/yt1Qed0+Cn/Tu94arCTW6ssFgWJp3XQMGDfb2wzcx
4YGMxtXG4+np9gVIcGyTKcowM05u31au1XfdI5RW0iR6q/r61BcNOofEq9bsWFpzOQiqE3boy7Bi
eYeycM0ShG5qollUzWdLCLBJAYaDyFZWkux20/MhU9rcPb08Qtvzoeyg6O3KH7nzsf7TgD1UcPhg
/AbF7RfHGlwKM1kcBxfq943/oqIYkQRcQYIkfqTa6dwChuRuDMiQbWIRFsP2QxU0ebR25a2pp1CL
CVvSwkpxGNZXHfp2J0BFsJG9e9T4/C3tWTeCWqUbbDTnWQ0AOC2OQVC06uAvjPX1+XotBJ3k5oYe
aRiRDPiXTTtqOghLpMrOhCsI/LDI8CI1fmHfE1rGW5hPw1gcKaq58v+/V7XcN2onL8uazQqgxPZQ
Oyt3Zz6MnlZxaK7w7ho9fkhPfl8NqaK0YRltNYv8JbryEMlD0BIwSmJmylKX+OXDmt3sr3kKbiSt
7ufYFeGLChWSt4r2HzH4tElYnFhdTesAoi/LtgguNl4hE+TXG1GQAnT3UDNBKuPTo0AzXSD6VuQ7
tOZFSczceNsmWV6bl6JmfgLgkRo9AWAYUJGVB2kRxpWQ9Pnaavza22cvjHQtQcY5iB+W7CqpAjZv
H2qvmozksyhfmziljwbcF8FCaq8MiDlVm2/ZY66qIuqj/b+DHXRE28+O62n9LpV+4R2p3WCTQxnQ
iiRbikWHSRDybGUQeju43Gildj8vv6iNENDcRCzy84o7EZTSFDmUV74He+lK0yZiSRDsXS6iOHiF
Wjyk5lOPqE80PKj1UYuP2ioOruOk/WZitEIAEmiigAdmIaaIoj2N4762MLIOPkMr1Xsw2ZddgmuE
dF/hp46dOfIt4lZQCa1uP18N9uSTKEQ7Tzw34vVPnuKRa2fQiao3BzwRxa4yLkH6el2E8uWLH7FH
QCZTv5Z0DAi3XJtsXOV9Vd6KCMEVPFj/8I4I+NbqGrlP3nq5P3/WVnODkWTLopw2BSHLwxpTjY8Y
UkCIUPEco2Z3yQIWywUtGcg4Uq4QJBAFKd70a2zjKFBS1NttV5Wg+B5whXEwJnP5y0IqwEwqrCjS
X9jct5D5pZIh5TTJCracti0L7/Q12in7H5mlucbi0e+sgiZ8wsdv9Z0QcomJcUTWeLu1U9XR8pKn
DeXRMDLP7G7L7/oWWKHQsnkb0IX4UQBfdJN3K75qPrNnduhfsFpyIWJPaOJthsI/EqYX60BVFJGj
fm54jY9jEjE1RcTqLbURC7cloq4g6mnEzdUFN3hIUnWxahOZWWOCZCKgc+Zwi22TsUTcaadLsgBp
TwNYODRHfwG+YfJvNissl8yxH3OlFC4/cFQuxKOGj9h3XJ4W+jQ0shQ3IhEHrZrzxRppMi994px7
Rkqg4nWL6MffvoFL7RoBgrZ2O1wQIVeETo5deBJHwBdXpMuHhm8+dbFVNqRYgElXsri3OXlZdOTU
XTgaxdoMZVOPzhiO28KQE12iHS/Wzk0+0nEhudTcX2mPfxHtEddEl/3HP8dMVCuFaJm4qisxEhCS
v5I2AUTWjEkuuxweYpYu6lpqpmf962jLs//75v25AlV76xvzU7fgsgp6QoTjcgIRVztaX4ktJ4HW
z8vaJn/RF/zGvIFPq4tFD8ccO/Pqi2YPV9e0DQpiSg1z0MsdgBJMISdjYngvxq19KNhQ4xyzD9wv
0G5YcLXgqJksiGuxcxtdg+k2TfseLbEmAXLBx9lFyhYEF447i/eb+tFCrk6XC5FFph5HVIa2ap6m
D8m7hQ8aWumHOvZk3aJw0tHKudQy3g4YXnAhjBw600g/Ez+Jv7ZxiCWj/WhQLAO4r7a6qp1vhoyc
zTmg6pgfp2POB8DWkZoBUy9/AGE0/XLXpw1mnv3x1jzVZKkSyACZP8nNfmytsStimF5nNg6fedAG
milELZMHFRcp/x9mMgpGr19RIMxv/zoVMQ3z3h1B0w2tYPm5IGMEewDq8FR3nIhIvYVyLo10IOAq
IpbsMiSWPhZ74uaEDbIdDVpG/C2Vw6LDqXNlTI7arrMEfF19j0Qy9snoDM6JEYx9k/qcJIy7j/GJ
iKfKQg6MJxZ/iVSuBZpvGkxF8yY8Ayt75Cwm1KVcQVD82YNqMuz84EGEF5rxptS7cUPjuNefPbOH
1ceAnbqGoSDIUUWU807naeFunPm3NXzhMRhXi+Ix2T8dEQoPyZqhTS1kkagxCwnauUYULgtQVNUV
emSTnEq//24B8QwypKfqODuBXQU3vygbQPMFgZ8bj6+xmGtK6vMg1wGwtzmmhEFv6AsIJOO374WG
Amw97pKvPhoCGfjXyZ5yexbmdSqLCYjkBaEAZ2V6QgUMSl7kqfxggXE5BOJNuw5cE7Llk3OIx01d
TiQs9NlN3dBStbMljRAIrynuFuvXENIYrqmjQJ0e8M48G+juHSsacWbYj+uUTG9/jzOvGahbS3O1
KAcNcUKlPbv7SFZWOv9Ge95o96Cs86ppCdaAsFEvtbblCAwW6twZW6O1NhFONA86tcx7dnNDi/PN
qC0NUvfIA1xjJ9P5Yvon4SS7+hVeFCMvGzd917eQgycCxJJjbv+K4PgffbPDoXvE8+zvQc92O0N/
AxZdN3kdIH+m0Wi16bjmK+Ns7BJbVN393giyGjyM/bM5bLGY+LRPTCsjYRYLWO5IhBm1i69zpfD8
mIOqEXEJUFZXWyR2W6X1lqA+M9krK7h5FdeF3Yhu5DJzYye78Ivw1NYoVy5kCAIVXUF3xZSYak0O
G9e0prJJ3aOvX8ydv215EYvd6p+w0E2HHbVevwalf32KO4uN86UmhIYG7Wo/itmjPeOKQKrOKX+L
1+Sr0uKTM2+hwg4pFoWEYgW2SVARsfTyUfJxxwcpsrIYELRv8zGIVagqVpYHgd7b54tykiOZHMMB
OJTsqAQqMhZ6Cz7AW283/kCE4rYe9RqqSeH1PDaKXEWgDnW2JiJLK8BZXfl0txMHuPJNw1GgQCAn
W6nzu/Ze4Yft0ApuDk315IpjN7x1nojDM1xOdQo1ilSQF1J6JkRV0sxGdXnMmxzD46fpGJDhMYWS
dgSzGRtmwTg01wOXwXVEt1LZYLFnkJYVL73+n8tc2dD53w/a63piDXEOxB84GG9wP7rfKa6+QPp9
N8qwmnhRQvKWUBAJBpdGu9xSNEiqiXAkw+Scq8IEjbd3Pz+k07b4Z8cy794cXeyW1vgPT4sV1jRY
0z1JZW2Ijv18CcuKZPue9CPCiyAgBFjFaduqszWEsIFwaFdWoR55qevFjIQQd1P+6sUYnzdRaOBy
z68YKnQNQLVyyEBw0uubGfy+gDYnv27etL7IOT+r+PxAeFT6NrnkwxQrXnRz0ytMD4XK/M1gBWdc
f0QuKb+1h7YtCvFtFVDwv6XDma6LZfzAb4giNicA+YEiQ/K7VnbP4ey+Osx6VSfyNfS3FyFfubhG
DiWuLWO25+4MzF8wcLFGsIzZal69cVwtMbA00jlnnQoBM6dcabbbHL+TqQ/ywRwBWm/jrchxpqc2
fQxZ6EK6+EGgWaqB+7zKCF9h4cJaI/tp7JtQwKD1uGh3XFe89d1eC71wG76TetU9pQBpOW81GjDk
VM59oqiWzozRLZ4EhvjVZSPdAPNCwdLWMAnMke8UeNssXNS1gC1pPs9kSm/HhtIqRrMdS2HuCdgE
9BjaLAszi7oj4KpfXvyFqZjgWPkzBqQWsjFgMRfoULqZTpYMWAGbjvL1RNFgKcnxQ4k+53sUyJvQ
e9WUIgTrK3+LFXXBdpncotL1sF8oGaEQmywI35NeYcv1yKus1PSQjFL/E+rr4bCp6oEd8993XbrM
dtD/BQZyOVHqfTCBl6FO78gxrPugzmrzg1oAWFM1FYuHLK1ogwEhrKSV9fcFjBof8dGryMfvYeHb
+dFu5ch5IFIb8vhrzwGggNialATiniA1c0pDJf+2iSoVkYr16egC8oygSHovmryQuhgXBOb2kpRO
GxpEICdR2NELrE8onyFVjxiARJHn3ehwSVEGnF+P1+1aZ6P28AUb4YCDZ2JglmW7ymUOHNuO1iab
Qv74vrA+AdVHbThigsasAwrtjN7A63EeDn6qBFY/Bn2JKIrNP4WWiKa91GFCXndRxJO+Edzn2o/Z
qJxO+h2Y1q5nXhUfLSAx+0daaE3CGaIGdcMQzAFotQogM9ne8n+KGXcSKp6WwSwxiluTEUeJjjtd
NCJrjVJf4+LVvmSrq2AePlZZOCpVzIJDM2vinng0E5NZ642fVrJH8BrW47V7ZRK/rvulIuC82fe1
H91jVDTQZlTW/qe3zKItIxrsjCfvFqFKr7zmu3UBTVSdets6Pww4qkwtDOycg6/LaLJ4++3yDxKy
2+f3osP7ZSOkuHmXTAwNPUkpGO2QuoSaXJ4Z7tP3O0ExAm0WKWDCoEIt2egE4FhN+ZVL0i5IhUQm
2H9Lb/yTq8ESFTiZmHEgrPFam0wWeoD9Q7BsTDEdgKeQQuSrFwGOBIZurJ+uPNeJtvtXQQW1zpFO
BxqUkvxSIw7Slj85NLTLvPaWTazGQjLuEVTRT3jJ7eFsYsH3iCNpZlpBcXLuvQPAelagZ00dOlAb
LzwxdW0hltqvMd27xFvI3b+jweJORzUUogO2Xo/kY+WryO0NanWaBcRtZSwz/2I2/AZHcU+kU5Rj
SngD7cfLG4aZRMoOVc9GpmMoge7HKeW7vBEGSvdvGNYyBjYLGUbDzaKIP5dwpk2xHMr6lP2+Qees
W47S1vvyNzw+wQSmdha4N3bL0JpCZcoHimyrC8SUOEIn3H4Y6+sngJ68XNCI75k9PFpdrpbROWqX
ZnhDoxTKXDZf+a34ff1EERRWzNm7hQO8aNvGuzmPXeyHwteUhoWEIUC1MlKnZ4NaUp0SKqe7bfnF
u6XA7aOELPBrRfo1hec0u5GLT6jEhi+y2Dr2yt+TJPJmy0w9+rFopWaJGJGdsA85kuDjKVK5ZPIm
hAFYKaLnf9um3bzmP9PYsWkEMWsv+rPQItqkh03Ay/ekqCdJh1f8rTyjkIemmqd4FaWT+O11MVbV
hC52GhoszHTeEv+VRFLbmoDUo4JPgCHeHS0ZmixRUgRiLFLcBfPJaKzfVQ6DXrRROSLqMMkZF/iZ
cLJOab28XnXxNWsnWk80wkhLwuYHLOH7+7wLzAAK7lFdGE5NWeyF1DcqGqWW3ajmHNAStwtUo8Y8
9YzMbbe5WbxnfpD/ceQxZF2nkCfljqyQYmUkF2hOreFZcLbnvoo2YGDDmaS1LD5cB9EinJGlqIyI
emZZ6gNgQFK1c9AunxO2sVPyMGL2QoVvGV4dNUdPNEKkVFgCMSATJehU/KI45rZhrJlRjwPEiL6Y
Nrr1fFEWaXKtYKib4xu6yNRuB6rV/j65WvDxWMsBALBK4swZdnD2wh6rpRKd2cFOm8jr1YTZWCWp
yCv9nP/Sd1Xq4Xb/YUa4If5M4muYYBR7SSGHjchMo8JhCIN1csbF+Hnm/4PzLumQk1ZYhL0wfu5A
kAnjZEWD8Bx+jREuh0vXizjXr814Mai+n03mmSXj41ZOMLncZi7rQQRyygG1589Q6AG9Te6g/LAc
2yqRy5jgCikPb/Wu4/Kk4RI628yrmtwV/BzP4DUJRPTVYEckr6p3pl7bUEzB8eWp7pzB9kPpH0ZL
pJySCie1uSHJ7GjxR6v7mTw6bjv1bONebq/So+H5X7iTWM4U8d9gxjhnftibt4jGRyY2IxiQuAfQ
Rz+b97wnc99UHMtcaSPLJS9aXRkO8k1QMQI7L/o04XzftT9LoHtGVSyEWRzq0vuQgsa58mLUz1tp
w6abYJLaYRX7kf5qDhKr83qdCdFRw4OOOR4Uy7lO0A6qX/lD7R6NeImxbvJpZsDDx+A83dIjRXa2
bqLqzAOANAdaJoB7fxtJDX694/JENjPVbx4X8+6vR4vHj5l1htV/3eCxONNuv/F9RIJXrI+yEL3o
sLvFhJ3PlOCC37b5AuSUGQgKcEKXzpMmdEKVEatTeffTWEQ3bE5gvobVNQE2rXutdANZcgXTwxJJ
s8qIxP1r4vf5o+aD4qvfgUFBPsUAnIFfYjXKFbPXLh+5RsyuSO6vSmsYqKRrbYxMxoI3+/COTKQW
FwyIIKBMpNmucDe7JYXuJs8SY7GeaGSTyLp4RBNlecqrI5B5YfGLME6qzXTK9E38UIenCngBqXqq
w9trPrwgUdqoCzO6k/HwRDkqowd/SEMx9gosqEk8emG6u3ijsLF4c+lgXnj7DIi9Dr00CjuDlW9j
OaHfcAeZWyTTJ/H43BQuSM/o4msdLVb96ux09IesZjCc02GlTF6HLOMXaD/A+obyzLyK6CMPxCH5
oj6MJFsXwIzvT3BfL8Hjl7XXgrQFYpxXpEnqwg/OwCX4nQXUyY1at2crC0qog3eH83gL2w3LSEaQ
XwhIjJK72Kg/7FW48zAZO6ESxt1I8tOLmcM1VnGGY068SGrlV+u/t80tXETNf4W/9UxaWVNhvR9z
6ECor6uY2jQJxxv+jWDRA4e8dp/vbV3xci7GGu65iS8VPXiyxuVAZ591zEs2V+CUEeMWGfJOLwF2
PNrZH7WGvVLiSzf+104a6eWkS8RfsCfXBgBNXDxh05N0WuptUy3WZD1Ion2A9oLhIFAGM5CulXAx
N7x8xePrmfAjq4Qe3bH+8CW6bWTJPi1U7414aFrz3tOWj9BFrMFkzrVGyxTD7rXhWkWzwOIpgIyL
CSC32yp0A9fAEqAC7koB5javV64moPJs3x8vfiZqXg93sPgJoNCFkrAV0VGf+fccdC7x8P33uzEo
n5i4OTVq+4qzJBud4M1LAsGamYTwavG2DkP2KnrY/6HvTQUlowkCsaPQU0JGQ7KtMgDF65ZxvQ3D
CaVtS/aOkycDVoyVhLQ0v9dV87Lj9vzNn2stxTDn/FzjZuUT7AL1TQmp0Yyo0Y1+RK5NzXwqo38Y
AM0q1wtJRGu/RgeuK7BL4y1ftUB4xyfavUC86setZIjEnZcjZpimRWpP3DcxPs6lENQewX3FcYQ/
Uc6pOcy/LeHZ9gIoIPnEUfQN8ZT9SIsk310FkNbRdB4xOcPcFJoRUL4QA4Y6qesh9l1cMSsvVXng
1+LgzWS9wqUwGKnN2O3B4L3KPzJjDho6aZ2sIyjjtPx5lE/kfgnrFHiElXpC+jst195xHMwhbS4u
s3OI6SnTBCQvuenAWpaukgW873y0X9OQBiqkKW8sX0asAu2+HnGDoLaBY1wOhAtMAOsxmxBKscDS
Ns2rE2gBq9vhBulan//21c7VRDgUf6WBhd6POLk5Cef8sKn/NZ8odwN10MwtfVd2tFi7pWJp52UK
hw7SUxfzPGML6WVuual2Dlo99NpZ4VYL1NLFDbLMIkuPB6gSy3oG4OskOIVGpKsrdRYLYnmVuyaZ
5HeMjso1OwdDzFTZEsEntvwZStwibl3q9FpY3ofB57ijVeoWnBMEjOiXjvLCM6ITKyk+A/1I8elu
jCkb7gD+a6/oQVhBmjKOYD1joPlP4Xtt57rBe1gBXNOowoDysTp9WQZWU0bbctoOY6b7TzGZ7n3G
2JQxjKeEfELNpuT8ry1svKjW3ZarhfL2TzE5WI7A8j5hiJIZGWoCRvNRJimdj3oC+bjA6gvLET+7
GRsKBNZPYcGv24rr/zjyoObiZl1LgsCr7y5ewzHSS5VHh+tUpyFYBtdACZGFnkb5FEpBeYyskIda
0wmhmNx6QSzoKkwPZa+lECBtOeeaSPZXYNtq/g9y83B9j81IkAtdnYRrPLKRXWSVlZh4r4iPh0kS
Xy0kvusc//aBLZnzOA3VNyrSifrBIvhDC9snjl3K6eqWjiSbKmRAy2YARWqe/ZXFI+lRwce95mOD
33YQXM4vL5tNK9S7/XSntq7TIZa2zc6hLRVPBWfkka8c5fWNeHFpNjkzu5o9QooX9uDGtZLteVxO
V2rQb9WKZ0tPw2b6Hcv2IrO1bWldyZmvexsUENdRgL7kB5mR496OGI3quLbuCXqWIeRv+YAVupt9
PEtww9jwsqjnApzrZD4SVIEckGGXqs1r4Q1kaXayAG1QFHhyblWXGM25e+T+EWsDOXYwkS4Uwj0l
f77ziWJunwtbfQezJvEOazrFOoPN+974FMP+3bNusv9fsQssM2trqSiTOBYKbkLCQFMnTDVLY3ys
PcDxLE3kuHikXFtrH/ajUgEOuPdEeKOcmqPc96KyxszGVXiicF1+fSRNwqmVzAJvenJGVWzEKYEp
s6UNd1yHbQbfkYdcCDXjbH5Gs/Mr/CPAO/YeQZYvYx5QsIBodz3C1dBrO8Y9i0aq9q7ebmWgwt0v
FZ4EUsYmX1RgQFgTHBRZUrk8IC59G5Xt+nv7lKDxYAL3T+MAyfe05R1Dm+o1h3/tSQIs0UuNfZI9
muMf4MZOEQUVDAL0MjecBoeozFn3SqdVH6FEb8aNIMl0qc+yJUZeMKxm5YGFnP4Fz1LvJzpAiKLb
EAG6pTOTu+BnYMaaA3fyXo1FRe8UKHbEgmw91m0jMnZgFqtTycuQNySW9g93ycxQ9RxbccJ8hot0
8h7b4bki6ubAyFZlD9HizIizKpzRoJ7sTH7meE1/ADq33W2x+l8Aw6QqawxvM3GDX8ABGQehnYSa
Ud/6uOnW/Y0W/LZ/b4zMDW22cVo8kceDpAQHps+HjDXpylJOropEMgAjCHOIkeef5tl8SYdirLvG
0SMjQMUm2Mgn3tST/S4xUYZn+5KtDS0fwICnQZg/Xle6y4fKHAAKRJbNBIiUibfzVl0NY9ReW+n4
PzYwjEovkbiZsEq8hlSqeakfZO9WKCa4mrL1UaK7svSbJ4c4n016QrPCFbHTj191xMmysmF7A5mw
b5ezSDVxjn0YQKfH9EEcuE8lNpdouy1pqQiWuEOu6qnS1CEwvQCIt8A3iHqrbnm5U38Hg2rhKIU/
Jr9/k94IP1KdtsPHUrgaPJXmrnLtT4C3PDBZ82bbN9E+eO+Q2RjMaMAq9nBmbDlQa8TkX2OaBRn5
g1q95Q1GmsFyz1DUGwMNgNcTKLUCMS/wmHCtTXkC2AEyWmkRlvzWG9QDQvPynrex0MSUyKBYZo0h
WIW0Yu9QaVCayEf8XZnEKAyLCr57qLSlBUq0GNyhcSTZTGELiBU8K4NsxnRMUanpEnk2ifAfzXZN
8fLb+eVdCBbT0j/SAg3IXNPJBtGHpeNHjuTpD51vHlQTCwN9RAh8vytzJRk5nySaBBaawsUI0wBl
IRDuwnzT9xAzmmps4xnilILZlHGlxUprlGr0TrjSxZmp38m3QtOsno2hH+RgO0qhqnIHJqqftRMk
d5jFs7Q2t1TPgKGmfX34c+TEn88u9o8jgZWEceEfBgXpAo+b/5SGcVR1T5HBEiF+LOWCi23cOAWH
pB8e2eihw8Ct9KxKhY2lhwxNpmhDqZQLO8IygobpZtSwZ1LmD7b+lPzBgj7SrwjJheTadp7IdiAW
LQxGhhDvMQh1WWVcJPOLt2mOab4Kzzd6FSob7iChuQBUVRPadQyaVsdI/LiME1fXgAgPJ/UUjXpV
BngefbSxKAFc4cOswHMjbqIGUhAnJnaOJfdR/i1kfE7QrvE/qgbiuRjAkV1Kcyq7rXb5NOs4oBF6
wEmLfbCuJk3PtvvVZRpekgkfDpx5uURJ8JSNWhrQHS+Uo7sQsZcxDz10zc2P22zC2JRIMhmxeh9P
GZ8uu/2Js39zQmXK0Ci/tcnd/q1LV2hKaubnFNhKdB3Nsoovbq414zkTEm2rsCz/SCKGmqYrdT7y
N+aE6thxo/s7EH8oG0NxiYWUpSGbhF6E1L1UA47oRdtWo7UABywFP6MHi24Fnds8b3zUFl0vHcxG
/PQmxX731pPBUakUyUMYxeRQLTCRI+rZhdJtaocvFhoEzN/khRtfeNcuASng+6D9fIBGM0+gNodN
fOEv/GbaxYm45ePzsbagBiJ2frXySZSWtOHv1CKV6f06O+vaFITacamufuqrT4/rdBH3vfz7Mjh8
wMKLJog9hD35pyZycWt29RcyOKG1vW9dR90BTI6g1eqYVoKlpMpnn/W9h075vU7vgDc2DAJjENHm
ry9kNlPfv7ECFPn2gI/udPFQhWFTOSiaUlyRX6YBhnkadwm11rQFvlQkeb/hvsw82hphZjFEGT50
VNDkDbXete9vJPr6O6vUZ0HKK7HpgrTIvHF6H4ZLkQQWOqmlyBSYBJnCsi0GWbYi5vzs6L15bLr4
5LlHayFPNTcRXqjtGDLo2jMuVjJqYu85wTSCwbeDDAmoip+Lh8NU0qHgua+iu+yYdRXezxOsbQlG
RsbFUzsQnnTY/ErPclqWjy1QaCCUFJQJw4aA4Q8R3CzbR/CsCJ788PrkGrtouPJtZvdmPSgTOKUn
wxRhAiRec3/mHD2rtuRMD7jSMqiu9MKhexbwZK1VlQHdQhy2y26KCrowqLPZIb85DWv+xx68qbrI
HWQDvMAQY6R/U1wtqESoV1Vbce7AFM0Nk9MJK4e0fVnAzZZUf8W7GQk+foB9dMiScb1yk/tfnevu
FknjWtlmU48LzYpn8BFqkQ7vRrXl9jZrMv6RXMTGz5hXtrDDR24d6mow6dtkHHuxFiMJcg1QZmoW
vyAR7WQVDJKgWsphbjFW7+msCSrmkp/wZP3eF6Ij++052VzeKTl3NFk4Sl0rZEpbqwHRW4k0IYz7
c2ax0SCdSRLhKXJOQRc+QfhAzOt6XrJdPrM31HzuLlE+ox+isHQUUEBHytxMrDqkN+QQdBJH2ino
GiZIsbsJTJuhYJ4xreaiIFSiqJupfXlK0KB3U6MgF5l9xDukacj8DTv2ewd0tHc5nrynwWpR+tmj
t5GIunJJi/SOgliXxMEO9l9AVOQXqFOvS86H/82QfK6ApQYxyEO4gSaPLZe6ErrSHJY3TmDWcflw
ehBmevsK8Dyqr9w/G1x59Etyj3/ouIbYEqFWQ9tq8YX2NMUkC4/cdxkRaJ9SEpsI0ZYlbwJIxepz
LphHp/RGywwZBPh6p//5bK+1LvA1xA/wB6PHAhgH82SiEqggvwuL92Zw0K2W/d3dUbQVebsWAbAH
UkkJ/XjTSjjEPIlI4AneWQCJPh0aGZG5wd183vY8cxhwbIx0zQj+c7zy7gmQmNoRNv83dNfJW5KD
sCqHEWCmK5Co9mrHDTxjGJSWIvwP4FHIkp2lc2AIwUjSu3y6/fITAM2Rkhedo/2EHQGMO683fH04
F8dkm7hA+3DtkP5ena4/QtSvglc0Fc9md02EkyDGGdXpQxwoKPvr5o90FdJ32qLns53pgAktHd4L
ChlMpwtPY65/S6nizPFgwbdL7rMw+FpRJUrDaCQ9LU7SmdYVxluh56LrqRnwt+HTZ9UrkyjCJD1r
0jtDqXYpNpO1KpASE+52Pt3IuD+uJuJVwAR7yOVzXBeG1nL3c8aknhIy4zaI2KAPQP6Olhu9uxuZ
avkn0H/n7vonk5l+eDd6l3MuItXHUvj+zmtd4QJaGPi0T6b0CIe8PPqJYoWEKpoM4aT4eFeaqueX
swlxdsOPtVlR4P/06Y8LtyTgueGDcryiXD1FIo32EOkK4EoDoWWMxRU65ReCSEOYunuGWzy9Ixlo
JzIspvzWsENpVEOjjlGd7e2Jz02x8Olu0wYxQPoNG8y1OG9gcUo9s0P8mFmIcWVGUeHhEtMswlqC
mtUv/NCahtaAVuu2lUcSEahYPRbHALneWJMqUGtpgjXi+dPiR583D3eXHlJPj8v7Hg/97px6hQLT
SeaezG9al1vbwT9wcD6u028N7eRN3+ohx/U2QgK6WM8theepWAU36n9+KdsGunwYbEA26GYWtU29
OavTfv386iG0yssC5RTSi3LRqW9WZCBI4zdI6Yep7a4AGuuHsZ27QP4+5QURWs4xFWKYTruVUIWA
4UzGxrseorCOv6lvEEJV8Wk7XRXJ2Ng4I+YnIrdqL+Trc9tK4vyFL63MOd6EdwhTTaxlLI/sDsdU
TrjmsVKyAH0K8oIzxbcNTw4DCMgjkDSMO+9x5OpW2tyspHtRwU28aqyNELQ4YqWYgBVuE1L6Hk7o
e/y3jsChs7xt/VS5FCLYPC6ArjAVJ++87NsSRomXJ/15mGnLL7JdsdGtvR/WFejSp19WTYVnTF/Y
I1JoSXt4jfxY/vzm1DeKcckl4gCQ1pBemQ9Sm2ZMI3w3ilnyRCdyP3I+r+KoUCMQrSChlhdwdT7k
EKzyhWgB9i9ggj9hNB+VzBr9h+PLNQSWv4/D8QhUue7qHDiSROdRYh4qjhzTZK/x2NRz38fVKapJ
Q4/20cg/a+9Jx87u4zKVO8lGyLiXeh4Mt9bviGcPqpY3GvrtI9llaGptJ5adH9H0GhZOo3TilcJu
4FcDSfAWbyTu88aX3L1J28KLBsvKC3jny88ZS63Lapqg2lypOt2zSKSuVyZCEqiODjlAiFMgwpCg
E7/afpg/GRR6ij+bsKp0DjVTSCP6w8Np+BMjaW3zcbv/IYcBBpJH/V0OrlXTQ/lsrc+0zWbK7OOE
XHlghQwKyAaLZv5XIMIORxbNzqsa8y+iMne5k5Bp+LuKq27KfnaBX7hpZmLwBuJ7yns5FhnrytyN
9Qpa7/LedOCfL96oCOZnMImP/fPxYURGWBe03/U3PL6wRAfAjOPJoPkjgCjLbzLFZMAj3fO7uVCQ
SCR32BmOG5rtncIP+JiuyuyWVLAjKnVKz64O0tF8PiQ1mj5Lp5nhMIuPRhPUkHRhubomjcFqEPFm
IlIqAff/foyr9KihNwmWJ1OhTRxySIjcbVdGGzC9qp3Q9t5PVTCn5K+GjBEVc4+PiXkRdju2gqdv
+uk7VrxOKVWDE218oZJnosyHs6Kap5dJVts3yhfhn+K8fr/D2ww7fLszCKlSlnJ7yxW89z2b++NK
uBeQ36FZFTB4joVLz5utcilzKfQtXqKkJGeBIcSXMo+nlYp2k5hX8SZAPPQs089/3DKwabZP2xl0
JOrsj0B7S9rFonPeuwPxz21uzTgCaO2PPB5Q9J6npbCE0WxZwFq3PgzprDeFKmbUE/S0jPX3Ybes
NWSM971qayIp8WchJfra+TEKpywtuNQI8yQUCSjGs4aCQgEcbZlZlG+F7DWNLvJgjW013Qrs3l7G
rfgxi4ZFpRaM2Au1S7UmC2Y7pHzRuILtYE94bpeLhm1GgpADdyalDty9OOavp1e7WIlmEP79yrYq
rL48BPRzIpfOV8UCHB9Ug27xKN+2PBk7uY8ip9goM77NI49Is8rfivcfyHbqw2nyrvZbyx58c23H
j5iekRpt8kbhBlEkdo2NOwnoT6Ep5THUvv48hEK7Anazw3BrvQHntmWiNvK+unKBs5Iunb9ze0jb
Ata3OjhbiwSdsrYONXDQ1FvP0FGX9DN3BtYf/qbVV0TCy6rTlwGgbtKgzympMpRbkfOqybSIDd+9
QCEHeXHfXKX/ZsRHXsTIRlFnoH0g62J+du1kJQ4LDtgx1QzTUTLsLCa2hXBGR+kFjaDeE0wQ5OoM
PN7wi8GqZ4f/agfuZth9cfKQwAg0KtajUh99KrScQciPAOGyW30AQ0RrHhM1aWuQfCGZqn2znvcy
UrzR3mYr+1c97c7aVhJtxZeUhsNMXAdFOpQTp3goNrV280bCK0FuC/Z8xbRtjcCSKFYwgaPBerJF
tplo49gqWeBDeKGXFTW8S1zmNZzHDZg0MWvpZ125zngRehoF2nKE8Qki5cdZ17uGsLUm38aykyPU
NLnmZCL8wxrt8fFsHN4Usig8e3DyO5uXWFswqsMBDkEg37fBKNHKyKMZeQeX75pH6IPJK0sLQD2c
fJ2pakZyZWx7OYSSN6noVLK/bA93KenQJtWRdLIcxsnuRFnYD+qjZRcQUVSU07rGkpK1axWedauV
Fux3lE39apayOpdaGLTrH5CneZn6uoSiDFME656bP313KqyRQt05jWzQHSrwnuszNeb+Ukw7gpQM
qovwOuW/Iqx/O6+WpyceUJc9kwFXcSuqhRIKum/IYvhJQtYJBVIuRN4AHdreQzMMbXFQPh2oClOl
il/5ebkFj85Tk8QltwFH5NZa8Z8ArkP+Sr/FOzdxWvstxCza1HIZVvQsNHCJBtDIxZljC/Z9YHiz
jadXTOToVS6cGkvj3w6dasIFWI3zwZxhGOHFhWZ0ToWk4PgPdv/7TcSfFz5aHFThrOIqG6ivmGdu
0l/MO+J0f5tcMz/woCuBQatVVJjin9+qrfCWiZNpVafLCGH4vEGOe/0SujYGuOyZWH4PPeciVr4h
+OaAXzW7HoPLzxBABJH9oBcxzqjA9v7vrf8Wnf/oLUGSG9zaeEKeNubHxUvCmZrjU/BtHLlhcBqZ
1JjttGenuRDZwrMyORKOQ+5RBpi+8qOJytwMyIlDQlTJ6wGCzYXDkedggBzjBvgpzFaxXrZ/+hhX
gzV7DF+Hne87tINufC0QI3V4hPwoU20WMxbdQq6xXbGNPp5ZTNSb2dXXSCGSiZcB74FxNab6TN37
iUe9yGKRK3PUL9Et0FjXg+Nt8KLkF/VC0PT8xBB5kXu2l1RKc8Mj17+yARHZ4gz3Jane3tqQJ0aO
jd0cXnDSen6eEQgvl17xx0TZ2Gx/+t7sRlO7vIFfvkvl7aPvH7ND7QNM9Zm04fg8b6RCV/uXmFMH
fY+9jhI+nMcoACjIHJUGc/QsCHB+7SkHzN0R19cmK7q3HedlyPMJi5GzXWFllBdDAn/fefq3fbUK
3XqheJybYhNIo3obQPpD48fzO68uYKhC5Rp9Ufkej9zXuLTrtVPzlaTRsaQ/oOnu2H25+2jIWB8k
8ZFGX+D42I3dMsVnp/aSS8+yGqdD5B5FSIKwxWNIMUzqRzR89Lk6sTsxK9hSUHZqOyTlULFy7TUi
a7gL1sxznrevRlYAjBmiS7JE+j5rHAcFCGwVf3x/9+THXmbE3XnGlvaVT5qDYBbPtkLEpaEhu6er
LTzhf1Igf7ZcJMJohx0QbisEEoI16HVGX40FEjC1Ys09HfaVNmq2WfRmapY4plsLFx4n8zZDeG5G
j0F0RaDhTWB3Jq1kF7T6skn6p2WePVIcEDGiidkL892ZiBeyrSozslrrM1xg2WUeRnSfscFiIRN1
r6pVPyRnjZdDoPernJ2WEXT3AR/8XX7/+HpdJTyPLYoGkV5cI8XDkBGv79vLab1a1wyhXrxGnFMq
/+2ARY5EvD/JgOJaP8A7l1UA1/C8YR4LqDDjinwvE0pFd6AYejzr4Wc/Jz6BmArht3Y19Baxn1Bw
27V7EfE+fgVc6GOboIN+Jh8iW7aCpfO5txQ/MPDAQiSv8Y3cjlUc2xT6apfEcbDOcb7cONdwH33y
w5ckf+uMqzjPkGaCIpA6B5wPzthqcDey6dzlfireyy4MNW+NsxeZWLSuy5E6lOALUbiIe1JIUhVv
wpR3EwP4x9oEyH/Q9d+uAl+8uAYdp//Lk2PFvOldZsC8TwnOUJB9owdY5vmWMdHxJg4WiZl9hddT
HwPLTEs2HdeMIZw4IBjBKIvBwz+S8Kn4ak2D5WtrVe0wF797dlNkZNHOQGZAbpCknL+AvdY0H2D+
sx8PsxqbE3BGlgGfMjwfFx+VQvlzktrws5hPevSFccNKfbOMaS8Y+JLdXv+v77je9gOJWS2UVvn0
3rtfvcpovIm4/WOpVPEaGXNe0ffSZQyHkUo5lkQZAPls5hWiHVl1VY+swhpukpdZFjZxIXQyB1KO
jjrjKvjzPw+2pxNtsXChrb7C+fiOJbRYOmAfYYofIOEhC4PLtwXRL8pm0c5QdLHTPtsC1xIi0gGy
H5ruZeoMMZ0pi3gH/X6wgr/fNTBNZyKVTypWtwaaPADOpzMDL8pZaqmS9z242sblZ+NYJG7bFxRz
cFYCKDyFxO+bWSiz0xkwjk2qcLtulsMb0d4m1VnHXrz3hIgRLAoEkt3NpszGaIDXRg0PwxgS0HWE
n7/bOMlfOGAPTkOFONeJEUyMjR3y9jwBA9aJ5Zpmxwhj13Oizzk1weXLMod+PUQx2mQsbdhd9mYu
wUV2P+M/5HKajeR/FrrOHdzLCFU+Wh+JmNsly558sxqc8Tn7ZCjtrTM1xeh9Va3SQGL8zjVRl4a7
CxhxmehnRREcHBne+6Nl9A2bjADCNQMR0qJQhu1snYNkKOuKp9ht+aWbd0di0vfNlZl+8mruze/3
NrU2ftX2Vw9sRbfqu2Wk2RD7yh47SE+KVLhTG/5yZo0tWvRZ1zJg2cIxHo6dnfPd3uGvpH74bEMX
hfKS+U5ru8b/qETp9CNp9rdtzk4cKHttLHdH3ogSP5N67BGBzCwejYEGJ2JXXA/RkVhiQuUGyBwt
F+IUQKaddnhgtyhwjYDPT+9MxohGRNF9IEbbbXEAPDS3DoyeK37bK9bbixp2kX3p2iqux6iOcEhM
7Cu7rH7ZDRm+sLL64nWRr268XzxQROJ/6RiVKEQgfK26Jiz2M2Hwy3zLV9/iZVRg4Pkllyp4mxGx
kRF0xX6a9xJbkK3/ct75rub2ahspfa2+KKLNhTNbYujPMxds55CEDItICusQgNl1LWFMBEmgRyrL
XJ/oH3JHXjWtbStG6OeZnyEYiqMvAZCI5IHMPCChYMSiDKHHfOkMd6rhXIzSKH3FnSEi8c+Czpyt
skEjKDvqqem4ymi7CxMcIVleX3ADkNRuxmwCpvKl1Ss0YQLIgFBj4QinR9PYA+yn5aJG6h36yxjb
oyV1GQ61KghAGJRBXRmIz1D/Rpyh5Fjekahy3dB75b+7nrxhKEbXimIV5Qg9sS5FmA22gWl7UTzg
eKG4Z77k2aqICUFa9xy1udxWhq5xL0zM4fWT5vjdl1d1DUd/LuGJQYB2JYyRIoprxZKRNA/+wZ+G
qS6wQdD2t31S7xGQK1eiVftxC17A8I9bK8dwGOcNV7XaAylFA75LJ+KF+FyE73ugrZ/EBBk1lAg1
6Hw1kTx4SjoD6wUz5P/k/Ucm+wNX/eoB6iJTjglsPgHcWvZ7r2TOZnA9V1imV6vt5akxwRr27vtU
Um7x0iuHzNUqJ2PodIiL3Q5hs1scf/4s+wIiYKOA6jm+w127QDzbfpoh1P3jAZ5sXhnW6q/xPpEJ
9tPhRkhhkV7DmNdW2FHS+61zeK7DyqOvM1XpVXhXQ/I+5L/Xv+/5diZbcGnFgGamAvL1Lq5Hve5L
HDoUrfig57CdKdUvkktnqyWrBvfQUxPUK78RKZaSl6Wjt4O1r7pa+L9yDlOGDRRcWO5foJqI0NL4
oyuGyggQCp9LyMvK1x/+qxZ5Hg2WaqMqNCF4fs4XcJTGnGMcxUm8N6MuUYuZA15iVyqLPxcxsl/k
c8bi5RwfzsssQcgrj9sv+5xBP9ZOD4oqsm4XBIsdrweXO+xDHBu9K3/5Vp4kbWGGIRI2k+AOUfVk
Wghu4ehznG5yzakSomLMxkZvPUKevM+Txl7DZNnaIDVzXQrN7LLZtcXaZpWSCm67vpYgh+P6CpOG
OqzUwXdlfGU3fdG+iSk1SQ2+IYVYRM+eQi8YYjFYGIJm7thmQ9jMeNUnkq1VB/Qy+we3hpdpzCWh
SZYgElCMnkAzNJpOv/MJIfIU7NObgqaHjgFGSX0pTvlhE+5vqNk7tiIKPATNbxZOWOOkQwlPsU0p
q7APXyVxn6ob0btKAYFBV4qMLlRrK9Uh0D2t373ot4OoMljVpGNqQOAt+NuhKhY5zyfGqm22U0eO
eGHk4mOZGjpLWJrsyzSSfFZcfbToSKdD1SF+JLtZTLNWAX+4Bo3OwvFc5WsZc2U0C75VQe/QRJ7F
jTCiJZ8DkzzsGZ6ipqeKgv5F3LCcW6MLUtBAdUMhimSJSyLCWJ36H2CDlBiA8m9hSzDfhGDZdGEs
4V2YGn1zbQ7fnWjSMx8wuQ4CUZfn1QQvgzOuz0Uvjos82YxSGAKOT2Qmd9iywPVcMiX90W2w12w3
at1+kU7m3ID/W5gx+xn3+cVWGsXU7gnwVE3aDzkvdmYAclywv8JhdkGAvGTZDwdEkIgAzhr/uE5O
sX8YkWkNTXmrUReqF7VP+7DFvSAdfUO4EIVnJ4jpJtfttOraP0y/dpLurcveScAj1gbT/qGZuutS
qF6FfpTEqbDTRQMH7A/ej2o5zTkV9m1KqHrVL9BD2eQdzyd+HT4/tw2A/eyT4PZIm5GpxTjJizK8
PShw1terKgu3SYuMujskM1kTwXkpNRA+PLcrfOkXEKvrZSAfZRLneRnxXVquLXTf8ME7CBd0ToVD
PdnMXyyM+0jvuTteaVg5F8OkZ6BuArbB2ALK9EbevUsjwc8c7O/+hCFYvU7A2rKcrIUHKFfi8NIR
qp4EvG+RFGJlFV3EagGVwP3gpt6H2H2QWxTPT64ayMKVaPkVqRHQ1qH9azCd357CcmZBf2DQHgu5
wOq74NJog8+is87WzJfz8VOPJJOc9/0ttO72/XbDQYnd32zyd6yvgjaWbsFdvwijj6WunJLjFzex
ch+1JooxuCdWuxzOqmBHpNnPWhc/JSKOxaLykQveAdeouR806PDc+oqtE4vDmmKwi4To32RFlRGn
SZwgelV1lgTACXANDp1269utDJ4J5alTdrbwtBt4LwjO4rEkDkWC5fIBBQAu9I98N0i27ojDNvL4
O6FiivG9hqGfFJAszbu6jaaBCkb2HK5FE38eSczn6LuE2GeF/G/1DGYaAHdJ5pWNv2zi6nx+1ZQq
kHnK5btdPC54PY4iQU1ro7oPFCzRS/ZYQag8Yey+0U2kFI6+jGlSbws8HE+1rUIWOgfzzZmwaS30
Sz6NNYZNkeaW60dxPbrIkjBtXSAbM3aeK+zm8gpoiEnvZ7Bs+VnUGOPoxOrplA3kKxWBOTEdB8bI
umjIwxLn0bQK024hZjUD7ZUlZDa3t9PXlSHQbEmi5Ph9AF03Cy2RFpx9ucKcIREvIW7RHpFJxR2d
ptbboWn2LKpcy/7bpTTf2ACZxCVbN/v9F7+wl6jKmVO0I7caEWmJjy0GTyg+IVh6tqGIow4i3fbG
Fjr7t8zKnkCh0/ovlRmqrJqiXyP66vz9nsvMpYbJ9r8UqXuyAfaSpHhbNQuHQTLBS/qh3lShRuRk
3kINQ8SrpBBh3RHdTq1D83kxKYJ+eRTRid87loy9/n3Jgfdt7skIdhB7cs1uXj7Y8JCtGaXt3Fpn
857Wh5KnmhaoeshUBi17MPK/j0cKYrmW5baONRCGAUA4NN7Q88mtLuINQnWEeieshusS7mQcn/FN
Lw97DQIjkpgI3HE3iOIyf8eA0F4oxExBS8PuvdBcBep/7g8uHrAI652f7Xfn2Ly7JDxQhJFPR3+U
EbfSu6rpBy7nE6D6ULb7ttq+OWpdfEBpRkfcD/5Ypaxfg6be71OJuwAzB07cKJv+rynzL/75BZLp
OO6hHmLhHb1BMW0tsXAZBYW6SGCMRzYz+av5PVcjRjd+LklOm08TIwuN+xiS+7ivPI3JScQm2/7x
+YU907l6Skl6DJC+Gw9RfFM4IxpYLxjW2zrluB1M+2a/unPJamR48sKVpHrUlt0GQ2niXhrzYdcq
VCu60MBAQd9n5KnJUmFbsVaAklcdXINBZW2L/JNRv1ul9EcYAK18avljgcZ325VTiQaR38Iug4IG
WT6RvqK8UwqX2kYx6IOMOcQwLJghUDhD1zReT/jYJPnzLN8K1wfavJjR6ht+wj8qG9cYP0f8kRGP
+G9f3hKQdW/7LqyZNNsdWXgZTt1voYqU3HyMzyHuE53CQ61z6LKCOuk9JOBNhWY4BPugZq73IA4f
HvydH6PwtkDAChQopos9CupfJNgLuYXje3MWRoS8bNUoUbAOgWffcMTDv38B760JHzppgPtAigIV
IfOEbgyNxmid/up/TR6NQOVgQ1Z5lcsewtMmC6a8Pu3sqiEmgK/+VDIJSS4dzPodTPyP1WR4YlDB
jCiT+mxV3S5sRlEpQqjxSOexikOEUEqHX3Dhd9w6PcbHb0+YXm1WaScSeFZ1eZaaVd+YNNoK362H
pJGnsyxPrkHvrqHiuGN29IuQ2ng8kmGNzqGXgd6EwftCGj7lB3F7sflS8mpQH2ZicrlSYXQEL24Z
xZTAwLVZDfPVyK1ZtELs2EiWgsrIlX3+g9RqG52gHHXbEgbh0yfCbKQ8NsJ9lzJEUAFlD1kdSeat
hvGpl2mYjZJqIpFzl+H+oxC7MOfZwSTxhU+1VfZ//cOe0EO34b5bCbxVhRlMm6dnKtfNSzhMknzm
NRVplPQjWgoWkcw4kYoirGcpedpK0JgstTmdUHGV/YrAjsT4mLoTKEmXSz5+0vYEWXjQoPZQB0+x
XAeOk6MLyT+GnBan63VouUpYZboOU7bnyWVr47nxrbk1kHU8Tsj8+8qj7NxWGQJzEbQVlHTGqR/o
zaBaMcNgXTbDGMo+UrgF1kANI0l20Up+Uw9y0BNhV9RslMqgpxCWUFpxMllMKDn5+zms0UcI5pEC
sacbD9QFcClD9z8hSVLmcZWq1focj3i7q5sQCsbEEyqS3ihYQx4efIeZVlCDNiPgBLRpLEuE2JDh
cgdYWcG+IphKn2MLd00/vuhV8e7be7ZdOC2xbs4CL+DOPhN5cKpZLmPSIw02bRMEDdx8j98pVadZ
u8jTceC1OkBdTBMghZEENmHBa96oWrejA7D4ZqLlwX2BQoaUF5GcNsvXutvA31PmDTIjn8iYtlR7
oxMxUyou4S+MSI8/RqpdBRom9ulq4i4h5LPfH4P97WBLZ0q40QBjM1DWratnaVknNxCUqObIZOZ3
hIXNhSVRIhVq7ugoFGmdTmchIVMxbvUal379KEriFh8MtTgJ2yOic3yyfjOLGhJJAjMWL2bmdTcm
RWRWaI3D7JTG5iUlqsgmF+Ajd6GppL4SqMu5Q05ZX3NXhLr/WQxQYtVowLD9nqJtgNUbwCAqcDSC
AYwxAbof3jJyJ7DoHLATqxdlKhLUMRH5tOBpTTw597bfAfYWkDnKUpGZ4Uueo7RqmXOsIBT+qC+j
9lhQitKph6nc37kCDL3UP7AoZ9a9OYMFtO2krXjzKpAYyDRVfyCsMu1AaWzTPbVnJnIZvUCfWBYV
xGQZjgA1Aq7v6WH0oRpEk5ir28gvZ2u/+CHoT/9Y3nPAzpU8aFBPReBPsuufztK0s158khVootL6
G4B2CBWiCi6SFRPrYooy8m1K83gVceeobWiI9SXsAY1OukAkiXudbGPYtH5j9oqeJbxVakck40N7
lHShmsvwwtpLRwZKKTMb0XopeAJZVmjUjWnt/K153X1AmhLYwYzZ/7ccUzY1ITtNEal7pfUa3HY/
2I0QSznLQO4fC6IfK5LpV1muWSyQUAGBj/YfFixuQ+UBXGlEkLJpTx5rlEYwwCvU+iB75puhp+0m
hqiVJukQyu57pyYU6AdQId429OtlPUuogQIxmj2ArbnI0hLD7Nju2YNanVzUZkCTJ+GG2H9B/GyC
bxqVHy0L7bP4rqS2bF6ilZ6Vx424yjMARl6LFo0OohC+VJV83Aum3r7t28JxReu2X0ZBrhkVMMGH
O/xoPC5bBnO5bmWdWJBYEucUltci+Fz0xL/rYyxxpGif15RyoGp+CEuKKZqzFhhDRlIGI9lz1kig
Csc9/D6IAsE0jqgZmPrBkPownBwq9vbSBjINDy11xpYOci/gBnctuZ0OCm0GtSYfdHlmbX6kmvWu
viWpXR3MyIjbAFlqs9OtjazE20sgKk48tMZfsmKKPtPCTOfMuoH4YEviPEm77dyQePq1VQxXK9MD
mKALSYJd2c3lmQhYXdvRNdq77LuvpT2XH3rNcim+baEpHicghVmWgywOugbtHtMLzz4EHvItNKT+
VI3hK64xTbbXcBYyxDoBzZv+WLcWy3TnHksZ4RbJzkvCUtVddRACPiE7TvTiPvI5Gk+r2gRh8fvz
qo1YL1l19GKxk65i/LdSMP4CDcJ1nVyWNi00sPGJMXqA01qHORUYKQ3bRpI3KXt+o+c5ySRRvHAv
/QYQIhPRlhVAPyFhNclRb6mKA4nmXlJQ74ue5jM655rk5Otqi3vbSn/FUAcYoMYsk3TLv6+IiRXz
u5MQk2ESa1aGMJt8/PhTmNdOXk6jvjBSdxwesfTXYmhDlE8Px5fJNOJ5AgK14Kpsflkl7sw5JGoP
x95grs0nwVkgklEPpCImwzE8uSG4Dnbmft0oRD8F1RHAP9tkYfk5cexc0eQ/AQQUusC0+9FxzhJB
r6QkciSrUDeV8kPwFC6FOy27U/Sfd0BWg3zt2lR44L+gagYQeu76ca9aUZZUNLFZ8Tn96s2asRD9
3ttTNB3CWg6obT1oW9ANlUuY8tJ9/ltacZRytNMEH5dC4wL6ejHW4p2mJCEj9u5yJ8iDtRyM9ImT
KeQ15y6vM8A1YDdb+Hxtlj/zEj4xZ8AMZpxzPrAVyu5hGsIQArXGyqBtO8eHzWXLOV5IJkrQ9rfJ
L0zy0bD6UYNOZ9A0agAPkg9lC6Y1wWJTHaZvqlKnQJqjE026n8qmpaqSgExU3V5fdZVFRx9sODw9
/o3cFAag+G8/ZV++9YpPehgy33XE8ZI3kt98S+2wvRYWt1bmvmeWDNjXbr7Pk5iXraNqsZabdA5i
BiIaqWWHu/EW7H4XHi+XKd715P/YIA/pue0X12ykHcsRPzMbrY4jZ8Vypy12hlgL9RMfcjE0/DdG
OL1cIT3sElYmrv1dKzDp304xApRNrGkRWs2pDXP+tDvDF8vte4hdMjkNMt/JRthkWV6hqV5GrY5D
z+sL8Gn2OiaMxrr9VOoiObkiUIVv8PsX++s1Sqjy/n5AMo78J3CPe+YwnZm9erGTqwmHL75vyIzm
QFzcE1YQ3qhA3UTuhzHzY0iKjn4eIVh+CX8VMm3BABa/P+/awxMQfLhuRMgr4N1aePPgMSfr0w0A
CddwwTl8oGgZlJBtOnvVB+K9nwaXSr53BS3kme+MCIoxBF7xR91BU9oRz1V8WZRy5Fik/ZdRYuul
qRcAy0/b8iUivA6E61l/yUBZenOUJ62Lt/A8ieG2/uNNXUfDgIdIUswpYxuVjzMOt3tfl6fPE6+s
z8SMTNhh1oZzC4mr3y4Y86Y+ZM/UsESncBs/CRDohLssg3bMxXGLKLSUZAZ9+/vBDBOr8ylYDyMG
Us6tS8pTyhQTbAMlDifWfp0xzIzmfh074+8z85PEKmoyBwXgJJR7M9egHRzBI/UtYwkEaZikdp+k
6bg8P4oAh/OcLrO4pefDROiE/zK1qwi/ZBDJ7qLcUJLx5V5BpXGTAmhvtsFbuNByMbwHnrFIr445
Hc+4lV+bfu03KD0WQwhnvk5Eg23cWa4DT4axjLsvhBTJ7JeJoshzK33OTH38tFn7O7pO8jYEm6Dj
FjeS+ZLhKckevy6v+aUGNDm2G4ls3a+UT6V9PtkKB5HQEKe8XlGmCep0bcFiZFJJex7FRStQEXz7
ox1rMuiQsCtkKZ4eF8EsB02KOJgT5OA1o9K9mRV8DnKehLSGZaXoBPjNKsBYNCJ6ts/gIxuFn/1D
LFkvZPIlbEE39Uaj1UYOMe8PtTgEHlvBAaXC7kX/rNNPLwKNa7t1eh3nlGCdvzswT1ArQs42n8tI
ifwpP2drG949jwzEFGRPyJ3e8+6vCx4+gJKu3tCwcJEfee9C76hreFoAUhJQBJRNa/lZcgnGKruV
uZuZ0x8SQswVbDuIdMUZ1IXqfuYt7BL6h7rJW7inzlhtKOxJPIobQOVxChOa59XmykmI557XJb4n
9/jguBjPaiNyB5fxlLGAxtNGulorXfkR+mhkfWtKHnKF6/g2aus0lQ+Y/ODIVHLzsbT3Q2NE6/jC
tXBxWIU8zRcEP9jO8imnp/haQJU+MtszhnG/h+v70A8QMZiVVBvcvR5h1zCXdKcNaPXDG2VPCtIs
SyHoFThqRDt8id6oBhQ5AA4BTgANwls5cUjdxEAJzwiwJuZIQJy7yw0lcvtS7MNg0yDNKKo0whkr
lv/tF19IOWu30UJhCullDSGOFus9QiWUABNiY8duesAbupQfc5cwdWeGhpkKuHgxKRvLQ5L50+DU
qnv1JOa2OWJcNJW5S111wllrBZ5gIGHH7YIQ/9HD2MNYIh0OaA2Bz25hS4AhZlBFwoM1+7o0RUX2
PNFZrR3iR+8gxgJ2SAw1Q/pDX+0sJxALBJd/bGESdU6nvTM3bG5ScIAgnZB6a3ippFATQpPQ2qTg
+yCz2WoYLi0/z5VsjvtxjzTlyMEdXf4Iq9gnOuPx+D5C95xDxPhgF9HUI5pUa8auDX+s06coEvmd
J/lbBs045Kgfv/+E9Cz5hHIb8gSpiI4Eo1P8ZxvsO7E46YE5m+3h7ontc90x0LPV9JDEOBO4W0SZ
E1iY7bSROuntB/C/eoe/EriXYOZKYFAfr6V/L/0t0uR+HsUQbnjXxwA5k46EkQZHqgpl+g1+nI+c
IPCXPg8D4ihsuXa/rZ77gC7unbLGsZvOZAOflc2PcLxLv6TbuSTFJ6qxK7mGZTlPdaDDenMM+BMu
DBOUGkLP3N61F+UnQ/5LuwSay24VEL33ZBIVHL1rBrGS74BbJ68GS/BLInXj88Fx+cpWMFr5tx1c
vleFuN1Ix4PgXTRYduX3aCnfxtDHMkk3nlH7voT0DhXNZm9k9ZzNBrqWz7W+laZGT4gDdRmuxb/O
XiKnkCi51MrDi1EWP9zGbUcVYjbCqn0C6cgC0y1dZXj6HJc0uKDrrp32MQSZ9Nv+KznGCDxrfQ1a
CQMIDkuoHpqTK2LOgCDwPmfOMmm8GMpXkvW1MbmQyk5pvQAt/fpuQrEQjEGzM+r6Q182hVI0YTy2
SoJn5dYMa8Ul4ct9lhF1bV0kz9bsgJamk+UcwdUZZxAERYKx2t7VCI9ttEYHNGqUuxnn5lpINOf/
gHPyR+nCkx0f+CwOFGiTXWnZ1bGTZBCHENlPb9rPCq+0hKUza06cg+sDRlPSUngqYjydChUKTIaU
dYLUMveR5/sks3XHO7niID9Vytd7Rttodg0+iXEGWTfoyN+/6Jm2UQG438zuPQVN3Ak1UWmRba35
gbx6LanvwbfeMV2LjNaHKZJaFExLfp45TkIS4CD4jHMYG1az+XezT5pmV3i1V+IgrB6034LxblYT
ktuUzL1QOgz0hwb6zbITyD3qfGryEbonpKuBYzwVVSzLASH/dXVzPDawl/akHj/TxGObOE1ViXyR
qF7/0lmrq61TGn8tu3ieEL/Fcb14rUOyo6kqvln9CPBcEYio71MpYO5KbBO5tNYJ5s/0D3JYXy4c
3KCWB0QnEAQZLKVAtRNh5suJIkXNUteg+Cov4Vz87RLJv0awGnR/GyFTsHZFyUd1/kGCjMuHQfda
P4KJ/L48Mnhsxx4JNJyxJPESHVv3ywhep1xgJClbb2TW7vsiW9zrRG5tCGAKEznoZzUM/2VC3vDa
8M73+Al0rXyIsM4QlQmDSld1oZ1MAN88cOpTDXMyzVge35JyU5bBSWmWoFg40MVmnvnAVT/adwQ/
migMfFGRZae7Rbg74ut8Bw2hc11YIDIH1dCcmOThW0tClDaxLyWeB6hMK8LNXDV5hwN5XvHVcrU0
f+hFipNCWRpWwlipu4iM/thYSeft/AqIOvR5cFpZF2P/a5NFMx4AXQ71vOXO+EJlRsMn70Yk5AVp
yLvoDUQA/ga092kxT+EVUS1UhMqw61uV1JUSOba28oX/vtDBZnw+pQ33+2GL9ICCd6gYn6rGryAF
+jQL6IqxkL7GceS6YvFb1sgAmujCveUnRHksIjX+XtDbul3MBlcMuc5nne9wrRbDM6f2ClrklX8q
6u+IF8UXNFZQClmFDpFuIIZyIOXGl5/gYvLsiqlGU/s6UXhLJmUT7+pvUDd/2Ijk6yHZIrYe9AXb
PyqZYB9byx0qN+WTjbyact0pmNCFNaxC8ZRyPGBPIigdHoehNcCx1hhxWtKqoKKwl88dH0eZp76M
GUnPlKb6o+EIwPSsPtEvtC3QG0W6wydQwTMhAZjwEL5+kah5lq841ugQtA179ahrkPeIi7KlNxtd
LYURjK1NfvwHmRxVkgE2pCp7vdMoe4caHJvrRftOEFbWOBTxCTV5CPScYAQplFvqzbP46QjjcYjy
Kcm9+U8QH3JGnJJo4HqjwAVKlsVIQIPfouN0gp2AhjRL2GcBo8mv0q6cp+2i+P4eAi560iBaR1TD
JjmX7SjEJWMZOU674C2EhLy5tGJYnp+QucEo2Hy+/zFVW1H0AAcHHJf+ITAwcMJ/SAcJMgyj5jFk
LDZ9SNMB1jstXrzoCK645XsfvzCCaIvCZfq6Z3typY11GQA02CBk7mpXP5CehUqrjN+XhSnlU9hQ
diM0C8riyrpAL44RIf7rpkXToFv2SARXYjX5DIei8bjADs7SSMg2C++PaQdAenttBOGtIZKhxQ4v
AfsjXZJXyCRkcbuR3rfSQmHL9IvJSdpbeDSm0LwA0qBm1Nzm2cHR9A0N3jxHQrfJz1y6bUq8P98A
DpJNMnfu8+oQe+frOnMmy9db4x75JfbTuupymLcs6k89ZCjzeTU6n4EYvbeXzOQszxNt+Go8sgrS
TYHqv7AfLB/0jMZmr2spqxmKo6kXZXEa/7syg7xs+zdP3JF3wOnwAwSiJxWk0rrFlptmny7VJ0d6
maUpez8wAOg9hYWVZCtzPmUMRYiD2gySJbrYJGa6elqfCskugBPoY7L9J6sI0SzoL3+DiyJEIJYY
wBGc1AB5vbWJyFEudYb/kjH/oxFXYbc+E3NbdXDC9mxt3CiUwmxROehEtOfKr6yALg3FNrqIUiWK
ClqnCD8mTKvxCQ2TC5iaj9Af5CCyg6JRM+E+PKNIFlWRszM3sLDNobK8AwtvHYRMo/uvYClU/htE
di0gE+gf3oQiKsq09r8O8YmBBgQw8YeW+pV5bUdQJKckI6Nlttk0wBsifH32NQDqD1SwZKZi4BDR
DidUAjqOhL/oOjJVmOadLNn+Kmn4c1Zl/EdQGGRW3b9YE2mrfh9D4W1wHmesy7ID5xwZ7v1ygKoB
ST+7WdzOqWomGC/SZf9kahOkejp/adk1iG+wqhdhfGWNWoKdIaWtxBeouGZ8gW9AbaEut8lLFGiq
CQSI271t7X+HAKrvOBENFJEIkkcpcBoLe6VmpOO5c8maGdEAr5V2JDE8nCQHa81fZoAVnhf5qKfr
L6po+MALXWnVS6cYde0LvDO8tmT3LkAmApCskLRRt5zQFoeacO/JQgvmFK1F/+P7TzQXoWz8N8t0
arEzh00Z9fjWKbByYp+UbCYvNlZ+Ge7daDw5eyaW2QYpeiyYRvY8lisMiOpHShk4QSwLR1knQKC0
nYdqnG2LzljTkw19i1xrji7Vd23FWI/hu4EUVNCBis0F+/y/CZA/BNPkORu+MsXfNVB2abdt0JwX
YyGTLWayrlqou4r6sT3QBN2ALrfTmOhc+A0gU6z9C0H4+ZHXhcdBRneh8X1NniQlrrrJcKJSqcF6
g47tbMh4na15KPYwGuG40BfyIrBipOXy2XjK8SLzRHu/TTi1TjJ1+GxGRg0UuJSrmTGxoPr/giCv
eMZ2adapDbW2b4D5Ej6Q5uNrnURRZbXwfSZEUta6EPtqr8sMCjRTKtQ3kcA/QsoZIPPtf6MLXWTj
ghWsOVXwxdrjFl3qBNkX8eRobE6+IXfY+hlrRX7MlAcDp6Tr2UhtAvQts0CTdBeie8lEcUdL9XhJ
gVySyDvLBiR0xrfGCO8XYVVchI9AnvnDvkfo94RYTiVLyB9JGzLUhL+7/Co6ysjRa4poLRsn4+qf
DiN5uwr+NMDJSdSxVfe2GZFntc3Hue000rRGPFTjapl77AsNJzcqtpRxVmQG2lzr5THWFMaQaOh4
8o96WZEJAWuOIX3Zpj26YuhFtCA46u71eCU0tyh1tx7YL9aVwAmMhEGsxVBmo4WP7mT8xKQPt2sS
42OPSPB+ldGdF8fpPmL/e7aT0Q39qD62xAW1bu49nyTsyfNiBTs/fE21+xH60iVRKl3MOwltL8SP
1HHyfs+gk8LuSuCCBBJfCR/nQHt+yXp6HxoJf2RR+AVOPqY+fLMju/rLRNJo05GfokcyShMujEZf
aGjOseJ5PXtPywb53BcvW5Fz6Z06RVtZt1XEAXY4nBMMY+nCkt6fXFeH5SjC3daekQ/HTHXyLdjS
Rgs+ldcgSXyOHoaqSyhUVHmFh+LdKzhtZw8g0UWTRQXaHamPprTnYyxUmnKjOmTVq+qlU5qC5yjc
Whvyh0XXu4c3L4uSOpD61GJZr8+JFsUHr88z9AMyebRybkDNGJMG5e6291XD4Yk2j8HzNuK00DFd
LudOxKupE3y7f6r4vQTCYqGWi3yE6HOFKWjUyYKzMQc9ttrSC/jwfq9pagxdlj7MloflcW2PS2cQ
q3ukZm6VpoxfTCxXbDZD9oDqMVRwugdvaPdidR454KVy7YRrUfyorhr+KSxddK8l7Tzp4Ljq+Qrw
mlpaQ1+Z7s5i6bE/9ltoM40+szUJEt+jVEMIZx/4BVrg1IG6Y3VO7lr/Kv1xsrUDNisS6g27oROc
Xzvs/Kq3uZedJhEeePt2D9Uzmg3ZpCBYkloXTHAlrS4ROYvbyp1Hh52BPQT1o+61OhFdOGrUSIVq
hnb+oGncHbsOzde/j43wkVJ6ph32dHVCgfNRzo/zzbE7flB/fYt9kUU3mX+k28+Z0yzs2Hyo9mDA
MpSLOZYbsYXr93gSmivo1kaZr/FOe2NzBnVAuZRZLLzruX/vEd1WQA1OPJrmL/U7Ky4AHkN7NdRN
3RQkRUbhFSOPVErufJsnIDtpot8klMqw18ub/h4x3aE37Scyk4bSuSLzMoTnSupX94tCiHKZNKG+
CWNLzGfoQfWkzKORz1MlJeFyoAQMnVs/+9qTbgQIskiPO7qWgH4le4p/hnrN/jujRIdFt5DZQZPq
yaNr6rMPbQ+oC3r4pMeKknfQRINM6nobDLx26UKrY/ZM6VUbh0btU9yEwT+lx6oSMuq4/vlYkToF
5u2ysQMBTs21GTAXxAC2VaF2IyMFqZ9syFvDTJktfZJNZ+Ydb43Cq4b1FUu6N9rY12ANA8+SvhFh
W8T0dz1O4RpV/1VO9uka23QBjeUglyJE+vNFfh1WeOXb/AbBskl4LGxPrCxnB393mLsPq2sLYmHa
sEZWlf/dxmXtuh99/isR//iFSU5OICtlF3feqEUF0d0xGAWcotHe5IH1m4j9eGVA0rml7TE3r/ED
zDXeuXDjh8rQO/mwswQ1OxqCbGfstCvUO0OSZAOTltIMcxKd0LCJpoZkCV7gau4LR9dkfS0qZmhX
/HeQEGYEObj78z0hmPFIzRrRYG71naQlxcnyByV09BsmfHBZqAm47kZucYaFN85+EnghIQ+9c+zO
Muy8WCsht5nxI0qOY/BK/mX6hRv9MfvjoZEAXoYAB1nZkfKogVzfV2ZEiaoBbeRppWefrq9AGDwU
YYob4I6FkV7QnDPFUdX4tlKIMucYzdV2hw4yoeZprsygCpQbzZm16P2iTpAYnpMcyZnTJDxmFszR
GQNgSDOVb8tmXhnZXzkm7XGkZeP3I7BCyf0JDvebnOdnKAOvyHHKB8e3UkLyoQpRpMOhe1j3svnR
TedNfLHJ+pjtTqZvyIJLa3sXzXEZ9LRQ7GPyDYv/Z+Q/bqg2arpWfpK+3lISR7mRPs61pfOYL8WG
lAJGecEZ/lntg566zhEUsiHK8qvSKBoZ8ABz7JIKC/r7Xh0kzZB7ae7VBC7NVXQuJ8lZCyLGWmhw
BAdoOHU5B2HWd1tisho+copl7aaLCQbZLdiCMnhNoYAvf0BfQXsWq+4HXQf/s/evT2JS31tiQboe
S3gqRlFenn1N8m6mVxDkzdrrElz/Q6dN2krptflgkr2zaKxJFh9TL1vbjmuxZfKSIVkDaU7sex6U
1A/4qbJf0Di9TFc2qak4/mN8HJAUTnNxaOukUDl2bCFs2r44CbhwtPrEu+pbaBMWa0lrLpzUpFoT
rUdKb5/EPsveb+UgG6VJgDRZ3SW515NqYIVoU4rmBKHEJY2uerTFFenU+wyuq0ySChSTypeLvR+X
SjXtF3BOhrpTyuYKYMjq9VB6sIpDcbr5+Vim+PFWr0k6NVf+FllPtR8hvrB52QmPPXeEwtAbScfS
glorUWV2b2cILYKTq4WFRh/n0bbzeCyQ1TxhPvCJmp1U4cOHqUoO33YeY3ge3nqQ+daluBEYTDvW
s0aAsJCgT+Z6+KpsTDYp720U8N+1vQiiJkegBm6pXKekyB2W4UMrCQWbbN5/P+TFrDx1qIhAjxJk
HuQJneLEMvRDWaffaszxkTRKZaAwQ3Vb9+xqlW8/VGAGXj//RTzXetDLvLTvzhgNhZFnI2/t+Mp3
Cf9bRLzVFcdc0vb9NIi9zVMAj/a8kaAHdzsINEeTgEcJrm8iFNbKmVCnyDeZgGUIqV7XzSxJDJT1
B+H1yq/DxmdJ02hs5BkRGm+SkpOhHT2mW99Uby76WJAOLPyUVbkDURO97iZsXDi/LqB/nC79e4fz
E8NAWfeDKmB2t+7rb3w5sefC+jPaEZKYT/9tiGIAgSieMhZ7+4GEue59giXXRwE+hW93fOg30w0r
5gyniB5WglWMoQ8062vS88/NlTvnnZRwd5ZWmPnhcU7s7nZXTyGxMP/aNTxsSoiw9juApb7eveo+
bBOjlZGRDfjrslBTu8HugUBaCYu5qYZhktrRt5mAU92gBEQu1yk57M/K+/3zRDJpGfdw5ScChXqP
KXD0SQT2jwKXktsbQKVMl0FsJ/DpDJ9n6A1oRC4r5TDnDvx5ti00S8JxB0UqvEOZudNy/WoX6562
L+u8MQdr4s07o1hX/t7ca+4ug9BwXwf+9lJita8CCtGCAprq0TmoY/jOSc3FAe2BzWZ3SzxzFcSL
gTxG3Mv4GSsSlvGqsiVgOrria4q61wbwfiTlHd+bhwdJCnOYvRZQxrmC6isP1A8TLno4QbPK4ge+
iKWK3Ei/buS5u8nUKVa8Fo3Yh1rrz+CmJ/8k8uXidCpx2bQ0/+6BkwRM3WqhbwBtlP3QOYxCvQW6
MqAkYZC4LPzI9RJRucWDg3jcwsHyM+17zQgvZ5f9sfYkQk5aGsri/9i1R6hsBIAhPXF2/12Wo7js
pmVOXQ8Oqt1UAlQMuYzWw1uMtN8zBpya4jiDxsQ9sR+4IcwIf6KMb9YmqLGt/gK8t2+/2+7ViwVy
+NN4uAV+VfpNbc1l5kH7jWgrEibL5yZ7z+Svi6fZ94Otd7Ij4/5tJmYF1qrQuOjahn1JBG7WVyBc
XSQELXfiYFzqvF9VIlvQsIFR+ybogljYO7WZFi5mdY42vUZTgAHAQNwTyxviOx9G+Kboo2K07iHJ
Z15GYKhyz6lcksuAty6bSaJNGaSrsOd6jCKuXxIua3c4MPzfG24J2tu9shgTosy2pH18UJlRUt8Q
ztT58G3aBSpPqvskhkOGuYPgvJlisITrDbtqvlENp+NUGmv/VG0847jX5QCeAWSP7OQOY5H2ThE5
M0xXf/YwQsVTnlaAGfufZvCtzvdu/ryhNlGmOcL8Q/vgTjtzH6rsgwtRcQ+/2z6grOSwT8rH0Ut5
cCaXpUaX1OfG2LXW3lLZVMI1SO2JXHAL2CI/WkdMQjdAD4t7EqIrOSqQyzsCBCOO6r6Wf7WVvVly
GD0KZma9KdvajigB89TPR0wSMYl0U7hPJQEYMkUDukiFene5AAoU/yBEEysfh3K8hvGSUGlxXIZq
OLJfgkzITPXUubkXCA9RwkjIZ9TChg8qVy7pv45E68qjDIAJL5wwSf47nNln13FtTxX6WhxFY3kt
YCR4IZtArv61YzNRDVCzAiRZgBWqnbQkSqxfErCwU/q4RaIR4YcRWc8ahSYCyGuUvzZmbn55Roit
yWHDBSQ85KfMmKrycWb3A0YC4YL7qGk6ud4YbOEJMu6HG/8LgI9vYvvoDoTH5/lDX1x7ZHsZaGTk
3AHgbrsd/BUguy2uhpK6+oD+sqXDFdoMJF6/L3d5XyFuBdc1RvPNT6RRj9J7ClPN+1Fk2TYfcKE+
Wi2hwOMdmOws0DIqdXH8+ujJwGlONWxUvtG73seNWc2/SN283/gVEXQXOgwKs1IvdgqIrmZvGr9w
29yqITuBXm9c1jgXwlQgl2G5/sMAxg0skvu8djZ88Z4R/HeR4qWEHl++xGHmaZdfH8QdkrG/gLo2
kaVB3KwRcyoTUN0E+K2yXewrJ6MLviYeOyGSx4J72qpvfhFQRWge9cOc4+717tbeMD/nnPMOMALJ
dgtSzpwFZasJhtxPvENcuuEYsGUt2YuoRlnfrH+ru5sr2uMqC5ARu2J+7a1anbJDx2cPP4GcTlXJ
eMzN9wgWPeF8Y6f2aZgV5qndjSlW5h9cApKfGzs3GKlXys2J9LugdB7KoZ8NOYmQM/HgfC7XFH4w
a5px2PIw9w59ZieQC4ZJwW7cuSNrssuSZGouJ11ET1MIoUOJtwYrZqJmmfJU3ZeTy3VhS3ojfcLl
p1Fd3zp8OX6VScFkg6KzwWSSi+ubxwXZ9jjGRuWwR91U0wP8nkx81VnLGc8Eh/WP9wsktqe1qV+l
Vw0wxocE7uJTjbwwnTsC/aHdOFMYBn+syMzT/TSaxv5GqimMZpvKnzBitKUavzqpMgwYysE41muT
fs9u1rbNtksIk1MySMbP3oAxFh64+2OS4CHqWdnxuOx4Vcb4M98TmjOrYtIOhJTqE+LrGnD0tow/
5STihPfYZqMfx3FErMtU8M3NOgmFIuhc3x13c2W1lPLYG9Er7/UdKPiLIFbiY7f7obwzpHtM3TUH
AXTBBFPcJKIZydHXP613NhPfVCENJnPUjDXECTyRn3GCUzFW0Uk972QkcL8Qu+Op7hUvs31KideH
WQtNwsaWh6Y/p2Jpi2/XsrjQTIjTDwRk+RriohOBRtPGvfnqvt7nHVfu6Ny1q6JDCepsyw+/t9du
1VGKZFKP/t2NLfpfQrW+7wpFGFbOkp8KRn/UdTZpvstltFLr9oFOFMGfWQLbRzYPTvAqho8jTckh
jXt6FY065YBZFUYvRsCRtJ7KgoEli62ChlH970ntBHoDcbE9rf2UHZ87VJoh0V5NarrwuOi6BvJa
aeXj+NiYu2ltYXjJxj/X50Gfju1FnPxVQRi3E/zklAqsL3xWLbhCquS6IR0y6pMa4CFnbJzShux3
XGmLzRvG6+bX4qWRAbDFA4CBMbVpiBC2LWLApblSq7KJUc+2rG+EnaW9O53Ajm/zXgDqNTsZNUnQ
ILATZkulWyWR2HGuD4oyK1QMosVzqreS+p7riyACZwzmP7cGKlNwUx8RB+tORI6E93Q+P4tKIX03
umTlOJ9OcsTfvTlluYVLV4908cLhiQwL3I79Sg6iT3q1klgvNtlAZqrGVgZ7/vYdDxmn4rLIS1YL
Oy23Dw/7FDXXhy5YTXsPqgTqoiR1HAv+c58rJ0Db1sKP+Mo/p1HTJzm5ph7m6AtEAn+j0r0ssGSk
Wfc8JDTz1rafzWGyCdRCFMPhHENs2P2a4Z2BaknGipw3KU1fdJjnBvUjqqTRsKYgjfHouyocjnsJ
xDhsT3XAPlwhvjuedAjsGF91bzcvNSlyFv1dCotMx2lvz3XSwKfOMlbWft+gufXwF/dM3/TgqAhn
PUR0+YSkhQasPkN60ebrOQx1QNRWSV3EszHmPkUjj2tQPJJnw35tkqRIUTj/dMp3hhW3/Nm1/EWd
dua4JZ7drRWUZoPnS5wcQo2F2N+sh3UaXm9iYeeLY1eTqipS+ianPjFChrIBqbp3b0Cf4UCNO3AC
Wjp+5mhi/RNhewZhliPS0rdVduZewJMvKt9UxthXZevMnrXT0YBfkNVZ9Dp1n44TgiXeRNQAVga4
2dLFoRTcbzAz6LtOzSl9Ia6SM3SY+Iyr6aRDVqwR2n59XuZUZ3/KdXjNl62NMwzhVgIv6L2s9fsZ
TKqhwYxGcwes3BjwQbWWvfj+1Kh8/Wq2NlBsdMq0z/qFfrojsPEA4Ms4Sjxw+DV5lrVNoVAUYc2M
duc1LFyiRyfqa6NJuHwpkVpUZj5J5uk0SWAHU9AlGkhcs62iVrkNB8EIvr1aV6YM5R7LZbIs27cX
WdtuQSJUPsC/ptk0/x6hWX9ZmVYPJ6/N0bcK5ck39PZ7KFxuTcsCRG0w3gIFpzlzd4jBLB3UNpPS
64LqbOHCeeZ9P/bvczIDChVL3hyYwAKKkR+9lkndVQTMObr8lYsicKGtpEq/W9jnH/ZXsRC48dUm
wVArrZwR38AhSlttkWPV5JsJykpJlfA3qCJMi/VgyI20tckj+7ofRY+cjbX7V1F4+JK7AtJ6lRQc
KqYuzLw9ap5+YAjaDd6H67cmejAHB4A6X2vk5tMt50RBxX7qk1eLSBVRaFKHhyl4M7ccgcEmOm5V
Hr2yS6ly4OtZiuTZkWhuMUKuS7i1kmYT/oMjjhToEhS8LavA7Y9+f3EwznWCWn3Ys2AgFbRV7S1G
QIvTCBKYyx4oQ3BVb53Hr9nABD1OcdulSX7lPbcoXi4wC6Y0NvZ/stuk7LgoRew6DRhbyKK761lP
u9BsfVzcWsEai+QkYJZdgw7PmD/ibrcCMYL/GZm9YTvJapwEQOHxAl9qR60lfqyZm0NKiHZ4dDDp
EyoKoD0IckwxyjFip0LkV/cGOFn1kiuSKqquUMr2p3BbArTAfjWF7v9aQqj+7NZ9Dz1NGdjelaWo
XXWx0UnbT4m1yKf4Wz+Fcs+5G42++lmIm6V/iMI5T8X/egEhjOLeYNJ77Rjd9f45f8sVRfwgieR+
ZE5wXWaJ5umVxHLIS8p3fyJ+RWsHVHW6c50a1R6gLjV/iFZr5pCvnjs+WPUYt/hvqNz4lm0QWbuW
prjXtRx2EcfiLJj4Dp7OULhCNx1tkkZMr6AL/oh8/xe2sNcAOW3HSJsotfVvlypCNtE7c4KMBzkK
jzE1nDSTEHo3IvXiVuHMQA3DYp1o/Cn7ijr7qNjWCHP7lWB1LfRN63HgH/5P3NCJVYJuN/lw3RnU
EC4xKMFqrvZJCZfPqVp/vqDGkKWYXm82at097XfEKyn+o4jlxhuNWpCWL9c6gmnfdNxOlVqoLxxD
ucc8Rs7zk/hzebGa2/4phlysM98K3yBBnrcuGEMv4SS7KAosbuSWV5nfdvsoyy79zFTp53z2OdYh
1ru40xr/efKY9ASWbrZMpczBcltbeWw6w/5elnZYJj4dNo4hNg4M+6oGEhB+jhHLj67pr9URjG7m
pzHvwRMIRvgQU5ful7HRrrnsdkVmrhY8t6wcFV8Ms8g8dYpvrIrTWmgw8SJDOuDBRqxmEYwcPNwa
GUipMiLkKS2zAz6KlRAd/tR8eu3KdlpEwNGkvELTGUrHK6YVMPNyoWwWMiQ3YgbT2Llfd0xV6Tfu
OMerlnzgPyQIoH02JY4jA6X5l7E2kbSinxAblY3V85FbVK7ETazF39XUJ354gedl1lqV4dOL7t5z
43SKGokviXjWcJrA+2pVLswHEALOTlVp8obOeqsd9H2M3KYbkL0u/Z3fMO9H5PweQgvUcJ8EIc17
59ieAehjddJisIu9QbunM+XRzdoP7bbbkDhzwq1LBiTrL9OQsAMh8heCunpNR1zo3QrZINusZwZd
RHAO+zJ6RALK9H5LXDSfhhK8ow9Esm0BR/ETB5xs7pBa8e0EdMye1M7mtWgqQLCd2iXklqjOGqRh
V4zDah1BT+52G74NC0vPUDm8QWqPs+b+GGqriZOq4b5i77m12DsOzLz0Z6bysPpP7yPLJoUMSVII
zFd/S5fP08WlJefBaKHGVdMR48L2dW+ddJ6de8AFWxAVRNfRPNrhlfkDtUpZhczEPgLVlC0MSEbI
AMLDR3NPt7Is+vTZ4jt+I3tbuckUV2vtYSoX6skoqKXVwgk7MUE63PFKuP/2mNy2jfEECsFTv+72
TYvS8K/IPXNE8T9gR4i1IDGpRKaNOl5tep5wZxD1H/c/ulfNzMd7pFSqR+cF+sb1pKH1/AUYcqkX
2IZatoD0M8dEhUInm9Rx3bv5sxR9DHQAYrLWzpJASOxEGBFe2R8rqD6VRxXvKXOqE1VeS2cg309i
LdJ7FYb7p1s/nUkIndMKj0AllCx7wlrYO6gcAa2otfLpt+bO/8fi2FfXDp+nTz+WbG7JvRW0h2gZ
CJi3ZfTNLsHYCwc//flHhh1O3Kjray16KRM9ROLJMck+TqDqc17vY8NCFLumKazRv2WH/Si7m+iD
RdqDauDU+8wxWiy0xSoK81xiFSpx+1VglKQHgn0doGtXaEo8JvxQokLBlcPj8rWXSpAEVgQNfVs7
ReqGgkxWEbHOY4M6/0DgOehWtduv/WNBttWUOmfDmpkycUhppKsgsPb5eGEzIbxDks9IMhBLBMEF
oMZwviG/6E4AjaLKVeJnxtTBMLPNrPD6yel6HcjM2fdxCmAmbOIT7utYAVRUpTwoTdTv/fXpObFu
059jIXgNDm50L2ZajQPAv4bX6zfNjczXg6wPyGY3b6gF0fmSVQx9UKXK4x3o9G/OWjDjOhgSrCri
orAjAT+JI7An/zqFhp7wDWsaZKrMXp7bXvbpObnXLQwC1stAmFzihBqwsSMxfbmiYKrkUxE8HTmW
qoV6YVhImk6Ea5Qgtz1bybm7jET2+7vP5P0LxlFjNZr+Ejdb+lSxeEtV0XB+OcKo57u3o5pJmshJ
RFRo0R0tVSijD5Zx7EzfqxCqT7Ejl7Gu3AVbZPn8z1Nd/aSHnAKz3SG0JYDvWCcsmI9G229GzQcp
83VdGQVmteS9BINBowbzxJOqNwFF7riPdH4Ha7mOSyevlYBnD0+qUCxNztrjEhLErJTG789Zjbzk
RHsgJ7pPEaNICHfA8ddGzI4tUFUaa7uDN22CPDyDG/9OysXcmTJ/GXXxji5+KK/QYA39n7jFHNoF
rP5aJH6TjHTQGdFPFsY6mu0F8m3FyRl4y/D9OSrOQwdy44w328fNwIv1cfXI0fv9ubYsKvcw8iMF
JVgLtYEbHMf9RhiGKxeTs4wK7N4eOGES20WfjippXqyTwuf1hMq/Ch5O47FxJIbZW3xYbHUJQnmF
FcUVtIyi37TpWfUJDcbCWTPiBfE3H/KOGAJSjiX9F1A+h5u1MhVgmqL8WNoysbhsRI347WlWVLp1
3Ej/vcVr2xWnpmAl45DOB/l94mDDrPikbrRa1uRKhEK36VvSuYj307DDxTboFJwD+FEl4eOmgXYC
PjSclALMTqh6eSJYHGGbBUGpQeEHFXEvqE4QKlYEAi01TVkESbTBDR1nuJd0TS+6h+Wnw6HUXfdT
Yap25bgVD7xba9df5YsdjSVxBNfY4J1m+kZFmfShUX3EnrztJk4LqdgUiHRby1a9EOi4c8gMsFAW
XmAtZXkXIZ6qwUtFYSwQcn9rEso5EvUbM0bHkx8ekndRm0GKMxXTfISwkUJx6aS7MC6breDcisJg
ZPyk6lpUJ58DOocQyyFrQN/ivxHLt5krWPDVZZ4W0bGvF0MgFY0tRqPm70f5nr0bdamAmkE2iFnL
GnArHy6dtSJJKbvDmy2HCeqeN77fZYM9mDRiJm3kkNPNIcfO8HnVvweuFKrsx33MEWHcrM26Zofm
ctaJa8gXUKXTRSm9oXg8AfyG6Hvfgkc1GOLLnHq0W0KXLer4IqGloPxSm9X85uw9trKVnnQ3P03e
8uNotQYGhsSnrNh4ke+BA7SgTyiyyg89hYni9qlPiBnYDhRjyavf1Q3iR9K+l1jI/ti/Jqs8x9cQ
VJbvoNtN8P8wJFVLd67SCKMrUxfRvKkPuCiYglhZ0NM0pPv4UlepGgXnzQ/mSHgqKffRn77APp48
3I1NPVtLElSt6I2yOIXyDQJU8zN15r9Fd43osjOxxImdX3vk4pkxjnLlvW3vhIFj0eXaGty92R0a
z51+rPXJg0GfIkrE1FL97PRGWmYhnVEfMNA+ZDjNo5j26OBxsHONNRWjSz0SqHEhd1UzwBZmEWnY
PHeZTVSLADNa5O99KFzBLwEjOFPSW5zuymzKpkccYybd0XjqeIZuAV6A86mvZKtDaOonf0tAIFjs
2V5L64SlYL0Q0UL5iNMzVE78NRmEnw/3IxzsV85rF7ev+xgpkYRdG1kPPqmJriIu1RWHU0QR8ekS
kbKBCgPu++Dx4bzREwpLB3emguwQHqtN1WTFKu1g93YcpstH5aRxnhnXGYp2Rv4BAQMMOrC0viX6
LHPuats5wQEX9/M5vJYtFGr7tTUuNO23Nj8/F09znRHWCcGGZpjzczuDW4+aW/QMidUeXAiGdKdG
HfpD6cIDouagah5IpE8AnrmrYm/vlUX0aJG/6vWNS55AmAXzh3YrDtwRn4ntQ1C023ZG0zOf727+
OCOOGXg4hjbdjd2jD2Quvi3+tvefMMP+yEtuVdv6ZbEIh69Q7umAmb59s/YRoh49QbqyWxGHzHd5
j4a2Y6UaM/iwq7x1XUInek6S30CIRHtTuwLl+kxdT4u+cpr10ixq8REW3bXKXzjSRl01uwVyA/lV
CqJxgiTtnp4/rC+0L+bKxGAdhTUQ5rAr7cTFAVfoGmtIr0Oq06G35irPFWkqslBTeMV5h7VoAOww
buSs6QN6Tbj6YGwa0mkui/JL2O9Rpdy0dux78Hfb0LtcsL/NULeQEPn9T8HeuogA2h9k+8vaUa5F
a5eqsOCGtVvR+CkRRgF1VMMOocTorC0iyJ4OT3dS80EfLvMqTnbBJnn43eItBucoPxNERenWGrM/
fo5hMt3hNUiViQ0fFj3e6TpDGo19Uv/8Y16Y+9xNJymbMK/K8Fw57CLyHjzoYDlOE8kat2/9DjNP
JM8csixKmcQqUKZ0sPUg/SEbeGH+cahrKXG+TB89kfvQK6VV2rnnaWsWYteD425IYk6kFr/VbWCi
EZySIfv+q8kv3jn2yGI3FfuS5jxH5b2P7nGPZblylJ4Y18g8rrAS1AHMfyFPtJb+xouhXiTkzkI2
cCh2h544W0DyUjMfuIjwgbDhuwArrqFkV0FIaYuaubxGFPBJJeLJmEu2r4hPzjdNTGScjbcQQ0VE
hLh7KDKifUUlw3AWnwXE0luv3Qb75NEOHMhQK/HSKX0FidB1K8p6TJMD604EE70Je+IFALFwxmdw
+AbAud/bb3OzrEIgjr3W7R89c0W55EFufZncenKlVHXk3kecm3GBSlughj2NeFIRYZiYjAlyphb7
qowpkY9y+aGI1Vm8HJ1PkL8ucFJa3EVZcntU5nLakdEUyDHGmIQra+lHglPM5BEXg0H7cfCB1YT4
1OEyVvsYqGpmCQhTl3wSp4HGfJr1iQsby+do7KdXSgN/ksI5LK+H1+5cn2O9ma3rcLNeHVDxemhY
a7WHIL12DXTK2D0w31S1ZAmBke21lvC2OFp2KagMK3eH2+3ERtkvn6ndnIwayaeJ8H4UIaviBWz6
e5MalfNfJLNG+vSPOVMuaTCOE76yTIL0kRZp06L7NXO8Ed7457Md0MIIUMzSCc3U5ZXSE1lCD5XJ
wwzbxPkvzPbZYlJ7gMKLRe/uGABjJZfW4qMS0zbn2VodzeoRMwMZQOS4NpBabyW1MtdSpO6h465+
f0SwzrohC+GxuE5ZiqK78aMmxhqVWxg/aYAqBbTYxlsJMTuSyuELfw3sLV1GMBOZyUAsFrnWAB4u
0alGLBHRYn+yDXHctAwJfZRHdu7Abx7JShs2QeE6qQm0RR8Mzo0v2dTWQR154OvJ98LvYYKZAdg7
U/d2nINBoV5aJWMfS+fLsqhWgCIsz6z6hxvUfQHprf3WBfmD7seAOpKWBdfiRcGkpGrtC5iHLxti
xCiZhxeh1g7RXP+tbmlulueZa2kriOIOIFYTGn2+uRA1p0m99+Wrm4siuJdBEZzxFznrpADyPJcg
qt2p+FoRH6erJuke/qc+JdO/nDc7z1pC/O0lc6sbDy8WxzmRLmBOpaX4Did1Z6gAoQge/QwUjdcT
IncFPWJPNJgRNTReXXfo0U1gPKRF+uqZ0Md1Qwh8tbQ9tbSGnWolq+/yKptRpcwPW3bd/rJ/isR3
DL/LRYxsoGKwtz/6hdU5UxAJlen0vWSVP0NkJy2o266iQp3XQnoDBXwaGWji9zkM0SDUu5526LJB
m60hgylbXVtfhgBH7Fak9BdOZAs8KsbFW4sWRzVbo+iF0HxikKt6GxLHvUNlUFnBPehaP8uOKauX
m3/avvlAhTTfbKEQmgYZH2A87l2ENhflGq0RVfr64Lz9FBz9Ws9DenBi6gxNfS//b+HqGnvIBJWY
0ShHLn+wslwV1B73zskzQy8RVqo/N2jIzMXXIsc2GEjjB5GZtH7BJLJeuSjuu1dP6ALO301GvcbE
77hYjud2liuJyuCUSVYfHPLUphVzh7J3O7G0hK7kSbV/DPbCMc9Sb6+FlGpG+8ru2g4uh/w7ia2E
kHOX6BN12HRrYw/eihDXI0KagMlx+0OAplCwwgRwh/AW0eEUujb01AUpnpejVWHyFE2PCTWDdaCD
j8C8GG/+6mVXGdF0W9+GCPKQtWnTmvJq8nsOIG93msqZB3CgifKY0AH+wQONrJQ/rVx8MrEukMTS
t+xwIKZ9LGFwN40eyoF/2TqpL1Yrx+L/t0eV5kqPU8lgCea/qb5GBwqth15G1T8zWVN0fiSUQhBr
e4sTXN/PthNPyXfOshiK/8x8TeN9EMCqwPB+1lLX8fw4SEIvGad0ZNj8ArDoSn2jAvAKC+AuFUTL
c3jU01cZZmaT9gvaGSwXNddhJIzgB7XOZb3uTlORekSzYPyxDk8AkaVynpPZv9GrcYHL7t1LZ4pj
Y89ZG7T1bzGtDI4/ncoLHwR1i4cPpXoRN1hKSER1lMdwRcRuoNGFbDcOOnXd0B2yX5RlUOqvfDMG
58DnrTSvEjfpVSm3O3IMNKJnbP12zv5A7WxzwE3mzc2VH4RU9gbSTxIj28+mtcFGT16p9b8FcOqy
opWkAw4F2iF1bcapO9I+qbWQJfwybermXl0WcgXRcFfSl9nRT1+y2EdYcBR+qDVufNnX61dialO/
r3yrAPcyvQMh17A6qYD0DuruQX2nK/V7R4QqA6l3+E465Vtslb8Sf7z+kwzQnYOB+7jokEGzY7lu
g3z3aWd/EeqT+H7UdDb53NUtAMvMtKMENm2uDCm4BsFbQZ75ddq7/7fNtaMMfnuPaF+a/jQliz8M
JAbpVhLG6p/qsMofcTTcsGFZuHlUuXXfb5tuQxsEbGHqrTL60fm2ZBZKPmYwNGS143cg52k39q1m
7cgG1QyHFHx7KUaZoCs2xAHgd5ezEuFxrHcJRuSAgZmYt835O8wl0e4UzmC1StR9MXvxgQeiSE0G
+8zFjfFMb589UvpVjp1bl++Jz3Fo4SxwKlTRBM7n30r5Sg/unwSA74eRhXQ1MpqjG4Un2hKjiS8x
Mnxd1Em4cdCdUF1JGHeMrAeyiCi5f723UV/gHGZ2FRvCmQqsgmwHLz2i3uXrkTuLX1/a1SUMmsoV
5RFquKj1kQ8rgBRoL8SXo0OpNaiiktRwhDy3vH/q/PCbE4AHiK2tls/fxJt+g2PjqmlksXwzmV5B
Oe+th0XFdRmxBbPxIdFC5jA2W26pUXF5RXDk2yto287qQCgNF7LpNiuaLrm5VBMensqM5usznnKK
vw7mgX5SUC/ppL4ZPUpJ/0/h5qe5YN+8t/411cVxWSMk2lJjIs7TFFuvewOIwqa0zVpdEk3C5gnt
+Hj7sM8XtQJA1OaShH/eFaDzoetW8qZDls4v1vGBdcTnVVgDp4gv8k8z3AXEsK6AjQ279BGqqU7X
i9qo4EJJHQhVXWYIPO2l1j3jqn/xthKmHvjwfUjhtELBH3ANFnzonHltWW7xCoe11pjjwNDg0x1G
k8MF0vVczcMCw+SXJBR7f0yOjSL6Be1s3L6YB2dYFPWZT38NJcKuh1VmOYTYV4PkWLfpd0SbY6wY
2s8LYDXdQtnHROrUVhQD8mhw13/hxyoJc5R/oSAbJcQ1eFc15lMjry0jndWLN/QEsC7p22b1qBzj
wMmU6P96U5U78DISJdU8V1F/xSAPEPw2S4NbeD6j/gv2GI/9BT2iS7DJ9YRfGKn5bQjlx9a+CREm
lZ86MyydXg39q+j0mCajBfeFlHTesfUj79GaPhTlCf3EaWJONb4HdmxkFDH3DCEe/d91KB6+uZEA
Yk9Gqa0BWY9wCop/ij4ljriTaFXA1a0ZhAyHL4b2KG6yUuidtYgK8yMM4zVy+RoWgGlisKsHJAcT
KYfKaOGhY8xdLh0Re/pwzt0M5e5s+b+j6QkktVaGMg4PoSjjN8/GZxtorzjzbyFbjWwbum1DDDPD
Unc9/ITFPFhk/AkfzxlGalT+J62j3QEB8hzbXLUbROC7ZIetmP2wJM/7K3b46kYtCxSb4rwTaT+N
QlVMkOl/DNYLKQZVVlVYc3+sZRRgQ9fXPOJ13y7iEL7oT97b/ODrcTaN/NJUMKW+V/TKu/qQeRba
yciNkEOvuu6EWSb7Iikxf9b10OQLnV5a929/mfiJ8thcKk4L2aOiFJDCUkZStIJzrFrli68z+tGk
tcszXQHYMQCfyjaTrLDrGFNd0JRNUu1LlcY2vCy0YSAxPjLegVIHidX+m4i72AvH0XaIIZSUHO/A
GmY1g2FAEttxlRfmj65atWxlQjplIMQa3GZyBXVGAPKbAWG2uc7594OToyOAs89P6ecMbmtpzllP
gH4DAlwVpoMT94+MZDYxE1reEZsQSiXKnltP8dTWMO2+hbP/DgDcFLm+Qp34RvB8Qe6ByAZhjY+j
HDnBJRaxw4XhqF4TopfNky2KYez1eQQf+PZ6IvZTzsTwLvnIvp/IyQlb1uKA8ruiSNtqI54u+y+k
t2suj98TPdiqnpKLk87dUr5aH/4IzPn89LGbO3J8oQwcu+9+vUQ8Hb0UJu0Ao4n47QY0GtWRoTyB
oJqZzGSDYys3TZvZx5j7aIRZzVtO03pxXc9PLQonp/u5StFriBnPIE4jF/t0/MWQhK8SHAqipp8D
SFRZ4z0X+MUTR6WzgkvjgKUlXRWiRfFCjmIXEioEnDwExpUzUo+pg6CMwrb0SOLJp41MxzpdkK84
0beQpWcEfqFCpXg9TS2Fh8mCgKMu72oFmnrbGwLBgYRT5AzBveaBVgQD4KYAWAAd0xhItZ2d0Uhp
olCSy1PfrB/9H1eW+eik51sqrpKYz/28KLlG1OCY3xW2D83bVW6xaAWoPNLuiCgSbf6v6Sw01Jq0
DpSr2vOQWrPtQAWaV42I/27UXpsvNuMQwgqJv/vLhhLh7Ing78OeEuX+bnAQiCza/O1blV7rR8fU
+EfskapcgYhudubpITxcuEfU+xERo7FjJWPsOiZ1HZ8EfCag0NsopVbAHDiXURULTFgNbMV9RNYy
4R9GRcv2dgo3hVShyzAssIwwyDOu4eb0I+K91Jjw91e2puSB4xv/Iy9Jl7MDjMS01w2+GgF3ux3I
QcwtkWUbrWPA3aedGL1Yu6Hn2W/itiP+pvQo0r2SvV49v9gVqwptQBlszfpxPfFMU4nJpw4uzMNo
jrnWCwlbWBYvCdLczxGCO8PoH8OqsSg0cOb4BxsMoeZBeccG4KF6Yw907nI038yxWsQRkTYWN1MU
2hv8mspKldkjcP88MrxxhuYQJvG8+rT8jPMfQELFbWTEpJOiFP/+IJYoZOXO7ktDGgz2zPUDaBnt
MDxV0boNj1fmQF9HodmtlN2gBnqFbkswJgKYCR2BcRhEuegGmVyYDyjUX0KNjl7RoVXARH060CDo
WzLrdIElRgU/IxDDtmX8g42QzXi5BYlT4f1TbaeNCQ0yyLNBg9B1j3UGF49O1/G0hOIPGl9qYLSx
VxgUghM23IDkkl/h1iOurA5YO/xq6zR+U1KsPENoqkNnE5QFqPfpLNHYoXvg1yJXLyVzmL1tw4BK
BaSVtqrykIeDSAYnrNlYM6KE8W1yay1qeC3JZpE22Wc+pBJX91YO0oL/G57lYgxOO+vSN7KNGWNu
wqKYfN795dFt0fF/sWKQlqhUiFXOd1+njwM182h/zPa9Ppmbj9qA5mTzDu4jWiYpga+/PfulwWa6
x+uVHyNuD9zU5ss9Hc3heYnPRwD03lwa5cSOPS4kLKDBsJPfMFWzSxRznISjz9NeSY3haYXRNkxc
RAkO+t8XDaieF0LjfRe5rKZ+8DyKXy0MnL117lEBnyUy2G9OpH+78AtDjJvmP4uzS9WLk48ce5un
sm0iMsWqz+T3ZFMAG/4QmjocN21gxCH3WeJAnJYItJH/4LMwkPW7DnTX5DWi8Sa7VywHe0+OW21G
uXkcdvw297RfXmwSIOxvV6zoJIHf2eU46JBrMN+oF38oYkbSYWgEdgUUntOg1gWlW61ra/wgrbLT
EQVuVcruNw114qYhzvmnbTyLnUFhvysExAyo9Y/B1Ibb42fTkELvFxJCqF1yUU56dm6ykTz26QN+
Jpm3boWPir/4fBYir6BdBcRAa2+835h/xJxFB35xQuTyaU3gG1oFLx/TVBPZN2/qJRZvWk3UFMPO
yhK1nD4r15V6i0DMk9URQgTXLTszBENL5AAKf4ga9Ldk7OFjmtPODAJ3/dp2aYUT8sAf5R5sBlrF
IcYkT7PmJFF59gOO+xnCigZUCuJjtuLb0U9pgg5i6Vv+TuSJJxBB2D9LDi8/rGrNS3Ft2A45gu3h
opIkjfa1W3g/cKN0mF6iEhERCtQR8tJEKgUAwqLM/3DE86GsfjRt7dMSJj8OT23vBNevgAsi2GdG
HGxljOyPkRcZfjApG/ODisXULLeEkyMdnFOqGEGbYW+qH5MsDdzxKU0hmDlbJOv0oM9xqYt76ufv
ejWp24JsR+XSE7rdc3Q3LcUksViUqC4C7iMlaoJAxQMbxhNfA5dZAfn4iRCgoSf0VVweSpxCideg
tL+UL6hN+a/usgg5oOy6k/VCZwuIvniyqY2DeZA9pO1hRiUbRKbvLfZire/PxDj1hlgqNyG6BZ9b
KAb1uD1vgwhHXW4jtGIE9a2W9a9AV/zuyF38ixpkJpz9wgiXPYHL3Wo0o+PNAfV3f5D9QcznoYeG
W8oumHj/YU6dEuElHBiuFVbPikWb/JZLXrcI7yxEyKemxKrcrWjFSt2lnLiy5BBaz+ytDKgFEbuP
/TPEw6xgIk1BSj6xocigQWF+Tp47TJaQgVxkPMailTZZxAsgQEdJ1vKWpFNcKkJ7Ra9UAXGekYw5
wFk1Mv6IZmKen3awq7CMKmFqEhyVS6niZRVuMZpTXrFJAJCdSJFZnLw5oV58rmInvF505CKQy+O/
fSS0Merqlj1jfXBnls+FYi/sXlcBVreZ/FGBSoAAxNCya/4qkpixiAzu+98hj28fV21jzF1/R+cx
rWqMpOZj9GXFeUmeE19Cc/llnKiXpzJmL3yjFB+U6Tc2d7B1QhG2k+bF1uxletkYK1jM6UPCOwfw
FUiJMUZpWMjA6xTzGQ+si2qapo5z55nyTVs64skFyNBWzsBp9kaVjA5ZM3wO1gFNXREAH+XFkl2V
ZQ/fe/4T0cV0JdqiZxTWNnPYArBtBXzWfW/XO7+n9uIh3xDU3AxtEO9L/W0xdPdYwM8ZpuNm8D70
+a0TVlxpNpRgZFkQIfQD39TMHlQFwErirUDYPUJIydwCbz8Nox+A0ExA+9+tVadeVIi4fv3545di
Iv4/9e5FG7PNuDESizZVU7NY4v3AKLACMzrMrwDYgKKGjczOSdtEBHNuD5Hx+VvAigfXVNc2oObW
nhQ56nrOtt2llXAbj5ujq0MbiVz7UChaV+dLq4uKddh8poD3mwV3pyb5ghgCFErU8ZCOrBoRgUtl
FHZcXFZoMYQPL1xSBgkFh0BNnZwPu8uWMqKd5td8VwI1XsHF0NJEVyCFnH84mY5s9UV//+zyzrNW
4TMP3sGpPOlDkBgWUEWU1row/z0O6YETjpICsaMJYT79lBfx7g89L7q0Yw0WxlPNOIVGD/ku0/kP
lGdTdMF5+A2iI7b13+XiMQOsrvnlYoaT6myF6RbpzFzE3oeQbdtEE4TGetJcVeGXbvJOk7F4X2o9
cOHI9cwdL3C6rMUcCupAZa3dgFlM1eVssuytPyAzvPhxgd8aPU9tXDnHVG+FJdS7puwoG9ZErEsk
AHNp0LPZxsSYCKSrV8S0wht/3KNf76B/IxCbMPKSZUFp2ToptrfCag0f85FcpEOpWSyozhw3UN3p
/9Gc+I6u9QOt4STdEQ9id9lK0XASq2bFiwIxlBUAUcoTnUTq7zAxIdM+01eVvCrQZ6/0Jwx9jTze
Vdj0cUo5KxKosUQj9m4wjgzFaywtKdB1pk35l58j6oirQRDBWsi1wZQ5wxTqIO2UjcSYermTi1wi
kDIILse9LRCAE6zf17oDvkz9dOt6a1oq9RCWlZx5GGRZIBNfj5FyUAFUMZ3yNbsGd0oiOr9Ry2sa
aCYC5Ij0gf8vqpgEw+wLnYzvoQZejTlePF8sYokwRZtHK1cUxtqT9GDiCSrU/x8GekzvcdB5pTxR
09wiZ4J459KCxKPQFwh+17MY1gdRPKagT/1ttSG+x2S4wroQfsJlz0L47gYEWhy2rql21yHw6bbg
12NkMmB8r7UlI1liErsWNg1Kew80CfmV5rviPTMRkGhvoxUJ28kBMsCXuzgU95KNPUWQL/ifONMA
trk15kaLn2hljZi7r3ARXg2hVShJDU6Jm2+8jY4AQzYduCSnnUxpnmJ36wcnUNbuno+fT3Q2mMYs
Qbph5Oxr+AUxw/Vzh32Yue07oQGCNbv6ZwzPAUP4/FSi8zRHEw5kRhhyB7DO4bdQUtP4Bsi1H+De
gzUbKxFFSB80h1ScATvgv0zL8ClHiZ8IGEtQOreu7VKy2E4rvoP5+yuzD/lvLCwHAsnL0b/w/QAe
ew3sR/0Bhms/UiL4SVIvc8QUV3ZT9/YIKQyvqvrbmZJxxc+hRuPpwfDqhPSro8y/rZQ1cY7HsBYA
Bmt+T1ifhhc1NQp4aTkI+ESgXenU/WzMEfO+Oi00p/0BJTg02Umn1lRpbQ7wJlt3kNhBMe0IzWSF
5mRoIpmOTZSG1J4ytiPys9L+kFMhxCt/MseVQF714CjEvrPFYX1uHWSkob1GwT5zJ6T1me6GYEdN
21oVewZWR3FNLS8iSAyMksAWFl/8ntnp/A0ysTfem7C7Ln3XYdZdAEsVQ0EUpDfWMETyXc+RfrmX
Jiau6DNKEyN8Me9qIjXxS96W3cFQyFBY3Q4Q7ctZP1EGIYZGwj2qpKeM7P9eslQikHlxmEpXh3j9
bUoyi8irNE+G39y82CzI604h6E5I3vzqPA9Mw77DpVkA3cP8fzAexggnBOnje+6QcoRW5uIkhREc
ivOtSzt/awz+B387JZv5rDHDHP4qiThpFNW9083CQKP3Z7Lh6x/Qq1bC03rdxsdO8zce5vpSvMmi
phdSSTJqNtGAWX1r9nmkByn4hFlNHGloUyU/gcsEVTvnWNWWbG2loy7y6EbuZoqKXEz9hdpTrz2S
xYOJFejKEXOi0yqRuh7MelHf3WrZqvBbWmwM6Rfe4OQN8i3ddkNTlW+DrHh9Xauk8iU0GFTPKa2Z
L55u8/ZwGC9b5ePfrWcEk4VGNt0B6rdYCyI/xwTFhsBvuvjXU5eu86W+3vwPA+VmfkHBtiXbBD3S
j4t/Wg3KmkB6gE5rlkWZSYHCmUsXWl3gZ5CL+Xm2OvJghfyJXmllVgHy///JBQoriWIDYNY69wMa
5L/TFoUlvu18wqsEhjpyozox2vphU0vXvlH5ahfc3ReqodcETwKfkKIyBh9erCqWmSecXizvk91P
cDymjhHYNwQPBbRyY5xU40nfszNK4uG8Jd3cmclGNhskII1J2pjddSpVA6ghupLj5bvI4N4cO3Tv
SNdYxZDvNyKl1pxyHJY8ICNev3VoMJxpmd5YiLK2AXxu2Pw968tJZNxuDwA7pfPJd6VtlNKTd2QC
Sf2WcIkaup77AvkgAyjAkmSbPhz+Hf4y9wOaiEWxOJvQXI4dHQIJYd/gTciJsO4H40THO1N/O/BL
i+yGANBae81mtE0fyipL605vPUwsLwK8gs8wWSrAdZIpJKZnc2Mz7ENvshvo+QwnpuK7cGXGXhBo
dWZAOJ+viMUtvuLWFiqNlKxdBUq9LhJIxAOrHDkKg4rp8TrsdwDKOk/V7IsCRxoyvLIYn/6G8xQ+
5xH0kgLjTRLG8+ridslECM91LKxYhIqDbNrQAtDHmvdcDaJQUJUVttj3WM6F/9jUIeJalow3ihcj
00KyhYUWXNHYFspldOJcTBQuGT+iUoa/hTxr5fiWTQhtcXuj2BrlCO2RUyqjpoj2v/QRcfgUtRmE
SRn9pmvGjTg1Wn3plKCPmJ2e977pcl9bAW2ReLVWk0jwfQuMBqO+uBa1R8hqRiiwi3SgqvbIy2Rx
y6HBZZbYl8pCzc3l0jWy9M8LAqFFEpr7GjQGWmQCMrik6ApUxZ05cNvvpsExt64LvB9z8APBUYV0
5OutX5893OcRzzhpTHDWf3OasFSdmsSjkPu0GxiAKYDhAgyYG4UvA1aQF4Ie5e+uVsAJNhpTAMFw
OJND+mScgIZqDkh3jbZ+SFXoTlo/fWDMo7otKlfKSBejfhzkPcyWdvr5IADDjrVnRzvrEQBWWoM/
+DR1EyAODhn0QTM6PJA2lBkPdl+/Q0BtEp1RuI62VAqXJDya/tBwU+aaLqI8NAsutrbA8Rz2cnUU
Tw6Wl4DcIdy+ljZth0QWntq1Sd7PFuJGVBGl9Wo1GtuMuEckz3SW1+KIBC/G+RCdNcXEjdvsuN/l
5dDQRFgcLSqtdjo7hlx2yTDha+azjQ58Lp4KzenjQGYvmDjM4iKtOuAFHHthOap9tTS4bwzoJEiQ
cN3b6/nd2bdffPgNIMoY+9BoTb7w30Pdv0lzft0D4scTJR/aXwYOz7tAj4+0t3cvKiRFemIIepZ6
SayUoZpDgyvfK+B30Oh1551EsS11eWSlfU26LBpRuayKQ+IUzCyLqCCtTCed68l6gaWRcps8uGyJ
8Dz7qmQ2fToWi2OMKkT0CJhaYu6mQmShpsz+2TBy3BdxRlMsmTjO6FkKdU8GxCgvuJCcd+nUXtX+
q2R/dHz4B57Na9+gsKgRx7JyYPUeJiwaip20y1l15k2pVE1HVeUyrlKVAn1FRsEGbg1Br7XN7VB0
2V9Q4/yzpy8RXE6Y6qtcfS2Qt+T1cqUgYJ1QJ9hJ0dciDU3PWSO0lXjWjSDkSyosAIvxgGgSnpYF
aqBUouilccpbR2JEIzKeIAw53FeFEQ+T1pryRgExh9c8d1ub+6BXaZJthE6jv4Es1hTfJtLIrali
LfBSHv4ATTqdZIEnnqnW3yyFviw7UQ7GJ0AueIMzGik6UL3OvzcOVC86TuxW/K9TaQo5bp9/o1t5
ZmWL6YzdkhzohtAShWwkRj2ksxHxnUo4/RipzdAtfiHkzn7EvlDl7kOePEoFU4hhOr+h0l996I7G
lAv5/EzXY5xwErkqdTGdDwoEvJYWfQq3J6Ah0X32LCe8HFhZzrqMFLc66UaiMaUjeaZrg6a8hy8R
QsgjcxbP1+e2Oypjq7Ju7XodNRAZZ4leiE3z/ilQwBJxOwOiUfgWORyYIP81RVzL4Sy1wNmR6J8J
FVWOvlnbY4YTN2LgVPqH1QiBztzizYPuCFCLIPTIuWPn7RnQdIekBBb0+zTKBQ8I5Tqae6l/0WWt
h93DLFkqJac5yK+s0koqMkcyr8sxl7wVX8CaAfl2CQgNqJ3+MrzfKMSsO55WckvWFqffQQBPqFQ2
5J5arjtTm+mCNWsi1V04DgrzobWwPWE5S/EOvFHXu66HyClq/K5IMxWWu7/Woi7FeyW2n0AB9trE
UlFMgjj/DoSVZG1M+m+OS3p+dy/adG6B2H++4uDxw2EeUKuKDSe/KfiIXAjY2re2yPc62+eTA4oa
PkNWJ55Ic6LTg9hj2zi1HsxoA7LbwG8U2HCRAlZhxC+BJN3wyuyJt552aSG/ObmjCzfQ/hsJR6Y7
FuHm2GMc22rmNKwbcOoySy6OI4cfFpEMcq9EYBhoIctCG75eO4rXuuHuK4nkYY+H4/jyPqNWvJ2J
O7TyYjzfrqIWFTDftQd6NkcgKX42IwxByMm8BO+As1jRjd7c3+SFqU0Bb2r+ElB6zO4dOaRQiPh/
tHPyuvX0s86QleZFyxUDOL4Cz/lAtzx8N81a3seEH3WT03iZti3NrzQWcEBR5JcthMBtW24YxNZi
EA9tKXnsnTKkFYspoMmRPN6nV0sinR200XqlVEsR2Pe6A15SAddj+F2Le4FH8SpDsNEQu/SSBtP2
qRaRpobAFKc7B8ZNCFn7rdW67gZjqGLPF66k1kjAC+EqjPnk9KCuQPXnP2Wokw/6rBjDS+qbjgmo
1HuvPyRkJJNHMe5TkeNc4UFj3TJC4lpnsVjWnhNe5r8odu/kv6tB18wP18uMRnc4j8XkxJbkrXbO
t1Kewt/565Jw+nS4XX8MTmukpNrkm1Hn+DkmidKuhWyqAB+1h3opj/LSeCDLlR2MvZ2hjbRVyap0
kN9mQJMm2rUizutofe15egPRR8nwUZBsrNOoyeEatw6rVSw4r0L/5SDVomUB1EWW0XPxZk1q7idt
jvNjNnT506WZFbaZocK30G9pdM9rI5Pnlz+l77Ygw90WAFCz/EBXN4FMSBUuMEKvAzL5CMhKWSbm
6IgMMuOA3oGFk99SJXjiIIRw4WLmXjy7rybAV8fhNQilfOOfDPHSOqxypbJddjbBmkv236at9xbE
TJah2vfGKKo3DKETCD+A3ehOXZcxYYb927n1XrBeIVr+FSAAvxJm4IiQWCRT7Km5YUYBv+K981Zn
Hr1PBQIMI8i37Ap/WEFR9LIPgcXq6RajivgwOmhtCSg9JqLlSypkQd8ZgBRWxqlEbvog2NfH8+DC
qAhZUE6cwICBZv+EwIQgRE2nVzkwmO4tSIY1hK4dpM5amOJFnhenHiFrB2ZNM+0jCkfnIOZkEGM2
Cc31xwxoF94CCTYfeJzBP+Yk/NyL5PsfoKRFvv53AHeOBQooNltmHh9YlVlt7axZshsvG0mvp6q1
1Qfu8DmnzKkuBNQgxVNGzGMigJXaZ8pdUH7mOgmtRHcsO82xD++SZi/j/Sv64eQYDeeX1WVIEdxE
budVNSpcku3SL2NSTHmXN8zPy4d5jhKq7Y60s5KdP4yyAw55JokM1qhTZnUFw1rdsGXW14BberyW
JqVNH1dX1Gx/nW70IUZQMeR7x9Qf39tizEBbDDv8e9qRN5vGCtWcyTUhtdBkOwvo/amuq4C+/W0L
HwJsDyPfv0BfjBxUf7lE0cO4qIbAYMucZUFZSzPL6I3J4WuOGsy9Zu1z89wej6mJTL3/4ix6Tppb
Joo5BEpMS3+KuRHK5mSGWJC8HLLbe5+sAF1hf38lFWaXTdMu4nX/YIWp7xjix2InSxLfwUF9OC6k
f6MG4BVfFlSah/FE4o467ngs+6LIcbAm9IgcbzoDPf2mwVs7blJfO4gQJoWKlZfkYFRnV0Obn4CQ
UOhMgtR2F5ngKWQecKCIaidGFLpfa8qdWXjOGq3UmRj672okKJlLEigk8twNYjJil0Ua1QHmPsK7
99xaG+dV3GKI03BpxQmrvQSWX4jzc87UMZoEntVUFeHQAztwJcZCK0zhig0JR4kNq1EnXwxSnDnd
hzZf2WCWzhPvA3KCbTDDeIfAJjBUMuWN5WieAmKZOd/Qmgia1gNJ4L3sq0W1OAf3Yyk1bhblRxTz
OCzh6CH0W9KRBxVDo3Ch0DXJajJg3WxqFBWCDvdOkM6rvQcrHR58u6EXXA9HPXUqc7sMlmFjS3JW
IF6MiuTcvbkWjMZ0hnCJ91mYziCzwT91qrW+MZJy5ZN3zwXzcbJlXNwm3bKkMNpaUHkA1LB/TgAr
GYWES51Q06qXqB26Gy2XBbN7DHfzGjLP6Y6bC0Xc2SdwYckVr83KKbSuzXaiDB7GFf41ttro2VBI
i26RAdAdZeu+d+8PjbC9bB13F1RhNxfL3RUlROxlKvs0jt+GloUrVvFtlrcqQEcerm0wrkdIa80v
QdBWlklw0ugdFEewJZ1xkuZmZFyIs5uqLzkP20i8afwX86wec0O611RSBBy2NJXFn28aNqaXABmn
xfbguLNzt4bRIPxdjXOPw1lf5Jkwi3a8KLCnkQKFEeXO0iFNiRCdtjFYVHRu/gLgbrxph2n76Sqk
FeFxEcdKq4jbpQa3+o2LRPpMoS+RVaNyDl/8CygEjXn3WXPEzPBnD2SgO3t+Yhsgzusq97i//pIz
XKf+UyS6NnHpmCN82b3uQkAmHTxL91yoylu0q0rd1X6UjVqiWNubgJx1eBjprMjfn88vJtNLgp0d
33tbobO0+GHmbxlGOanW0mokFsqMZ2L+YHsf7437vhLOLyYIJLY0g9DoYnEGE6foq0t4n2uZGYOA
xPmhP5TTuZZKjBWNd2Atg9cliMVKtW6kSJOrn9vOS0+joYKs1MRNlKyeR3WGWOFb83n7234Rc2gS
JBwARP50qT8ctmFU6bHtdfXpJrPi9aU01UBkztchG9qTkyJ0qfroCEREICxIdQpWmbpFOF66Dniw
07q8yCnNeKgqBGpKXwCEr4o8cmWLxrirZdk7gYEeiHMdUTXRjQhvLCpQWeWARJGKvRvx/EJWZ9GS
E8MzzMBiYUAWBWV+rSxJKA1l/JEANZjXhD13R0v3gBuXYdRjZ+4nu1c/BQXrSejutcVnNOJawWTB
pv3Oil8vi7GOlTqjUOJwmT5UhkzsInILxvvmKJCSlNj7fOYn565NIbhp4lpQbeZsZNPEzELqUnvi
CHKruHD9wMc8p4200Hu+CByBwq/bPuDbJfZpjqMMk1cqpL6KCDR/rDBdwh+IV/9R+2ng0h8jRoUY
X00OJJ/ZCBzmQjKp4wIYPveWaVu7Qi3d7BCNwzIpOIXBX16SMrmYJaJr8qGFyI6xh7Z16ixpVLRD
MAdJl5L6Tw9AT95b0pwIUeXcsvljHRHs4E6WZS0lJZ96fmWoGTJkP6o4BT+ZZoHuBbxIOm7v07Ir
pnAh79Qz2xoo0w7qtGcVQcokdYlL6Ova9t1eKgoGt/U2OrZ5Sk6zESP7VNZTnT5n1BgJDPBbZ/rX
/ip3ZN7zULxW/fAwFXl4Im/SUBEakben0iKw+f+Q+WNvcdZ3DjNzHM9/13oThyCiDUftQNkZm0YQ
RMECkapxeK92TvmDfdQoVvZaZJPvdIc7cGnzj46TbMpl1DzuYZYk7Z0nzQHlS3An0zN/maqeFoRo
mN/ftktX0hcvs2DMdXu2oZkmoqavH3IeheED+K2RwBk9gjzq4JnXYnDf98QXmxITTqqidbxfFgnW
WCMmUXnrTCP2mmrEk+fnFTI0YmXosc4OL/0O0sddptdq4EzdM2cZhheBRQ+w5ofkJNxcSA94X0pu
MhsPJFvNVtOOSGMnu1aDXMOVqYtudA2ImAL2++4rjel7wPuajOUT1OhaNgr3q4pc3kRIZs+RVSMZ
rQNqXwo8w2ucpSLTfJbrzGaxJEq/fEvNTdD+06cRO878EvnGc1Wg0digzRBGzVHWo5iZv6P6RAOJ
IYJcit+N3jztc5ATXsKAMscwzgf9qwe17syLK35wrEu4ypOJ/qrnwiHxBMUKxVtk2xrAuJg9+Dyt
B6aXiodaSKzTnoQnZZRkXmbY0O9klOz2iqRafJLgVtR2F1ISxBCa6BksmhUnKT/kZteu+Nqxw0aQ
hFnyulDOKn/3ZG7+V2TS4R7HVd/+db7HZXKSx/ZrWkDVv5ndY/GyVruu3o+MaiQFKLlZSMbwWO9W
v9lnHcZRde3UxFzHVfOp+aPP+revKP0JaVXGdN3WQwY8jdQeyXvO9+sLzLSjmW71MzDJOFsRgjvd
q6+HUsRLjeTu+7ASZIhlcs7mpo2xFhWi/NJLnL3OL9ykbLCMtgIpOGWlZt37OF5Az3k/+IQRC8MP
kYPo07rZ5sOxyp/uI310tvUpWzTwgyKydmQtrMP0bV6WTpuQoajAcABHnKP+LuU8VMSAQbSVYJby
YxiTC09+3JDcNniVVkLO5LZf5mD+syOZ5GY+iagfJiATeW5lreEzGY2i0/fLjVQkdZnciu9eE8bT
C703fjoRFkm8cWFOqH1I7FhREYWy78IOcN/ugttktVjhO6sLIgr1bQE+gHejEnqfhy+P1CcDGUi6
1ECug2YmShTadsr62KF/69RNLoymBBnxJkoAHzQRTc18DKR/H8nKvm/IK4b+TK79tuwYsnQnOqPa
No78E7Yzm1gvRL8lGJQHcnHuc1fcGpDxysXdPQpv5WJWESPgcTjJ5+X0pb4DLYW8QIEaS4t1+Ylu
cNPVaAYHfndO0bY2Je6H0JRnH4k5UC1wuGCFNn934SpZqL0GAwb/MdhBh6KlFZqYsffYFIKcOEpp
IYOpIo70JS0W+ND+plVvnwgbGmBOPHCC4LgoZbrAUUUXHOlNAhNmWwxCx4R8i/8M3T6ISwRLpZQN
PY4OCB7pMqhqFMnNrxUhqAlGlpBoGV/sKvWmzmMYnwno/GLBOfAntU1iOPuEPPmxi+eMYfyZWmac
65CO95q0HKrvEoji3M4LMDBD6PjXth9N4UIRWylkOJOxNwafgCiBXcNmN+l4WfvxQKtMEOEN4hZc
u8MkU3J6TzDdKuuJ+zj5ja8QgXmqI34FaroMAT7E0LZwoQf8hnt0jHu2x80ykSFt3y/AzR0tWMXX
mbZJW/cpdbAhnsR155g66AZqlzXE5baQvsC42kX/R4Nlsj2xJ93u+Rq3rE0OVKyaqw4F06DbDe5h
n+eJRgS4IgwhF/+qZaCsUDOszDHkCduv6Rlb4Gtmowcz/Hdp1ekbHMo7/uX29I1D6eJ/O1XF292S
qtsD9Ety9uBXDXxt3w3kwSSNBTrcfVajuk9Iw7ZghsOb5/yZqsOdDUIuyhW6MpOqlQ6JUKCZaCpo
ZeRjl3IIc/zAdGHM4Z9lrfnL6QJ1ofhQIsOf4p0J14giGNDYLjaANADNOCnbgcWw15mKJBjNyZsh
3thalQSOSi22VW4GMAEGEuSZM7+OS7BLKWlheO45ig/6oiGcuUAM9m+S+WTh6Nn497jqSpEjLTlG
L3E61iwJpPi/bT7m8v6BCmZN/0hzLWfHLKBbZ6iYxd7ylG56HM0T2dnbKPi2Y+UqI4LKEORxJF3c
rHZt/DQ4nHfhmKDbVM9pvRXro26yXCkrOq1uG3qApCQU8aNHr+ZGBHbQ+u6swdJ7Gx6byZI2L7dS
T7Gtn+mqWZifb2o/jAOheYBh5PcLqxpOGOUX1gZ/bRBuDkU5TwlQRjzL0tDM4GStGhHKu3ENwAvl
KMMHlrlOWFifWZ94F2Snh2Dwzgw/yPZk/ViKp8mXoydxgMIkC33aSh97RMjn/ILVLwcMcd6kPvrX
+MACzbeUjaOD1csEqUMnKLppIjhUqwi4yHL69BIjyzTwYklrr9Ye3yVR+SI32EWZ7qH4DE8WGJ1W
1nXgiq3uF0zUAeRisCUuLKwDSbFZJM6Q2ElQv8BHsT6+M+ksm9dcwU5Q8bKVAVaL4UrNj97Y0/ja
1ZyX5z2Tx64yVgNOKrinUqI6yJjYfvzpWAALQGDC+kzNbq/M0cXkcTRJyREINSDnMMGZahlR1oTh
Vp0BkyETbrWhqaeNNAZ/e1DoKWg7EHq5Cv0V2I8VbE/UT5QI2lemzk3dkG3NKYHEkHoavJacunUL
ZXtyrhHs4DZyWzPlZPqLop/Qo9bfolzCGkGC3j6ehadWDT66rUj8YwFqMgCZhItIUCd4I6W4gkY+
/d+9EkxlR3YG79303mqE1M18twKDVCtDqY9qnlxmDHaW3LB4fzMFeM1Yl8ExkMLY/yWluGmqnlJN
+vdSkv3q19vfa1Ql2UjMnFXg6XD5+aWHBUnFUTH/R/QGHczvFKxVGhlLnLfZ9w5ipdLp6hbCvJxE
7XfcSgcYjrIKyHPb3Za8OSoUbWg6n3iPmPwoEuwtawbE/dAvEk8WA5SKuGzk87LTez28Ecq/oQep
ADd5WxHxELNdoD3Gpdusffpmb5/cULr/2fnkpnSi7FSr+QGqDLEg4/GzI8DW0VuR4S2VBqMpG+lT
yk68Juxhj6VtOmKqhVqkJm4T35jXy2Zyl3ukiDQybpG8QJkHz0IWJkMs7BPiet46sLyI5xWOUamY
bNbVthvz3Ea0dENx17GEFyS0HVs3kOX+mNdxmycoBemUsnZ9bxLmqldYNt9gSaGydk8oB+2f38/1
dHQMZugy/mWu2LKQ3lA51fSO6BdfL1kQ2EnyNaQZlWravgV0SaBGzRizZxXXYCPvg601qazLTxgT
okGeO2j/2F9UP+dHoVOh25ytNqv+bgmKtfYykgSuwtpCjRWUJ5ZaSfI0J1rJVuRC/1aBX+btQuwd
sn1kr8DDxGoCzs+cGQ/bII43GTzPA6mLI+0/oJJ5fmHGk6/ULmk2X45osLjFD80Skt5Y5w4Jqtxg
Tu3yNFbUtdvobmdYL/C+nQVlLDYKdGPGOxF1eWB1ALe9HqAJowXl0SQ9ecs1KqxAdaa9VFLWhWUh
J6ftw5TuWgvhFpHYU4Vrt2+fP5ZedEOvHa7NtNCV/Vh3hDY4WxqYuJiy4oFebnKa32AXxkWq24Le
vbmyFwvnlNbg7ThKAJDAP+C93KQNsCRMfwopa+IvXMrAS3QODKx15SAZZfWkTTZAzeBlKlmhk0cJ
W2Qi3uE3MV/a2iIqh46mz8LbJheaGDfnRb47L+BuT4GNN3pIAzNvZhDqo36cyvr4RVoZsLthXpYn
+mVpDcl1mjcpy7TvbI8jQ6SVbk1difs3B5KlzWzMCwVk6ujsDx4qV7pwTAnMhOlCSjbYvoXmc0HZ
eWbc5qkLlU102uygCMCIXhyVd9ZtA72R4pb5SOJh8Oavy3aHasE24NuaZkCtvkMuEvvj1+UtCN5f
rZMk1JSa8ew3hsOvm0repbF5nMDUyApqlYIoKsn15PLXYL1uxCbDIegR9q1w2AqjuWoy+xudJ2BW
UNUj9rwrJnXouUe5jkZZRvofzn2lQ13vtZK/niwbjg2Ye8WpoA9X0MOPSkKIH2lEtQxh1+ml9+wR
GUp9wI6KqImF8a8zAPwx2TJXYnS4xUfrh5+scCZqMCItXafjqN3t9dZwDaRbFxSvJUQdEQm7wwnS
aOb+qo8b0VDvtIvf7QrWzQ2DhTysdUpGjicT44ecoiTKkAewEHBlDWu29wQ8kZ9W94YIm7rxa4Aw
/ada+u1gnzBfhrscI6S8arTr9+QT6i+9Im8IGBqJN6iX5GPnygaKNtgI/L1ibzTrh1xqy2slzo9O
dAGmzX8PvDO+cgzz6U1aqFbA37yKk2LGfEMUdlXDdwYg2VqjQYQAi9Zm60b0njUd1jJ3qnc9Jluk
Dpjx8oThQ4+FTqMsUkBHuFLSSql18bW+Btz/sJL6xz+9X/ktweIpDoh0qiUOoOiDO8086THiXeet
tpqMvwFxZGHn6GMLkTGST+5pTERqJrJMTwxAL7cwY2Mj4X7VR+pMPytt7DKvR90S3Z/BsUH44UGH
uXafrCdrEJ98s7iXL8t8pWZ6TH7BrAiBS6/EG6i8jVgvuCmaC0Qt9qXBRDs7MJ9aOHrM0tuvufBY
UDQW1VVOvWe9XqZUy62u1EVcrItSZjSsIhwSd5QtU3NSJDLVYbqQIoxldIBkWc0bzP17Np6N95kU
yJewHP3p/EyL1mNUT2mdvrk7/KdwCO1lsJHq2Q2ZaEPJuxrjO1Bu+HuPMINsvqte5PTB6jZvIRSu
AGfD67Pqc7ueOMnKYSpdvqoAbJJ+FMu/uoPa/+q2j8Ie2PXPFu24U4eulEHc3maJ3B+dS3A5kqN+
5+cLA2k8l2ZIfLcNjgK9+pDJgbAuKHWJyVW0DvcuRD0zzPNw36vVUcqAsrPDLTVu8tb5CyJ4vGR9
979/G15PbeXJt7D3ORN6537upbPy4Wtkmb1YLIilf4MadmQwcEljx3Yt05FnIdQd0YezntPQlPeL
cRdqBb3YKeKQkQKZBNJwVYhasRx8miilv1Xi9vwlPZMa0MMEngWy6v5shR0R4gTmawVFofF7NNO4
WIwxo0AfUP9otIBfunLsD6J/MtVbR0ylFWD2fuJulTU9e73A5n2qm13niDQYeg93rpuN9PKaYvCv
cwTh/V57c4h/s8GgwW/trBRnojMNMByZT8Zva/CKRaOprhCXAz37ZqklLwmY4fM/Lp9RAi3KGzWh
c/92ragS6F8/S4VJisnFg9uQAF7WbGCF9mmjKWzf/Ed7J3/GHo7lqdsQhBrUBl7PAHG96xGeCxCR
WbvuM3e1W5Y+vZhJEV35mJ6RdHDlINR8xs0irLdRLm7PeUXG4ga96fbJyfi+sQK5ytHvQZGli2Jq
xn1msPz3DY5wIUvHRK3uKkz1/hEiupUWlsE30t80KicsyC/1qWRMGGuMLxeRujqV1h9QU4NNTTqC
HPMkBOgF9UUr+ndKeEbyOY7HQBEug5HWozw8yxyiQ8z3F5REelFur2N1Uv7iCSNVG3qTgkEP07mB
xLTr1tzfzGfEE22V+epp27cV7VX9iRdp8srlKfW4Z2XsTX9GcE3RAClVhCSpUfLRTgfZjk1lWNQ6
cdYzoc/vFnw016a924avdxYGv7m9ThKOmCsJbXh1riiQA9kt2aVL2H7KQaoWmZHAhwtAT0TYQpwZ
tKVMrKvs+uaXgYO6JDKlJHY8KyRH015YAo1CEuEpf2iGedkZex7mce4lIFJoPJx7fyZBHfDs2L9l
3G6fvB9rPrFcHIG63AI31WBobLf1CEM+4wTkMTWl3FZeMPSCL67uYr/guocpFxheyBwieDyk3nub
ncFizhcfvIUooubinRy1GMjr+DEwk/67NPr6gkBGhY30C66vdWDgESpmVknHjddltDhOxgIxvMir
I8T7abJxOCEJqAQ30ENiFVHNwwdeBq1T30IjefDXhFf4g7rMmJ8FXX24h8BIDAnKxwu6mrYAGrPd
GKPzcxLLICoeBbjHGdYovdAMcmakyM2VcIzgh4IwvfEzGGrL6jH1i7KLJktQsWt0ohxgRYYWtcQd
z4JqeKNmZNcCOPUiPEYFXrIpxzTiG+Zz884DsXj+M/6c93AGV5mMmNhp/h2skjXmqY0pswQKgTva
LMACBX4uMgICSpByrjS1NnT9WwqCTWhqrFRLeLx3ixmHHG+VpZogEJRbWb9G5cew3+m+pElhG/V/
tzZY/oy7Z8IGO0GrX+bs2T41d6gUaClOJhsxuM0m58ehx9CGCVfAuL2N6ngWv8Sc3GJY8yrWEWZc
WV8/RI4/ncWPjksLk7TlgYEbliQUwwU5vQPtklXixDwN2LbO4UzNsjXJPIERBqWEYrQvGGhB5BGK
Ijdr5Gtv18Ny4kptlwtK6Z+2cnh6Ip0oVYgJuZ+JIznbWeGjd6xKOybDoXHoN5zGku9mSTzhFMHL
6tpmkEl1vUFor/Hvt9SG2Y150Lt3fPUgUDj9t/MPYu8EqBFk7ectk677ha0sD3cXkAhqvb32sYVz
8+zLiAs+a4lSz3HPQ8bXvpCeya7FktgpyKCn8d4bEWwzwT0DCs1CgW+izkuy1+jER1UaHkAwHdDK
I6BK3hBstVWbFfGCUpqKKBGUwDRdAd3joFkOM5H0+Jx9lKEv7juSUSRSM0pgvJuoSFfcCDpFIKdh
VF5jKC88yyaEc/N+wr6ljcGHAlCDbqthFUYnM5p5SSWfPolk08SM9vMMn3yHnXUmCjfnjgqHqknY
kKT/Zv5HaGHwDzXT7M+rBPC2J+VNfBPZXyWMo4RQKTmnIAvtERyxRlioyuFXHOLyWX0XK+T9tGln
XKj44cksbivGe8VdMgEeXLTgAMp542CbNeqC33zZ0BNfgZEoN8NnlRmTvIBd1ZHPeV04vkx91yEJ
lw/jNvgdRIwXRzxhJtHSlShvTaw9l1Ss2+/B/XK6M2NzFm/qimvmGbfYNagAZ0uedZ2n6aB9mavK
FggSnthnIXRqxSgUuLfjAbneN77/NbEXcLkDfR06yrVNRaLqRFfFTQLMB5QPo93070KJz/ZtEhQs
mPq4/jBFIKEROCuNuVCk5hun1vfIN70tpIvueqtr6q5teQfff8pEqveaNnRhHh+NciMcKzJqvGMk
Y8308u158Wo98yMExV5Yu+KELEXdiETgqxRhLxE0Qd6xBJ2+Jx4mqP8SSmSfTHIsiKs6r9QNVZzq
4fOrKcZc2UgajDqSAq0zIL8AlCtg7ENeaMjjIdfVYi1L6M5ks7b74pQf2ud7oZcdJVIKgqQQCvpM
lV7hEPiLNVd8ah6oboyqIoX0ZkAuyVYRSb5dTb8HA0fiLfX4W3aT2zJPoxzs1TC+KwXtnYjceLIP
Z7FDyGw5uvzsbC64cVnWsigRRDbtiyCpCobgLlZvgm6DXB6uCvJxt6YGMf31q9hlWoZziOkKHPS8
ZarMBpthRQb1soiE6/YrRlxA2EwN/81DM+I/DTjnjh9JLNeF91NqYUAt19wDZIcpQD8CouEITkvV
0edGjcShFx+55COvYfAQi68LQgoQNUd/ui6P5hbCW03SJbd9nusGJMkEv72D86M3ql2avq2PfvwV
qFEm9hWauLqyUwoxQsJm2QtrlZQH9bfiSE0EaLe9B7H27Kpbg3x9sLUKKWvu5Cvrp4WFoenguHgl
T2fXOOEmT0nY+EeksSiAkcta1YX1KnsXA2uiVQTBqwdu06fHf5nd5Y0ZiTtcP6G3f4Ff87asgVL+
/Op1lJHBCAj5nMZ8w08V6vgbM6oqaIjzIkw7RUNtEooIjMEZgQwwgYtC6jtIzIl5UW0iPpLP/cn5
L+XBemLT7CMK6lQrL8hIdE3xQiKwV2vyKUKsPoIHJB4SRZGoOX+HGtKMz1IJ/4cdOBcgzIZNrBPM
RJ1cfIbvSdPN9jvAeP6yrn0JRxvTENfLFf7SObZIZgbN51MZBl04qFQPxokG+hDKoaBbS/USot2g
6BLbUzTDZXoo5iEKCL3il0EnckBgTFsG0PZakvHqpo3lCTXVTbc/r17zfGK3ZoITea9vM2thie0w
Wf4MYBNI1KZWfoA+R/aOxHV6cGEYknwSgF18bJAZCOiOa1dlKehe4sr7r1h4xcGsBfSwNirnuZ1l
WdzZcYkQVgofhziXyJbMTf3BPmS5g+5AYoRVa7fvNotd6W/ioWUEoM2gu/vejEBycequUcoG6Vn8
pbpvqPdjAZOQ3c/8VLPdTjVllOsDVapElqKnhb+fAh5o9q/JjxSILP6waraK6kgJvBBQCqgqClPS
FyamhcgO/ly96DDgG4Seesu/GdGnQ0n0s2ciZ0J+YDTyWZpahB4dqnvk3wTbeOm7oJcB9A6lPbm2
uITUU/EvLfhPkWznnlAA2pkwdtYYpLns5UXmmeSMraUU9GUCuIbXE8paFGFKrTCYGSnM7bciJc2o
8MI0KI/gLrZQp1jl+ZC+rpTsA5Q7fmabJ8NabVpoihwpxm9v6bFegrUjWnGvDwNW2RWlIhMyym5A
oDlVTNaoaECv1MVKVXl5i0r6KWT6Zg4Ud2ALyC67T3Q9lY+talrCVUPhQt6q9sSsh1XuDVDC5NvW
ThEA5/WMjuLH4Y1gRib84NMxngvQ3BOd8U3JSK27GpRbSSa/EfCzZHENzb4PQFhTfeQ7OpvJ8ii0
CFPrfe4X0/uvhOjIjvSp03NlSlxsEF1y85OQArOXHSpz7SIa1i5qFifKflpqhCxsp5QwMOq+fhjc
83ZTpjLP8DJF4lD/SGNpllt3Dho+kIF8i/WuoUzcnh730E2wYPpJO1UgmYdQ6lngs3X0OeZ4Q10W
UskgTAeZB2DK7tL4WUnvCDBUChafb8IjkmWDEXIz7IC/gGE7e0XBAxGtrfY40/uG3MYI9c6ze9gp
fdNKq4eRPWG2XiUtYj96espzlmo+KrZG348EpfXyS1e+842Mz4DnZTNJGQ6avrZ5DJ3oOjDcCu5A
Lw0ehwbYVkp3mvlcSAyyRHkSvg1v9Oh9e3UVMd4fgIu9J8y4416IRoGCa82wOeAOnOrm53Yem57y
5JIvD2qkXu+YSSrlagKPw3dzirkHfHEvHBL25qtCrUxha76gqN5GR5P3InBnWRaQQgbrHBFhXrGu
1zyKjvTTB2JX5hQJZU/sPWMkBDThs1RZ3RX1KOIaCTzJ2ey4kxhv+M6rCk19MItXErzVGwd6jPu8
SQJhUUTmvL4gccJf6z0o95R5me3yO28qkUWlWJVOXhzN8f7nWzrlPXSoYcu/D7kIzJMUoL/h9YkJ
GIcowVwXUu6xywh2vN92uwNac6ZtscrDZeMVboI/ZcVKNCYNLt88MiLpPaKptXFoopX5Qpd618SQ
dIxJUc1zkgy7HaJ+xkJshHf625UsBcvXasFUPRtPViAbL+vk78T9k1ikPnmjMpRfKt6Fst9zwOw1
8rD1MDlBPEnRWLlVCfsX8WZX+R+s2BdMAHetF5oJ1JIjd2s4fTlGjrUVcMMUh4u5+XukXXIwxVON
bixdtlD55lP8FDAr9egYLZDcjtibV8pavxyXTEHYRnoeJdZ4aUpqVvgi38UtjEw5gje6IGKM2k6U
SjLSJbYBAXHOL6e1jVwM8gz3hduFGYkpup4O/SAxZVmXaEkbVL9w4TCvBq9/3JBQI5Q/jruAYH7o
6vrXmd9kpHE7HRXKduNVXgK6EfKwj+GgkoBrOK78tQ3U0QbiIm0kPMDltjcVqtYlo+X8Pabd45gQ
WPZf51j95gJ0zkXhMDwWIvkpWSFQAQHMr9jY6sG25hq/DOb/1eV/6EXXZa0JEtVHdth9kTQ/KQdO
58d4MXHrSgXX05vxor0ZT6DVMYfnWZyLwPz2vgXgYvSwPFCafZi0mIwqmdlmkQgZGAiEJi+H0ajj
o60F1nUmRvU0GS/188kwTx0aJ+lX5GOX25tAGBXz9iaDxXWRFXWOCnlh7USVfI4+9pQwi7ycOE3U
nMe9ovPz8EOIb4EoPY0ofFoJ7KK9hhcgsiGw88GWzaFFJvtQq7v/k7E93Da623FFC9f/cXG7DyS+
UmZZYRQXIC8vlSZYdEEGsphKKjoDlVt4mxam5cFO3BbI8QX8IsAiaYbPKR8gbOONOPiv2qG94v+c
naj0z1GeyP6fT8BPF4hSX6jnLngc7YVYQjoaTaSVmA90O5DJa16bUx+SysFdeVrfpmgruxuSdsPD
bFZyKYkMFRNLdGZGApX3L2xl/3OHcC24Wo30CwwCR+dxgJxfzzDWG8NHMVdjrfH92zL6Nf2502yI
k7Q83MD/vMNiq51w5Z4RD3D2ZsayW43P623lwp/wyhbIGAl/gUgVaPaXssUyOnrPPmoirKUq5KBW
Brg1lcgzN7mECJN8FMTQnASGLNjDFMyXyWDYESf+ZJo1FzJBvGgFz4zF447viuEOTSGFBt+hP1nk
osbWTGU+bnN9UdvBvPRcpakoMeFX2crquiyXzyUNhrKPj2EPgTPy9O8m4RP7DHccu3yU8cntymb/
fHmvXVu5Pq+lmlLaSyFwIYus3hqUALpPLD7EvEKPdyj2K/1KwATaVImTH23fdu3HJlC7MxNZRGHs
sWiYFp4dgsUqI3k7kJ8rbgngqR2ksiDEmaP+lFbTshFItsoM2c6Orrq29LcCOLSYXGy+l74d1Vww
+YYtKOSw2lCxUKJPMr0ktBBWmE1lKcOtgs5cSZs1PASViJvhf5KhE8wOBoC2OEwK9YPU/+qwhKSY
UoDEpzbLsXHcg04lGTAl26pJoHXA7fpOUFnc6p9dRpA1F1/PvwKAFqOauMRLgWZvo8v0Y2Tteo/z
i9sidVtince/R50xmFs5VuVIyI1VOxYx3UaIip/c8BCVFZUlIVdeha2/LGVVulNtPNybgJNwUNk5
qnjQ2cyc3pgUsbi8BDj6oR3SulGj9cYrcZuA6EfIkFAVdVRVRdhDfv63nvygHAibrXpa5KSUYJ/3
3fHf5ZLgKM/hXrlko+West6BWSXrbkoNPGUVIswxvqS+Ym7WvApsWvdQ4slPZ3waYEULKKOtn35R
qUUgCHDgSfRkgO0kwXfguEyRsv1T3q+y4Dv4qJXW+fUCLTW/J6JVdaRGbIBMu9jfLfnWalqNyGtb
xUPzJ4al6bDgUic/dKpG4RpqEle2fzU7IzyHjvgZV0/Zy13IQcd7MiAOfAiaT+0uzlyKbOsRye3Q
TBZViZsHV8UaT9mPFHv6qmYLY/fjINQL8E3QrvhDuLYP+94VoBqksj2VGRgF2MDM2UDMvbA5YMGN
kdhlIIOHDrnxf6OBHLPLvAL57zlukJkF+pG8155e4xv4vhaaIkmRzeRcXgCSLg9PLN4dxjdTrBm6
yNZaPMzdtS5NkVC4VHPdUq/GR+GkwiPIgAz368N/lQFuqu1vrX4HbxsyP6ZHtwBI2XKw9eRW6d5F
Jx6P+slQXGZzgEdm4aQuzdD1cS1N8az+wCQt/zPm98Z3VBaN11HJ5wnRb00Z59Tqspi/r19333X9
2npk+uiAXxTUVgwvLW+bdfbNKCJRRFyfGor1+V5LEfxZa+43PcOlSl9f10EbC0cZnXXHGw8ExhZh
a0YvmiBz7WuSQFd3lCYH+CQipMd0f2bDVB3YENceVYrMKdBcFXGxyL1HkaB6lPGhSlFd/KqvszMr
bucvVTH5ZzNsQYSmMrXuKK4qqX43Tai04MmtJ+d6FBxUAFwUAvihPOfNri4/ysgbDTb0CZWcr+8M
XKj7Y2hBKRMA1kP9gsMtpj0dWFKRBioNU6Cg+jIRWle4Yp7FF2oj+gNwFKCpY72VD4IMC+fSU9qC
tK1MP/e3usJBnTkwccmF8/kvYPcfmjRHIljDDoSE8yIFh9N7H3i2qUTxFW87Y4DBWgvyUKtVjKZK
19oKpPiPdq4suyakf/bXI1FBcTU/xZH6Du9GQW7rJFEJ05tCOU0xfxxV3Qy6I3C3YMMPdeH1yT2T
H46SmvMLsmMfFkPFEgm7fyVaU1TaQz8r/SoW23XpAC/9wPApw0OPrYddxph9CSs7SNl56cEIi4Fd
xSnQRfW1le6RDidq4kzYcymF32IV/9vcK263BWonV+fesvrvVIq98VHAOQVaRCc3gzY+4xmrCBw6
E8Cv+jxzTCjUa6EJUDVyt3nEswEctWt0xqRfFoW1WRVagix4rz2YhgItJOVagvgUlLlTDF9HhpZg
IR6J8iaH7LZ/NoWdYIAo/NRo1HBFNbCJKGnladgc4srkTbe2WqDnCGR9noutpzKJncZkrIVkfU8E
6+iVC4ZjvnrfPmpZ4s/Frew1bMh7BtoTOwntmK8VT29lx1punuyMcXlbzCCzqsAFI3QpohybAW0V
Gk4YWIRDYLWHb/Rbfen++LXpq2vEQJZvR1qdBUhAzJTGMxKIpPFwEeBTxk1KHvM7K3FUv3iGGezj
SV0LzIyR5lb0fhTGgLKPLRPG3K97gyS6bHedGNktsSMT0NrgVxQIYm5nMcBW985/Kb7zXKtDTiJf
YNrJi4XIqTdvAuJ/pYnWS4cfUsAgjjcjq30WsUeEKzcICWZEO04wRbqfaspCDJfQVVbMuDe6O6F6
fsEA0uehhPQzjFSWmDCztt+0tjTKmpT0FF/rj11PEhxJwrv9vizywmtdr2jZZjiMq7EluE01Ca+S
gxQRVkmDo1T4nN/0h5Nrk9xldl/92D8nOujF5pckn15ooyQqV2RyiFcQi6gA5v9H3CHHfczVBhIR
ECXOISDfYkpusY6qVezSPFN9mH/Ba1leEzRcOioMbKcMKHEjuLxYTpcGMPQ/lVyMgZk04japc3WF
OZKJbM+jXPLV2+OxGVhF7s01631Cp497OnaCjRf3kN33eXPUK79fNtQ90fjQyLueJ3d7z2Q0D+wq
xVE+rsH5HOMUFhRr38I8dS2dpuKOJJkn9pUmz+V2dPPtAo464soe8Od6tUKMOW3rzDisE9VOo2Gn
mKnwSDJWJTYUVNotnPpUaI0y1U3aylmjC6epb6jKsaGwnTivpTxpboVV/S+Z78/O0q9UHb2UNC2E
3DDyjwZt7qNH9WvrLfidLoZ8ugBeyCbBh0BzfdMLBpCfFy8PD3E2ZkQEWwNF6Kt9UEMYzfguRD3v
RbO8B6F1DgWG//AwRh6xb5ULJPPPF0LEN4LNqCul8Ae2OQmz5fi2DXD8+dsYCUQmeEwZLMTI7hob
H+Z88t9G1SkzsbU3o5ud//Oqx8HA/HPZyOfoJ9nb47vvHMZjgTUOpL+TiSNMsAJu2eKT2aImTB2h
ra1F8yeMm27hWw3ds7aWDVEu+ceTHuw8QduY7RXXoWWSF8qBw1CqJWRRBOFN7W/0XZDpRJHTd0Dz
Z89HJsm1w2ugEH+YFjp3HdxQ4RpUoLDmvmM/9L1FJCpFwgt+7aF0moMu6w6OgN76U6zxB2MlzuSm
bAxTSElsmnJes1Xtbkkxz48KZw4tRmJ5fQGQLyg3XXPgAlkR721BG39WO/K5yiKtR0lJxfkMV+FI
/dcGBnKJyjZ0QMxE3dNriNwkZf/pbHlD/iK3eD5Vak5bPodLe2zyvkEUBXAqdm6Cgc1X+hePbWZk
sjhAHmi2AOo9R/2m2jV+AG/UCfHyW9DQLR4JvZVTcgnBK+8vafosP12xri0Awm+pbI9OK6QRoMR3
ri7suO5OMSDHzkmD69iKn+r5tY9Yt373mYgMfv71OsKVPov7rEC3u4FR4ZgVdkcAV5MzBsz8PKmz
ik0/MSUp82oDonKT7f+jTEKyYXwVi1cN0THV1q2grWTgMWWpnVMie37gxc47ASPm73wrEau/Mtw/
hO11Z/FFZ+0tOF0I2iL0j9oKyGjzfhJ0Xl618JXrTp29qzG+eyJWZB9mGgZWYwbfpo3QxnAW64MD
fwxOLOkWT4Q0cuPs4aPBNkre3rbmMvTea6DNgRQUezhg38SlgYIeEjCZBIhfEHM+bx9JK+d6N0ne
6qIaR+q3rBwp7jcEBlu0HZWGxgN9KGhByMBC0xl/B7qT1k6DxhL9TmkGiRzSmRJqT3Ndx3HToJvT
2d63lp9ecbdeDcIyUYgJgC6iw8Riws2EHVFXkTv6NRweP3E0Nn2JXjhZf4nf69/IcqUNMLdeJKsI
+6QxwmngeFExaOZT1ktkBawkcGQbtzSaXPy+ys70HYVOjnf3JBI/mdR4O0OfmC5lGma5biiSj/AD
w3IiSoB9ZqnTZSZKM0Yqdgf/KhJ4Ig2glqjFaoTgS0zQMM73dKvbhZTA8QOQ2yQiDWc7nBw4WGyl
Tw2vZUy9g+Uv6k17au1uC4X7cmYIokUsaYBHtwuXxgztX7a65hPf7DoUyspk2LJoU3+ynZ+LZrRC
g1IyQyLJ2UrptnxTXa5wt9WSIMCJ8hj6Fs3GcsgfWXDT1u+4nRExjluDgZtXml0hC4BV4fmxtglI
3eF9J25GQyhFAOxYvIPBmOFdyKPsX6TUUyhLE0WZhQJ05XhhjxcXHQAkrOkQFx6az667tMYuYmh9
Hcw2rJskSUofxD/Wka1HSwhUT5Ch5IpdIbf/gVB4OSldQs4WX/jDKLVG07u1j3sN2xTuxJWF0H9i
Mk2XsLg01asdq7oQSpZXRVWk9GEUPIZkDLWUApy70xEUaR1MS2N5eSjQsi9Ve5BDlYyyImlPDpqU
a1KovzayrmfBCqZxCkcrgFWbVn2VJdf1ImLBiw31gNKqMYDds97/cJR0SRvNY71ciyca3HcEJm/h
d+qF1jc75W7s0SsRIlVYfSwKCsISjDIxoN3SgJ9ETODyAKbfjVAlAs4Ya0MzMeHwkf5zEOgt2ZkR
DTXMs/H0fInTYl/pDqmXAUH0+qSV2MhN8g4bFEn0bL0lbyThch274cwUGVRCqjEhIpAZZq8MrHyQ
ywnVYmOof5ka2VS/hFlg92+GnOivDFT3Jg5xNh29j498GFfMFAaHeB7U+okq40rMeKRdsTo9qC2C
rlpQqMbbgvMlCmIfc54RNi6Kkh8hUrqT92i4Wfy+PXHERZnoOKbVAHO6BzYY598A4NoT8O6t0Fj7
ps1OXS+tO+/C7CRnrO3p+WkWQvMqGMg89aEvZVnLU0u6azJ1NtkAQsgKsjBw4pjDIJpFUNZmk5FR
IxZM5DFU0JBc0jssgVfE22IpM4ZqOv9XxQV+Mh1RHA3G3NYeAbT+cthWnAGaD7FvZoLpf+/QUKds
mXKTG4aDLt6GdPHhSfDn29QcyAEwVJ5QAa0axGNcA4KQPxj/oxuiNZYV1N0DDKzOTX2/K4DI6wgp
HajwGnCH4Q9ocZ6vUnJEfuCmYbqG11qYLb9i0G4emXDCdm4TVsG4jDcN1pktqHg417C/5XMGkXHr
3Wjol+P6Ed1vgNgjevwMuZguSdAc0SOYyP0qfV/3vxmShdYdkTGkqYCjVESYN3tSONriJ59boKGn
YqCnqNbES8hNrczIhJ9PuHT8o76mDTNXVRCz7gJjZZtDEqWh/srWERzzJ0be9rw1P0eIQWatRJiI
fIHGJD21159SRoPnaIPpkbxMqxDJ+18UBkOYDK1cvvLYg0YHszAtkzwrZVAz7HLVjv7PWCChBTXt
HcV8GolQhrKQD56+m3kZFBynYwfZ9cW55bZB/SUH3vCl+1jhCVk+CR/IJvWQeWvFWhjzsanbwiSi
dDD1fttPR8K6MnWsrX289SiYdiMs/opclvq636DOboyRNkzDyU78MmRiZ+/sNDfWM4mXFbYjUr/o
4Nn5tPfXREAvVkGhjTaFqhGmw2Ytr8QZFhiAY3hEcvz4Zjvy76/Jilt7RKoLKWZWINvbAi63wI+4
N24d/clqP6clRzgTQ6CtHmgyCQjyn8dKu7+sqMDZjrymIHKqctlP4Nw1+qx6PlwTUzI48u9wx/x0
6XS44wHBGhOl0MR6cung0twzsdgY6tSNdoNHhRono+J+sBQeWzTaxokg3CqysWJCntIJeNEqd4DN
gEm1o3giWCgYNOIKGVKptf4+dokQpjxAri6D0Saqp8gbOfFe5o9vRaKiXJal6dwK6nGzss8LQ9Cf
8p+8Aqd3YtHEXcB9ZiTxZUDJniqc8/KhcrUZbXDmegtnj8jfx7XuPSE98xQEWoY1bbegZKstuSmL
Z7d9DMdKGk1kzuZRgiwHYhgxKHoWYoP+A7CbBwPsWMtGikeodHjCu1DzKT0G33Ji85paig0xl3Qz
tzbO3Y8mpRhCEf3BIdlL+QfFjG3LqewNukaoM03WxMI7g/KTHXmbr+fKA/0sO6QQIcvrE4ZiCxnI
ONzw7s44cCk/j0xi7ntDl+IJw8yfmnvx3PNBHOfltsJ+OGsSTa7L83qPr5q6bJvydm83EbQOMHp0
Gl8CYxBDN8T3yCFCCzyuHVpP67tprpOoIw44hMkXygZGQAu1k2MifGZclujB/4BkGCmruuStjEp+
N+tQXAlLaimdrazIgEbPP34GOH0UPN+XXMCXqjPwz5qbBgv2ZFvCeVVOk2g0+ijlYR71wV3Ja/al
nlP7SHIK63O8lPEVLgj3mfwbRdSDSeyAW3fxUEYNF3oEguPcZOfYGyE8+BPIDIz43rpTtdkiO2qj
DQCOxVIK27lwnQyLjjkThp1nHuMtAGdRcG9DqjEj+gdQG/ha5R63TE88XY8Cg9uvfW7zbpqZqdAM
XYIfK5w/tdGvW0AFmoVuWXCJeZuCrj5PdqMpydkkzXeqIJOzaGoIqNY7r9L9MCLCG5h7tiyoBiF7
SXv46WXtE5BcLmTzev161uR8ZsONmvNNF90sMfTE+ryUBwPnmnGsW8JX7PK0CXfZoaraubUEcDKN
92U8PfytIz/MevT/i6DjHsS8i65O9lqxHsZlo8lGBZ7knzu9N0EtM0TJonyDoU7hvdLzblVSsy3o
PrtPtCeCpwWKMPusqvVwkh4Z03SfqFuHhCZnJly65fw+vCb/wuJpIbusJ81nGW0XEvBsvINyvo6M
dXU1CNXxtIvSqoj+SdmIqiCmMtpNPnaURCohJETNH0Oxk1YvMi/dj1PoFqw9kpfe7SL6qaniQMc4
MV7bmlaCutzuNEMiy0dpJlpv6YhNj/d1CnozaZRYgp1m8x4qSyKJ35vNLCNpIrdeeZWAcj3UvzyG
9/ohD7BA6ge53K9qLjTDZceXJzLnu34QnF4RT47VVm/3odGqKR7jqMumdO2PfL/HWsUMObFmXSlt
fzzBiaApXHrINcWawz5a4H0+qf/KzwN45g6DvNZA2pZ+zYyfJlPVDrVeiALpqH0QiZyPhxyVtn0c
DoXeTirrYF8PinWfYx/8e9MM9XhgfraHINEL3uBmhmUpH4Pm0rB+E+Sw+4Fh3UTHHXBWwXnQONXh
E6Y8ixZL7koSmE/Kg4PBnzMtxjWrmkACAiguSOLMVcPi+O1dE8iEv8btRCvlQRjA/8Mcl89H0i2r
86x8AAmet5kikkVEUtDaJHsxjUjuBWNlnUCQyEW91ZsxwruLQt81YgXSdqt45hlY8trXXx7hIscD
hqYj7xZcmPHNZJIcKnVdgofFKu3cZ6PvJAKORFzDQXXJtud5fv/eGRvgOPiL0dupIwHt5LbrgoFb
cNMSutoBOAJDaIlJ0yNl3OlRFGLI72qZAX0wSaUyozn5Vfj15PtVt1EzBa4dEKuGOH4V5z2ei+Tp
oT9uOq4w1UQOZX8lIKf+PRhIk5pvod3u7DdQiH5gVKnV1IaweGg6Y65MIqyWYh0cNRJatzO8q6wF
Bmr2dqc1bxemFCg/fuoLAM5ObGjEL2gjHVXfyCj5aVGHPuSfonG05OsoKsmeRVlDQC1mcsacPdIE
X7FrPbB9y4WNsw6Ovg3C+ZAiwJLXaUel5c2l6oi7D5BgU30iiTAskPYSg7+HfZwaGNPPgcptCggr
9vDz60uEvMIWgV1oDdRbLst6XkCOsPIODZRSBElE3tbCFShxg7Cy7EKLd6UXMzRaqgwnxQq96Xe4
sJG7Q3K0OLhsdJHbzwNDhvQgT8ZHs2lDxOApWfzw535ag3IrTe/+AeXrMiQG0Qwimz4yZsV81sBu
6379/e87eCASU35vZ1QO9UgeXyBIE/CIrYP3pIBqZt+sxlkRZ7UQA/Hv4wgeDddyn8rC5ZN3D+JC
a1PzBcihqAudXx5lINgXSuusa2MyFgAXtXRGoAMSAv0ihaGZMmJiQvUBSrsgLRdIjlOpw5Po/5zf
j3MUaAe1EsLOq+rv0EPR7I9oQCVAXTqPIKaFHMxuNlXOWea/blCYlwM1LMaABDZ2lXmNVWUvfcDA
fy+LmSKZrYxdBO1q8EKpAc72nb8iLa27YxfQIURVJ6zR8+dZmrcWDoWhltYKSqX6GYeCWIBWlxea
51RT//FDiqJkpJUzj52KeI8O/EW6P48tr0rlHDh/VOZg8MpuMI/mHEEEI/LBKE4w4DrJ4bwLBUQ6
Y1Gn5PPr7/549IxCrqGPAYaRpHOe3aiTBsoO0k0yw2yc+cT970iaQB6TftnZKXpmGGY2mAc+Mcm3
VCvbEs4mM2i+U5ztlwWILUSVWtikAnoRQJa7ZrszA/zABWVj+3O9ItNfKRYK5ss5isjToi0r4303
s9z/VLB761NqPu0DiLYY29W+coXs0/3Gl6b9O0bvgRYe5450JxfvAlmR3FL6NZVZbn/TyjgxljBC
Y0gjwN4jpiti6wvyOBrNk+eA/ynYb9zbMFZ4xWSvK1c+fbqGKjuFTLkGZeVcmo/fp4BsBlJbDAWz
S8awFVsO7P0pKkJN0pJV0WmpCqcUCGZelMXw2LG8yG/5EFsUeULVXr+hoIjU2AIa83ABVJyoBMxB
A1yNgCPfLqHUUun6VqiPo9A1ILLZ7ACg00XuwzzjTSUaONRnOswsGDzCf6Ol0or9djsobrpTBChw
dHkeudpeYGfZG4eL7H4An2iYWduVUs3iVV19tmJNANlZBUFManfkTgCKjOc1ZBrEFnXVvTlSF7bC
gxUIg7b/kXVR/qZocA6Log3wSBFEkRow14+MLxUa9xELZoWPqBbyQ1+Y8bhk8KPizuXvYg3EhjEA
CjYmOG1Hf9FuPF9UKC4L2L+W0Luh3FOicXzMzo856Uof40WGiw0DYtiw2w9o2jQItEoPzQJEnM37
RGEFLzDdX/JpJb3QLXxpjS8/RQ2WkCkeX/7tEFNFdkhW95Xi47pe/SMW8Euh3wlmvr4qq+e8nGlv
ppOKCaWovLXncjYpN+zZxeJKjxqP5AYbPYS2uA+Cx9iupn7wTt3FUJZa0ZKxWgQaiMaIdlxwLM2l
fnumybBulU9G4ae3USYz9as721DfHLO2kS9nBakPdZ74H0Ovt0Dz6Dn+S0XzGYpggUZYDeQf/vN0
CqWsyKW/ufXItMysCaEG54TpTTbS7uwLNsB5b2QZH0RQAw8VK9neqSHv/PxCCjH0p31ne3+fP3Rv
3UTJnr98EaJGIkmGoDkLn8FOZ6p5qFkRH7PIBZ2WXr6b9VO71gzI6HcSt5IQzmbgfaVG9Xhcm9S2
i6Tsn0rivGXIiGToAPelvTB7RCIRhSCLBEFxGBUceks21Rs8lamK0BWuxYmGQaMsUr+rJmjl2nAb
HO8k7/IgemI4suNqejl7EcB5Db7GGkx6NKQPA/2xSVIuVitSRaf0B42pfXap1SGatnPY5RsnBYTI
Fr38vU+2HosT6XQ9wo+6igHrhd1REYvPq56xMIRImJaMJ37MPaShaQvL5brAlhYXDyIU1KAaC/k6
OyFLkR6uMh2vLc5BGeX6+p1vWhPmv0XHhJ6IeYu383EiEF9OAYoCWAhnnt25IFVfGcVdE8gzww2H
zoS7X1lM+IASZJUHHF+qREBEOSP4uk1fBAdoF9HC35V2h2b4wSCxtsQLa88gYlH4XOv+/dP4SECa
b2G8kiaRDLAO9MHBYqdj9h8KkB4OvHDtdNgDxEUzUsU9wagriTW2RDat7xWuBOelhd44u0PZyVzr
Sr//ahfItm94gcGsvMtA5iBme9uYUHNFZzMg4W+NROJTUbfpI7TuzznjAnR+Y/bwcAs2m3n2Jkon
JdNW8cLLT5IsoQLy9RcxYys+Si/Xao7e3/uw7OVMhg2XfWa/g8iwR3IaIpVNMTVXZENzl/cW6ml5
9lcaJMcSymnpJ9WHJV4FyuJrkF0+ZEAwoZ2CW+1qgARu5W+zmL4QItD4eyUYGP9tpmVWfyA3KKzS
bXOGpM77qbbKrlne4oOHNglK92t4wMV0XLMJYejvqCEUu9LJfpxUmz/ACpAcXI0du3pZjXxjoepO
rZHWVR0SDYhjFVLsGP9LB6cHuhzs+W1UIpNfjRg2/v7BHPpOObTbKC+/HlZSKquaQHhMZGTukhtz
W3hnneg+0fbo8ZFmVsUG7+7vXePhz9X888G4rOu8qm/EWYnLsJZWhovGBXvmC+5Wxs0VKeCkF8Be
bqLhDimRSzPV7g6RtZDUdDJnP0i2pkkpblE0Z185qUAXENqqCqD9JBNDfjr+Zp+3hbupEbxG9tNH
BpzAlNlb71wO6HPQmagVDfF7P9DVP+RbPcu1XnlF/5CzOcULFrii9N6Zc10eM16BCJl5eoaUiemO
15zG8N3VBAy+FwrJRswkrxE3LBfLBpD1jbBfmZSZlvvBO3YU5N6qz4VCyv0c31WqsGyFWDToRj52
ld9K7nVY47V75BqrG/JgQJ5Jm201s/0QELyaTeIcQkuJWZSqfhbDLLdFEPS+gj4QTxqcp9Zvilhw
WLB3w34Gs/blOVSGyb6ym8W4P8kGjUYqShNbWG15kq/avOSdzv6+rQQ35YAqcI2TRLkOYU1/1uPR
cCFL+O8TidBJH2wi2/YufkGm0eNNmP/cw5V/NRucMC/H8XLU+P5Jjk1o+ZVUvyeGOj+w0XRQ2SNp
YUqsqK+3jOUYRCa90xbS/Y/V8rokuXkQ+PXVJ4dYeVecXgpeLbfRoSOYUtfAIH13p4KgYKSmXMbo
0zu0MH20KkhhpGVNhClsL5AJmQm3hy5WqWuzmWC5e9kTg2QbCZsT5e4Zz2Zyflah999z7xDY6a/8
niiQZx1XJKnb9iF6TwdW/9e/OeSLqfbAzpOYqE23+T9q5M1vnUJ28ac5ZcrjRFo5N+OTuvSgMp4P
dte03ZA9dNA2hru5KINWn9mHuH/JlHAI5lRD70JoM3Pp3KQybIsZnVgvyg+uL5+jiX3sKJScCaoI
bmJP4s9q+bnTAPLL1Dg7trox75C7gfXKyJKRtyZk2gNiyWlvJfY/WXSXo1voY5i92xLEYU0iHJZ7
2og9uc6othE8zW094v0ucdKQ3yVCKI9MEyWV89skN+9skMsibp6kj5q2GXWcJ3K3UBjl2AFmeSSJ
nvBtQIR0v5aH+UpQdfGiYxu5RRLKs7GIBlalmIKpeNU6gPM906ZG/KUHnwTLsXSJEab7y/hw+gZr
MSaiopoF1lNuDXXqq+8eR5MyD/pdf515W3zs7ifDSu2UFIXatl1yFJkvOE4tNE+QWuyZlESWtsK7
rk8Gr3bp0MftrJIqda3mBLWmmyuRsYNld/Dgof5DHXBE2tMA86y4k7m/fbIGejUKoi7tgbXHsTqO
iD6Fj1w7MllhvaRRu891m6Ju+9OhfVWf9Y3m2IZtDXyOWnF8Y5HiLx2W/2Ek5uoXfRcdDuevv8UC
WBZdtJhMMBDzdbcezYCAZ90u2xA7XargJz0VVjTZS6lwaCP4G6VEMwYkcjC6EmmwUaAnxGBqhB+u
MoeaGAo9OxixyyGHMv0b84VLaly8eMhGuIbMieA8OXx6NKtpJ5f+xQ3W7ssDvt7gcR41tXtG0F6J
9LbuVsRNCwqr/VbunoGcZG+JPdspXMghG3Irx1nFYJBOYBuIAUKnoTq8NqdU25vkwJRro75MKkx0
Bc9hYqPNV9qLiJVpaLJjOe72Q0Tkd5EZUWY8u6sojCsZ9Dt7wW7c1/F//OtN/x5X9ccR/bzO+LJh
bwug7U75HBP+Zr2WYJDeS3wtf2uWhDR4p0hPaNn35XZYXPyD2Od/aYbFbQOGM0QlAHJYmMTaZZYu
V0yprmqwI+wESUSqT4Sx6RSZ8qXoefvF9QQjOhBmfsVMEOvKvxKafR4TfWqWhQ3RPRGSswdizgSc
hWu94aRX7GZc6Hc/hkahoSScFw+OCVSPgJr/C4pLHxt/QQNYQuWf9qWRG5NcUvzQwwOTZCEM9H9f
E9Gsi+NMIPdjoeWOyYTnksR+HgsiaOR01PWUdGNKLsUK+dYhK8CoEG1Hvebe/AqE82SRkw1U0m0T
EH3uJrFDA/YCjP4C3SMm58SatxpC+j3ZcLigtEDxS/24OI+JHlS/YRAYvy+2O3CB94JwyXLbLuAP
Ar/42a6WPWKdERkhq2cbn+bbkthICURbs/pBo9oH5RTops4Bw41PhjbfInjj2CpfrWbQwTdh2V8Z
xVAU2DxvIK4lHse9ijxKIMl/WuBDFYkR6bx3fRbKEfKd6tiApXMIXN7djpZN8cdoD5Vh5Bgivo5X
0x2wWyVwAwiBt22T4kCnj8CLmPaWTPIhhCAi29UaNSyBd0s7Lmc7FiByEUODtr3mu5TQm6ABXo5R
bWDJFbMYNOucGikZrwXDiknfkAkcdQvL1qOOq0n/tRickMPZGW0Zty7YK7tAKc2FmxD3bwW/jsOw
TLyaNa3zGceOG1QB5k8XUpsvKJhrzwYlDXi4TU5pt4KqrRrbRDzuC2yBzjUeJxO+9MmQ/EPCMLf1
YVJSCxftF94t2zm6/HB40JB4j2hP8fSonhSNRyERBEr0eN+PXIv3unD/PPXAnVaIINcP+vVLTf64
Z2HqmOm9XpMt0LMkS1Cf8lo85QJTQmd1rMhspyofCv20D1G05rw+URE0FFeNYoX90V7ip5WEZZ2t
xV6fA0qbX4LyzuFUHQjW/akkPa3KJpJv66QpW6ltWtW0vns6FCdd41VXUduUtQaXW/3v0frf9snf
Yk858PYzib9lM58Luh2Ceodurmp4QHmRN+9UXi7kFeG8MxYTUYRF4meXU1YNipIA3k28XvmoalQb
ERgQ3d9iebXfK/WIloPTIOsWfpNBq5LZG1geuof8F6hME3dacJMOyOnTuzCrXwKoe/VMxdMQP2lL
bsi/Qrf7xALj4Y4r1H2IHD3ZsAM4dBbKcL2HjAZw88pnCQHUrUWqkjxVhs+mq8GWNtjT7d1j9jFp
3jzGADNWF6x6DxjghCXLbt9s39viEziWdFrAPRNNzpQ/OF/ks+qcYArlxyTX7dFkmKHIJdGAWsqA
thH2Mnq+BjJMFUQY8glen6X2EIrFwam7tnS4bYdbl68VwNPIDNkJdoL8YkL5IhtARNpR9p1/fjZo
Bb9F2PvWTEbVSbpS8hpLTiwe6p/tp/vr9pkDcpjfVVGsBU1hyWX3lYDlb49sfJRskEpX2oSYC1wh
PFNSL1Ts/H2e57uUNZ3Z92BpH69B54tRefjzXWoS8AcjA1ac/a6qgvnkbvnzV1Ml4/DRrV+i1XLR
PsY6eB/q9Ax49zZmPG65YalpISeZOXm2Ep7h/5BWAUOvXjlIcDC8swKk3NsGVSPL9ypSdCOjLs4K
v1M5kP9sSkXeNupUjSE4sCbE+Toefv0YInezIiJ9rHkLbImpMXVMqkokm/5sMG49htXxXIlIxqJE
5KJYC9xd7OYUw1RXs5FoaCkLW9SUzlTybyzaz98ylNLxbWcVkW32QIjr9INoEYyyumDeNr9O0Ciu
ZBEYyxV32uIXMYKUg0Ml97l7vYOa5pfxtCe/FM4uYn2wRGAfD/cIXroWlaTws3JEylr09QxAutyg
c1fwvPuk0Y5+zEw0l99S/1PPbmM/dLLvkg2Yz4OG+M3q0XsxYJ9BkY2Nsn2sjo1JzvyAXRIeVSW/
lpk90bt0puiB6lWgZ+hBBHrwvkA1V7ddbVvWrBEbeY5ic8YnLHqFb4LWjX8xAidP4ZdYhBIQFASF
KTtmrzul8xJLoGVtwZyeLXsgTpM9xYtjphIX36nCKZNCMMvEUIFWooo9LHbrs5DNsGArI3ZAccfD
kzAEfNnCx8Nzd8DEa1t7vy9dqgTQooAgj4rL09/pRe1VIlSv6KwRyHcfKxygxALPzXE/IzgHuP1P
crN7A6V+/B+W5luv+LbZYD8c4tl869YAFnwsj8yAKuxUcx4Zbt2OqlhWJz2Wcov5dO5oiW/TkkcB
8NGV3ryZyfwCcNhO/oD23IT7uJgXQ/Y/d+R4Pw5JuR7Xa01UOxCYIDn6lE1gtS8D03ORjdu2u+oi
KpaGtxWjKXjpTAI18tvk7pnhWJf5/kmcYRnktwsbUBTXnNDQUCCdqA8mHLItxhqkdcwLDRrT1c8T
GyWMX/YntYg0RVZCnYszXNp+kzxdvBjqDmksshY1pc1XCzGeg1oRTnCGa8iom1WyxtdQdiYMkXeN
eCf3np9a+thw0NK6a/2iGcfXQbo5YPE3LuP4xnVWcEOJ9haKRiv6QNEW4GwbenkvVHMGkDDhEmFc
7V/SBjRYk/Znr3hwdbaN8tQjdeyGNfLUD5Ss1OjB4XNfF+wTSIyGmspiBE/6u83LzJzg/UBapBHj
wzPZEG6uz0kXhYehkr3wv2oNBK/RaooTqtOAQBSHImGYbqJi+AykuLCNhRsx/JlHRgQEzDX/Dnzp
dO0rnEZ3Y2QaerTCx1xAEI4HPa4rv0bmayzB+979ETYWQXzKBWEaRF1llvQ6ULS287A82B0pcb61
ZvCCIuGvl/CNjzYC7Fwnol/FkvnVd6oc+W3fvanh92yH//P0gzSMcg7DhtTr0HZc7bkVvNvslrPa
bWqWyg8zlynzcKfq7b/R2r6PHVGyMhx/FNxPLcYLLsxgGbMpy6u5kQ1KqkZpRTbQimkPnriW/VIM
yJ0yv/MCZuH1R8vttwhN+UPPhMSjmN0+SCtQl0WRfclDj6x2mWO2g9WaO8KaSjhrUa3p/OClAb/g
eSrddd48yIlv0DRu/xzLN7+YKSXfvDeuqto2w1PZ3/v26a5ARzRrr1/QQ69yK1Db2TjCVX/duR9l
a0v66kjVcbLGvEURs1bZU0X5pTOHwAWK2Hj28rucHm3IdL+BhH5bykDOIBlQbnGGD5V5H52R2fny
t0Odra/LsFmynkuiCUWNvZim0S82sK2vMR67B0kmIzfrgZXwOfDwyhyOK7ntmcpabS9kvvhbkJt4
xm236lpEVDjOzdnlrzBJi3tp4ZgxXraxTVwYulHWHGYBnXtUNrG9dkGyBkiRibI4uz1Oeq3RGGpQ
ugXEFZAvDuH+EUA8G83Ot64RkIctMH3HiZXOYLRs2i23PIZzGUSlPJFoKx3XFA33ZkuSVO6cH722
GUANb07ErMpjrTKZ3EkBlA8l8LntsnOva5CVIRO9qmNqQurSAsbNFbXekJ9UoDINpQXVsp+KPjL9
RRsWG7vBFcLWFFxSCVKFgtPJ9n6bxG1UKO+2tq/3KIPXO1h3GBzVzrBzFR38R3dFiubqzKagwEjA
I/qUygmOP0xG3l6K8lp76zpKuh6fUK7KdumGseurLnWcR4+eOuRrQn4efwyBHea1ND0PFk3U864F
qZMPTcX0uFMurgTGBnGS9rUYwnMIwPG8KOaRJ6YbXwColRRyRklCxmpsmdaLUsUcjMv0mdFMLTf4
lLM7OWs91BPBkEIzXy2XCbgxNBj52wnNEQJNsd/14l2ekby6jrHohiHvbDzbIj+To54m/Z3KTWK4
c5OnRMKNSv7wIfC968o5FrCZjWI0vrTLqWt11pJ/4PHRTd1zXjGvxr5SbAiSUYpBBighxV9Y81le
O5Djh+7V871EC7S73/Yn76npV8AtLdEs16oUNpUuXvkUK/54qThTGbPpzLvX6jyWBIxPXraHme2E
xkl8/xR/HT1KO/LcZE3RPo+2Gxm8SunRjGzSX1EnmEwseYOojsO1YTOtnA5h7gFhhVs2x0Sh7u75
KyH20HMcR6lUGuHm1nBgnYy2o2/02A7oSEx+Yjy+cupSrkxRSqnJ+3yJBIVrhs/nZTAL+GIDXP4y
uZGLJPCubj0Mge2Gb2x+/Ey1enE3uk4PdDqRNqC0xNA3LXTbIoiUDWpPVMMbPo133/2Hxli7YOHS
GNlAysgxuhSpMGZYn7C1mt93tE5btDXhly57mZ+LrzqRxOLfKWrdzngFZNF0sFEDZfkJfDVH4IAB
nvyt2Afy2MnK0BZj3GTOsJw7EmPO7hC0thY0GFe0fyaipfFRpn1Ha+OvIptA+zXcMsIpXPZaSJwr
25OY7AB84O0KqrhsM6vBy/lu66yVYo/dlzHq9jwauQUh5Bb68sht1rVvJ/xeSHIzcfopEwZpz1NL
ndUN3NNFCndGBAwJ75lE5a7rh79J5yhhdL9ITDAsGvQFoLN38cc4842yNJj0LPIEM/VXKNWiggNH
1ZAHto1GLcpLw+4qWOlXYJZNuYt+DhAs1oKzE4g7MNNWCXf1xfv+smDRHf6ZfqX9urEBU1zGM7Zq
SqBefofDzzrgwTzcOEatkXGaKF/Qmiff8akX8Gu8gtFzFrezJmVorORAciMjdgY71OIIpXesMdGT
HXFnz9/vwEYAaDQCgLIgf7/cehM0r/EZs5mGBpNyDGru8FJR+S+majLhR7E/u8D07ovBGBUiwPP1
lcEVxDhM90GiQKIE1eObb+9ikPq4TSoBUD+K2uuva99TYmLiLqVRgS/s2KWId8GJmwWV27kD7XWg
c03CmWMTp1SAHj1dho9z/iHv91Dp4GPfAmECCTQ0aHP2GDoyEyZNoNwpO3LsL6eUTRXY/cJWppM4
SzLlAtE6sNdMW3j/eIHeLRp64nSihNcfw5271U6BTjqb/wx9Krzbalc4BrPrledICRDZNpg7BAvB
dCU1y7pEVTMW5czflEoHXHZCn93BIgC6GA3BRJJBx8PftQ0iOG5pk0CTt5ViGLhH6AF8JcNU8ImX
FMfxLXIKppu4XQMAkbdjVM5/OkocvM5MluNZ90kzvSgSpR9a6rzL9mwH2vTSvCY5mKWa3MRjNOWL
4L1IO3TwXAzxykfAjYiVFlMBkJpIyX1D6kl5IkhnVuwdJwRpdU1Ps15M99kruJAaCJClH37bFx9q
4n3VwK/T6cyTkkZaymVdx+2iTd72Fawd8MEJfPb2ZMvP/eWnFW3DniGAnnB1ehWXH4kwAzUTA6bg
4Do32nNHe2G4qgQmW5kLKonbU3qY8uskm9+L08ugT/0eNgmdMIZu3oOfNVNnr5ygAF98V0k8hMn5
oPV77bJPR0isnevAVbcRb+5pA3y7rLdfHt+Tage4FKZUW5kLd4tzc/wesl7G1Q8/f2loZbVuEuVI
RrdN+imjL6eWhZ5Abir75y5nY6S+al3fvmDF+mNAoz3ksQoIOKDlUBRbBdvsJq7yPL1axBP+ODZj
V3fPuwO/1SHWVrwYE+BCmA3rRtp6RTSggWpEx93GhKSNNNqTL3+FGd6Hjk8mObWrO6gj5HMteTTS
5ew37ZBAVDoM32rsBoaNyO0zJE/v1f+WChHEobrj+xZJRcdB2k2eId4/DSwLvvxE46PSFAQTSDDV
ZebwzApQW9nDDg+B964G6K7ozEh1BDoaPfi944bIBIi+QpVRFW8sJLy8oeblh7yt/UHWDDZGlUZ7
6nuGmhhx4BbQW7UNIL2iSA5Oj1SG5YaYq2evvACXwslYdzO69Q3U9PMHZemCrZXXmo7yoqUbR6Uj
8pFljtsuoOsBN7sqgzLt5WMSZsy/wYBrn5c7ryc5QGFO3Grw0X0ASXep3MdM9YS97Tc7KqtOTI/s
RYDs2e9qUgp7xBQfY2UZkC9gqDJUtxQyXjM6xZBm49dTHzaQK7oEIxD5rF0y+aGDgh+dnbv+YfpN
Xt2KdhtWAVI0AMvaH1N+9ej+V/FYkGndHADsYbz7dk3mJoZvQC26+MSs9LARntHQsPcY1lz4LbX6
X9Vxn7WGhmLZCfV4o/zmb1YvgsP8OPqsbK8Sy7TAkX/rVDw0B3CTus6ektlcIYGVdPetCBVug0gX
TRqCUjNxJzlKGmU/IplDJRajHs2xD0lGr/U5UsrQTIw0Ty6zFnbCYSpzBmWDmLazwHkNZs+BvomE
tFP56aJxRoMqoJO2Hnhh2VWI+F6OmFB4aZuYuxP57XHf7eILFdTA4CgSIeMf8GhF+qG3jWB2cJYx
cSPtoMSXms5LU84GLliinaR5a4ZIsUKtiKcGaVY0m/iu0miVmUCE6zrf+daSMwqmrvCxRZlJ2ue9
v7ijnTrD5FDU+L05/zaBnKH8Uq8qiwHZMaWRH4YHwwd5CIeyWKpGLgq1RpMBJkxaYaTI/FN3coU5
l/mCv97asv89B/RT2D/jLvTow5LS8R+6AcOClPJzkikqs0CyUqy7g+WH6Ha6SHGidyhZDRBgoMjN
ZoN39qJ6/COfLuTllEIvliXwQT4ztDJ7EpAsw/yXEfUqrzFAgr7Y0HmiKbRarthBpQW6YrYSxJce
hfQVQKOCDPiIPqlk4ld/m7fkmPu1aEiGPgzEbuIryIRHk9TLoC8mcEFXsaNTO1WTAtiDv53LRCBf
efaN0DdL6PZvkFdnDYXoJ/9HFleAfb48KKF6XXyLw20ua9c3gHq2mPjemJtCJELPay5J/8oK1r9C
1XrjqEpdR3iBFCu5ZSo3XBrLr4Rbh+tygpdCX39bnjyyEI55VKWZMmqiDO2PuKmsl5ws7Zjhq7wn
yPVnZ/bnx2ZWWmCt0/UPvmRfzguiGgoYAwmM4CuWHsB+pVEIxB877LphpqdOlINS8WhsiLqg+htu
Gq3MTXsKqiJVWSef10k2ZizU40UDy5as3STvh/ytUDkYe8H71Kzt3PKPVn6+TCu24Gi4YmlDSdKs
vkCPb0+FykKobex24iTBOAwB1Riord1PJEAgxS8hFkHKn42It76BOKBv7bVI1E6rwHuwZWSs59Ml
8HApwaxa3YgSeHrkb1qAFTqroB61en5qcKWvguIe6fd0dwxy/s1iipERYgkoaH6ZmEmx3UEi5JIW
VopIHeeEueodhklEg49XZWOABCdI0DMaz/mXgVra0T+TAuNWGXB00lO6o8yNOJsV8nNJig7Fju6V
ZAwR65it0RmIh4fXqU4Jc9bKNj8CSCVGZTjrqKrRDJZT2myE1DMdW/IzLk7UKP1LxJlwkeYjHKVo
rNF7mXa33IB3huEIDHTsgF0by1wBvlBAv8CyzjNdNsrjYx2Zph2O8ElTaYqV/OaknRhp/cOpk/14
LxCxogX+6R4HMq5yV8Im58QpGEWzGZ8kxLrMRw5M1w7F5hJcsV5O0iLCtC1UmrDbC+wLD1xEugC2
LGUg/gVq6V0GZbl6hDNZ7OWD6NdKA5OC653CSDNED3O7bXy3d+ii2KXJ8iEDqYvxAM2ErFwyB877
xuticQ2yEytgmUW2qSDR5ZV1/fMzGDa/nPFd1HOVvLFsvGZprkPqAe4nAB91ueQLc9S0pgShGj6C
wQllZjf8xNB7dwLK9eXu40/M9CqCLhx7+jjPkRgIrZ0/TJT7axvVsWEfnKUclpBR1i5RWRYK6Khe
nq/j7qJhkpwo+nFY2IbnKnwanm7HPcsNj868ntxlQKN7WZn0LvC7H5PrIfU4C+TLQm4emYhTjg7X
OsP6p9ZI6Fg+Vk6IWNDgsF2BBks5mNGIV3gPl8iGq/vDaLtFcHzl019G7Sa+0NlAmt8dz7ILoELJ
on+5jq1hEYNv2smd13jdy8R4yWoupHk2W2V4jearoQK/WNJKHq/JY+oImvCz9Lw5VjnTE8nrLZS4
0v1345jODjZ964vh9T0y7YHDGVJpoXcO6omCMlE0IIZGSLyZMQcfQ8E/Gwgv+0bbsT7SJSqP+UpS
+vosyteqcf6VC6CQZ4PUgLLb75icpzcyHH3SB7U2124/t8IWjCiMr0fPsXmee0c91BsB7b2jq8d/
tdysEA74EidF5bswDpnCzgax++Q4seau3lc05H11AUfj+UkUPgNfeve4+2F9ygI93ldDRmZFBTiU
gitOiTeXEkJOlyb70EqoVre3RsshCDw6YD/Wun1yoNAMx9638YGj2sbOj0whTa+p7ZjDrcUu4Frs
8Z2LBB2IsSLl7HCBjhmU5xmwWzVXoh4VJCgZhaa5z6jMba65T5nLA2uYrF1218v6JdjUf6jZGU5k
nVyV3DiJ6WQdlj2PNimPV8Hyr8ja77p0QRvK8UDnYwkK5oQ5nyZHVJjBcrIp2XQCJOXyrsYMqbt2
rqefm0I9y92Og78V2+C8H5sBIOqkE1vZU062eK4mQFjI1ZSPQ3+PSE0WBidkNIjBB/FxVmEV+VH1
TpJEv1KkeYSrjGRq6mPKepNh/VMVXZocG2VjtwGPZhOuUFaMaAt6AHYrTSkVSAxHwPBxX6kkuwsK
oeyGKkTb196HcsgrUt/+4XaTpk2yMOHdAn0E0lcLiTv+XAhGqMRjoQrQ7wNZZvkrM8n8ywJtjrLi
mv1zmvdBTU5K9z6fRJL0DjZuRxVnDGCvKsw6tQxmdE4L3cQV1TlzgzpSTFhnpbySfOJk8XsPnjfO
4O+k5SaO6uiFPj31gMmExGa5Zz82Nt2IFZFhRxNhfnfWjnU3NWteahsHA+MWdZP0M4XD952mvlDV
5cXaaUc1kNk+9r8kRIQe1LsBiUo/KBiaZbqKBDM80nGzEEsiCzpGMt92dUOM6251Ezh7+SPuqY3H
zKxmnKGznHyj/K3UmjFh7ooWcnRTa88LJ344Qyie2BwDOAVYGHHMmM4e7pbT4PQJNxS/HgB1aAet
uNPKFFRQ9XNbdkm4n9wysuBhTB9HUqXCih/cI+oTe30TshrPnbPv485VvDCmUaVzSYxPbaMlxkMM
9HiadGjPHaoj24c1xcacVti5/640GBe9QqIP5SW4Th7Dhjm7dI7F9vYAz+rAFYUZIzaCcHrnkzR+
Ar944246EI9hnUDgGxu7SkYuH+1QUiZtyshp55nOsEY2ka/3JzHCLMbnYnggwZjCVljgwBy/7OTL
OEqkLEicJW8bY59wvKZkoGIJFeDwsq8y2147iWqDFvHaPOyRuRa8TCY5+6EOCn8lqTeqn/HyWr6E
WV85Ate2+51alb4Zuxr8O6Pp1Opx5VC3A2gJN6aNbO508umoQCPlEp7eTIWiIaBxw2VM4KfzslBQ
b4sFR1Dg9cdYbNRdxi/cBUTvAcL5bfP5qysq2jATnGxoerQOdHxVAsE4YbdTO/HxxYtWhJoYZGuD
pENFudOp2Zn4cnZIeizJs8CSPA44MOrwlW+9otifVPCnDPOWXJoGc7B/iW8dN8GOLDpIZk/STHZG
2Nig5hw2LY4THF7hHBqxIDPizfCWce+tXsuKoJ7NEDbq/gB/mnbBhb2gnMgc/OrVBghxDGRnVx3G
fSA8f4E/ghK1T4Qx/yHNHRJ/LD2A/mwiH6VVdSa0oOyrC6bz2VHIL2nD+JunN7++ipHtqaEPJAut
zw3+5I9mitEBYvLqyDK2BckBFpnTdPtHECzfJaujIk/6/Co2FzBh2xOPypmZsxxsnZOBb+UobNxS
CZMlvrAdSYMiY8M0nAh57qqgS/EXbmtHXFj3URqTPJA7cn4XUxnY/DKhJSJN1rY2GvkkA+TXvAze
n/CnLer2matZLkgl78k1p6JEkhCNYLxLktU9lfEWwFlKHrQKIdPX4y8aSu7G/JugYpdHmmLCDEzp
NvjBOdHK/fOW1HhSw5676VNyXfK+SeSyCe4UlGoeI5alSyumvlI96wsUBytJAjO7AHyLckkCcDbX
wGMGaLPRc727BUbGRCtLV+SJ7PXSFLIyRJ6KGFauWTec15xXq/pmtiHpQHISf6l+rKD6du9+f1M/
rCqPlkO/wbhNBk0CZJ4bKyE6INaA+TEDxTbNXmUOPel32TySVmBhjmpphwR19qNyUrUm0aXkDu3z
ZHlBzhKycdCZxut7hXvxbZ92xxzaSMG1I9ywrMCfDSA/9qbWsA6QFKnsYqecrPunAWO2hSn56N+f
MH7CBEapQ2cRwBBSMJoWRc4IkN8RyI/Yd9uwCBiq80/rw7Y1e2Mh5EkhCOmQv5qKGdSuckIXdoqJ
i9xV5+z2V9Nyb5yRCdkdPmldCf1Acv1kbNtth7MJuq7YWaepkfXDWZVfjg2IQq/+p9zW/XqD2eRU
g+FHpglj0rUDSgzmd3iNJ5qisiBqvm7/WfJDqKLbt5R/pZOIhaC86ihOA18+KQwjtJA1t5TNq/p9
WLuDkw+cCNQZ1p8Q5YAUCvlS69NIgt9aO2fKhlFu3+FX3+mTll7/Q30NJWA9kQ/lFhkwfAFoxTCI
KFBrjbR9hpZkhh6CjKZMoWuQoqGOmEMeXhVLNzAXSRMUZDAXtq38HYWP5RT32Z7pXpqTRjoIHeOz
9ubqTbGUX8tV1jXq4f7j3GyzA3t0/OGtQ/z1tbZQBR3w3I0DXjKFvh3RG6oBkXHsXVijxiEiQ0s3
6YinhuBzK1PsqM0PqHsu/j7RPi8R9noLb6Jvm4GubID6OLQI6obHtDIEw7Ek5FhdbB4m8OOM+c7x
RZqoduLMDHABo7wgbb8oSSGT3pdf+Peb2x25x8D/dsPLmZP0vgyBgvHM1YscCvWcfLyzLicZgEZ/
BFZdkVbZgITKOl79jViRHAJXbaH2eciN08IRkFoHhYEWNOrtoLThICFSwQmcyKBnoUAgw1JyBhNN
JPIk0scIbm9aP80i28CGxKUwV2HCjBrl7ZLxPGDodg4XzpYyTR9GrTRs7LWdCQ35ZrpTI/cfpjfR
u4SD9+Vuzz+iYwFURgbxofgO7s8Ch9wATaVJGG50ej5bXBhGgzYdOJcnSgbPmVrHi3R8ByunWWMJ
0NYTYyQYIF6cJNCQ1w/8sfZ2qes3y37/8CU+KXxUS9b+RTVS4YERL0MCEaPVca5MdFjBD3ZDALXz
B8g91OeDJzZtc8e+DqtOEykqTW+T5OvLPb0GQnmEHy5Fc4EFSdAjzMtrwD5Z4xFXLSHWVAFf2Ygq
/F3RWUACwtCzDwB0HeDS/tTNoGzg1Hz0UGzHEUMVsSUxETgThPt8CExnVukzDlsZwCvrYcwFDj6H
nlCUgA8MOj/tgGRdIeGv4ZKxpLfp1CqZYDY0UU16SWDkGwXdBtleLAZ3z22+B0SrRes0P0O58g93
qur/fY8lsuncoAfTPnvFMFaOQmDi7VdY4H9U50bcVxgVVnvXQZhCIyWrU6238l35/FZvAO3F1mzc
he2yI7Gwfng/S1z2VgZAGklZqeJd6JhE3Faf7KGdFm2oKQ8ouTtHN87yajXOeVhlWvkVt9Fp8KsE
/0mFwR1CvCBIHpC3MpvwehnEP/YvbNgWh3bpFCzy5q4aMAqE+/pPtD3kM1tjGYOT4Rg9zj4Q8VZW
7xdTl08pUFY3BNBEFHxMyD9kYbZ+7vlN6EJCXa/TnaWFM2LGBPigbygV/JheLJ13exv8yRMIIiXF
04XooGtsgNzDZiDQUUF5HUOGFeah217m2Tv4Bxwirs15tHFDtBJiLPCLF4nwT3DyFN6kdNKuEAZ7
zCDUYiDEDIhHLQfyT6ImydzY7BWG59A8esdlNCZOJ8r51T/0PFfbhOmaB6dQUYG1JoWsYIJV5wyI
hFQwaMOaFMSIGumtnNdElDhWRY1lXoIcKa7XvCVrD77M1/yOfmYaqZQZYPwGT0dm62znoamzH/L7
LhJ0ZJv1MoP7Gc7CVDLfS0EbPUWWUeXwCjiVu/I3w3ffJW15OYxlShFsayWHS4eB5zeW87xaJ7j0
Pu9LjCuv4sZNFmtKeKFu3Jtkteg4ln0d6JRxGOySrII6ONMGYhfZS8MoXJ3EWDOMwX4vj25ApvOS
u1ZyGg8WbxjvFgCxV0cBdjH4LgVlABVMl/w6PKP1OKQ+qDi2PjT3UROd2s7W112CsYsO2H2llqVr
pqIQtSBlRZsIOCcRNsoLPSgUXVICl3nyz/geWQs2z+Yt3+E4Zte5b/fqRGR15QR/e+P7hlgbvgNo
8AgGYb8el7E95AsZS5Edy+82EgBwrNF1DKNui97fHrOeBhXNkksRvml62pbvH9jXURJP4V/WvJDR
FlTYd41QM7jqsiFc5581ZGqAXAKH5DFGABmv6C+ZAp9KbYXCBKHgwt2DYvhSgRqrigN1521lgpqo
w2sqXBrmKA/dYhgXBGcek7MiDPvtBsRyfReCyx6k/jZ1i9qTFPyEcx0CFzf6NMtK+qBtd5ZwSWqI
pvmOgMUNbjZ6voQosh8G+DFtgB43TMRwj12DRv6o7fGglNYarw2MHNH/2YwDX5MOCsSMhHFDnjNJ
Z6nPUIVdXtq+G+fKradjENjbC4GfJESR3SkdYxzF3yvLSAUsNsZGDH8V9eXJymYyhWLqmAYPACsI
+yo+2Oz9AYQhbyIBWphIO1VRRSIIxc1P0/wqnpED3TJz2FYMNzQDNa11jN3Ji3FFjbn+JuJn3aHp
tk8WB9kc78nnGNAH0K0Gy/JvafcdcGpAu6GzGGvme9oCbBRkspw42jtgddQvv/dlNJxIo7gKJM+r
7cKxAqAi3OBfT/l2LZ1qeuGWkhyowV+LR5c5B+zv9rwwrBQgGhgUGv0ap6XNeQkStezEQKiTCm5c
A+QiE1+bewI8j2jqNxRCW/JnXeRTivHMAw/aXfs9GDYbxuCLENXkm6S2EDakudcFTMdP2yhmuYau
2zzOUIiZa5Fu0sGRM1siWa+SCPlh/cO8Zzh8gAQpOjz7yO7ceuvXGDeOkRveoypdaEax4fOcDCEk
q5ggnIG5h1LBkhJNOb00CDg5PswT6G3g+JomdoF9by9CrmLznRtyv+bY7c+/y8VakUs90s6mzdnY
YK3Y990ZOn7DQOl04RW5BSdAz4Oe8Sf+dwC10bbVN+RJy82w5mNMy4WkRGRZe3pycTqd4AsGHXzX
0Tf7khAMIKREehGS/1N5hLnApshT1/TuTQKDBV3tekONALgKNwo7MpM6WduoBtrEVqFRVm3kme3t
00R52Z42Fi15tMASVQ5b+WxEQ4zBEEwJmg9+WyiduUGqSWit0fVrMN4lx0x9CB8BPMGOlgnWaKjW
3pVLeSGf8eySx8jeTq/ojgDmfchPGPO2vHjVzfeF4X4S/C36KGO9vLYSuz6fjghf1ok85ns1qaMH
YfF2vgizcVG5LSluDcNiljbwKOiBu1OTUJA/c3uaogGV0H6UJf+Xr2/LPBXumP84d5bQU9nGobgx
Mw12gbQOD/KQwNei5qMSDxEt97+zDi5sQ3KcS0yEiq7l6ztz0ay+W9Of0MX2yNyn7wGqkFyJuzJ5
QgocGpzGg6WV+VecHLFjm4+iRTz0vJzImKFYHhZYxcKwa/ockdw6Ev6nsXQCglZOVrL9TaGX4tVZ
ZQpnzeP93V0tANnZitHaLyQCjuR1PwmcTNM70DcG2P1xtjsPFPxw2q6/UDicx1wWa41R3YOkAN82
vK6N0DB18RgSiKoCBxNBqZpIQbDuleASIWhcFFSe/ukupCa0UIXCjJZt5sLMkWZgPV3M3hTPVDLP
qGDCr+yf262N/v7s+QwamN2xi+G6zXmdEluTHNL+chn0RqAN/HLnt519A6/5z2qKCFrMv5khDQRq
JlHcKrsBSuIYnGgBpCt4XWULNWiQ9HGz4/aVzuQk1ixMA+RM1E/QMiPvYMwLZfrIJ4696AqQhp+j
NezRVDejahugTHHtkrw6n30qmwTecRC6dqGqVDq/cbV75nXk2rWUv4yJTKabVwZaNvo+fRtieP9Q
GZfP9wiIi5xfe7uY4CzpSEzMgBNt2Dp2Prw1X5rgjwPilR0WtiiR1skK5b9KZh+tMbqPtU2pjPhZ
Xiv/Uo//+Dj4RdBRwEs4R7rwA/SCaK/Q2PL02i2s+ngPT6rkgY1Labd+Pl3soAIsOqjwIFH2HjeL
gWhTefXn2XSzTSBowIAqdySkd4MaA5pC4+4aB1+wI0l5T3YsqPkez1N9NnFXgPXSlPyCE0keg83b
FeulNp4oTr7Cf5rqZtBs1VV/osI0/nE2UJr7U4Cf/vx4pZ0EBQCH6Z+0O4VQ+muH7w4EluvHlZc7
Spo2EdDNAK7527/6LoD4khq+DkQebWZwifC1nQBr1SsBP4x9srcrSnyA6hOeBvipkALZuu/yU7d7
nmxIMDaiEjYzHsjNIKnClW/yVh/udsA+Ebj7D0DjMo6ZtMc90NDowep083QQ5CCjfGZFfoyAewNI
zCxzcCcyixLl8z5JDjcQ/KAglt2DFZhV0Oepgqc8mzA6O+akleSyNC2LAH2TKsie0DRXFmg/2o/v
ur75GVUkFlhRdZuUvKxu4aOAzRxibr4EowllHJmYJVW5zIbSAkXIMcxKxhS+/ZEhX5pCB9ktV8ga
t1x49s8Ck+Mzp0p3XVGZt0YfDqscnlQKhjarkFZNqY8Mx3d3tMrm9sVg6wbjR2utRuhMjpzWdJ4s
OH237uWSFBfbPSfquAv5cm8YOeOkxFgwDQjNw3/xAx/1pbVuRQSxwGedxKtJ0zACICvFekN1ywGl
vPralJeTa/PIffx1DHXEktMKZ0FGIhJimjpq152dQwL6yymhlOe4U66nFHUqfM5qVitvKc+nAQ64
MqrYiJ7qzCY/tz+jVEUHZCBJBdGrQF682ihmM5Lj718g0ulrRMYVVhtGJ1nzKViGDtnly+KWPa33
hl/v62kTYAFbIFSA0dOExdoLpxmK2tiBYcl7XHVGKElNeFzc97YfmZ4f9gmcdsYf15hRClEwKTy6
KaQuvYSrFndfROpYGZKOLO8dEltL2RhjnndYFLLG+tv+3hBVXgY1ZX+GfRzl4ETwv/PXZBqhFEuB
wZSsdkquzryYyoBh0n0UH1lZBjcgGmwxHNFqzT1Op3GfKoLON/81RCkG0vZCv4w2pRdNii2cL1aa
hHuLDLfrn7/cJkNuADHsdErwhLsmHdijvuwHQ+44ydXnyctVfTn4e0WqvX7Le7rKoWYW+qtp7SqT
Cx75wkbcxSu9OXqtu3lt1/MqraHD9jK9B1u4b8Oeq0jncLDmDEr4I4oeyzk9rKh8hO5rhQrylc0z
/hFOlCv9l2IMQVWY12UlZ0sI3pvPVDBP89iaepFheWvwE+5LhODAPkouHpnFFi9xWTPtOdDJI503
BXLUV81aNKnGzxZ+Tj6QryMM9NcEkncNk7h1LyQyaAi2+fTSSsehGBL891ancyJ8ytIEuyiDSUvR
Z3w8BqYiXcsm8iQCdN84WiwcHAS0ULVmZ+cN3kdQTr9nD4F2gL4H4DNjgls9OaX+ye4Z0t588DRB
47Bl5RgSYj1NXmftLOEQbX2dSqfO+qGwnm3VtqZJzPb4iJDz0AKWyOy7AVP4dku5Xpy8Y0ONipbw
fK0MbmUCBjWp+9KU182xh5p6+UioALXAl5nMPaZRZGIGVut2t+VXi1W948Gavq/Z3hWG1QVaWgMP
Ub0+42UID9ErOLNEd0LHGqcS2jKCKsBRM4wiYASdrdRxxg0nHQLn90ByIfWGarvcHTBvNTUyuxwj
9Sim9loXQZMPZPmhr1F7vaydVA3X34/CpWeQEs1qi3TrA4bLaPqsZI9EH0FeSOXHl3UA1rHdREeK
Iu9kg/BUrrV/cabL+8SX3cwLJHldbikrSF7jZ7Hanng5VhGEkIdkfgjewYMXlw2gzh03ODJTLubR
1Qby3IYeKpXLOJjhPTFxNprfqCpC0kWa3nn6agXr5oCkqvYz00Y82F1QP50o0pWBhpx0xYlghJvi
8D4MZNXbmCHaU4hmZBWftDGQE6ILFKuW2q/HGRuhBH4qhzb38uAMhVhdTFng1B7lc5DNdk0CctcS
umnKxAnruY+utb3zvFN9PL4ssORi1mCp+Rl5bIsYtRslxmjAQjr4etUi116efAaFk7TjhZ02/deK
yweZBShAhKni9/7NEL56Doo0SzfhZMRpUCMzjB5Qv1MbLlcjPFVpP47XupihvcEqM8Fumq2YDMQb
MHH1YeBhQLny55vLWGil6qftNO+pJM5SDeZ+2k2uN3FRdXcGZ4wL9XlOOR9+NvQU1RUMMp3OSycI
1wxVQDC/aCWJFz44dradzZh+sJgRUwtj3nMmWz7W2iNIDZo5tff4g//a8t5eNFvdUOSsoQgbnH8D
LqHQfhpEr4zPlZAJQCKWs3xiPc3ujVBd9zln83wrLlMHrDGcSYb5+BlzEpY9AL0iAYsTBb9GWUsD
isQkcYTO1QMEfU05R5ZsUy+8bsZ7oV4iv8V108XIyT95fcjDMXlu40SCaOBK7TFOKd7q2ONAzwBN
uanE64y/1Ruve+jjt1dsK9s2oLBxfxnOfKPs4lFCqWGzQg78BlRU3iqTIIro2k0JNJBEURe8qd8B
ziUdDXEcIkysdbvK1ai4NLU10ET8lb8dXoarCHEKVk4kctiAlyhkTDMFphmOR2vT38Wusj/3qhvo
lMBUe+nBwwNIGnEzqT71mZMopmk+Jpi0jh0I7sD3ZcRZ0307Agbs2soku+7jhzT7/YWiKci3rm87
8eJ2cYcntuvo/qEGHhUPZ3POnc5kc25/qow7sYZbv2alvPWJVAZvDN6Oju3Q1B+TDwr6q7NoSrUn
hL31LgMJ0hFvy+ATQA9m7vOyukiyajMsYOFUJxRMiPKzVqM06uFTP1plk2mCC0M6sWkQSbxhOSQK
bMMSSlPmdcRQrdNWgZ/L20zqw667CRa1+pCu/LYRdGC/KXTzwNAUD3ane9mtw/gGW3z4KPeSxGMv
5QDuN5Cqa6epPOi7PT0i1ElVTvZHFo4nIFjKkYimC4tgJZi/fuxezDDqGV7D1veV2QozFg1NRsQE
vyzciaB7qvPTvpSt8dwTC7EcS6S1Ly5puOJuCP1nLcHPNU0uynEplx9s7gZ6/WDgaVqVCoda1u0B
QbBFxjFoMeiKjayR0li2x6ZTDZwbxr17c3WgyRjTJneMckeMb30x0gC60B7LUiImZNZaLfc53gMg
bQDobkkEa2Zv0Z60i9EohIyGJnw9AYQ8g8pmCTeh29sE+5Ht9iz9eUjoDJ+c7nRwMNkZY1v0cdFj
a0zbfWa0kVOiHsA3MxClORvAeVmtcGH8d4VpMb21XcJCM9kGAWC3+oyMrCeq+XkOOXdfEE2QdT0P
Gp2gDUvHu/p3HoTjnX0AV4emAIwC8+fkdtFDAx5BnbokIF6KEtmNsHufTH4tlGtDf27Nx1x2cFP5
cPZx8tEnCPwZ2SFOMOuyZ0dMbjjaQbE4olwQNl6SvHsvzVQLVSAtQdwB9igsV1qqKq2QBE21Y0Za
g8Qd9wwMCzxmI0JV7SMxiEmyl94Elxe7pYy6Xy2WZ+DaTqtEtwXPfq99EIa7S0cuf+0J6eX8kbaa
9vYcxapet1UkCImB3DRrZh+CXYCN8chKRRPQBnrTRK11mXMrbP7rf8/OQEFHfN2fUD8SMKmeXpds
R/+fLFqm5v3Jz7nYbOl37dB9k08GHoUDwS+hLivqiHa/aoIp/MNaSJP4evhSiMCXida49eQm3z39
HSRUhaVA/V9xdUJjYFYYvBdWZ4Om758dDoX7fykuGsMB2i2uFcPp1IfCV8idhcRQAOzkKTPPpY5v
5YuZq/30M/klATtmQxCHcIRGAeN7ZoRHSzxbOmmODqGmulkUMEoTJJhMjXl6zr/24uucvZ2ipr+S
KSbJQMFqf1GOOOukAtFwMj00/cou2ayIbmJgRd5oknNIIwHX1FVVY/Nm58ush23jR0YU6kU/GCAH
J5RhbnXTINdg4W7bq8IJCaNrXEuM3ehPBBk2jeNiuMTpN49Bom2ZfqCCer18kCKwZtEbD5aMruQS
pFe7J+mEHc9eG4pw6tZjE7rGBbolJsNRTg7Av5knMWVu1x6zMyfyZVL9mOQ2m503P6jQLdG+HIdg
QyOUhjLd9Uvu+GIHLPl+Bey6n0frZXVergdVzQo9QPkw0/9L8kHydx9D3Ytg1JlYTFntr7Z5H7tR
QaeD3lpoHiQkA8i78CFVep0LuGiabxpNhKic4xdlCsdlidV3x3ZHiYC/vC9O0uegGqGuBIOP0jfh
vkW/N15h9Co3BoBE7iO98W4GmFa1tlXipP7RA8jPCg/2BsaLMgP6l7g6YBCeMrWVk+c74W1Kne0r
MPqU558fEk5Aqx2pJq3ITaojJymJcUXg6VkWw9b3XqTZOuq8LGY3Jo/w/7YK4pRXJsKLjTnH2Kz+
kd3zdrbjPxow6uQX9Ld2hUH9Wat9FxnbZ9zAda2fx3VRbmNJm25Q+dljZ6xdVRATMUoi6j37V2L4
Ccur3ujs5zo9ZPgWO8J6syoG+0XsneyrhUfqbVVsc252vbhisKjptdH9HyAAb4qaVTiRRhY7/94D
kJglPLs7qoZ9wNsc2YZjxEZsJaX2qi9ozmVho4Lst9SEMWzsBxgdr5Ub760puGGIeteCPSix47yr
cQOhKbRfeHRTm3uwR1n5L1Rrg+Puh1SKO+9KK7COtZ47OoI6aY61UET25832aZA391vTSU/4BcAs
Ccs73KZJ1tkSkhw5TBq51OTLR9apLe0s2OKXz71NNnst1MtuZaCDAtVsxJBKB9HiAJS/xWpgHiu3
r7yzZTuIRjEmaPU2hOKDTaauUiUgaVtZoyhmBc3+pTVDcoicubA4WC4ELLLp+Co5lSrudH8hPJxY
YLwOq64wHawVjGcBfr1oEs/PJEhZe+rtKQzDsW7eWhyUHD/7Fyids+je72FWzV8wA4xuszedCEly
4l2BM04GSKhDmgWp0+zCm2e2MmoTov4uPsI+6T5uvgnTgqfAYYgSPwh+Rx2isb1Es+TH9oJXag/y
agSY9F8td491GLc0vjuKn30UTEZQwWcnMX1tRpZ9q8O+Y+1xqs4aA4xBJxxD85+bomgjsvPcxLzz
BMxwtRHaMoWXQS4ECYxnwhzJ0E3toBd3thGCqS8GeH3FwQ9zbdZK/Ol1GQ/92NDxo4S0fV8CaJNS
ESEQNJscRfa8k8nCyn0YHPct0nyVXO3aLIVhiUgv3V9z+H4Gdn280sGYlv34uVdVWPNNPoM0iBg6
CDRxr3KRNz6tt718zCRwo1QBWz2I2uEXs0qVnn6lBpFz1wAqrIcImaO7MZDYxuv61NECJQdJqGql
KZubm3fblgFSzEf4BzzBS+imbdxIxS8v2AUAER7uQAgPMPTAagXHae53R+sLhEdmvj80mujNWmqm
by1bdTTdyrr9V5TluVrTTlghzbyGk5KStoLbBvtnV+2NiKpF+oQ42c9eRbmxvgioGfJElvCy3Plw
al/qHcN/IiNNW5ton4c5UQIyscV5NGqG+vQMPiQaTp8harAYqUPMC9pzPwTqClwGkAz/pO26QuU1
O4t/wVUUYopVD6zRiEzBANJEGz+hMFKltdZKzPepWZ1in7jqFUKZXtpmZ/nDaS0YYU1afDxfkCSS
7hdi43/aTR74wyS6Q9kBmxiS5Y+zANpz8mPEWEZs2t5kxeoGUCI84m1/1+w8dbKYHvDuHyT3MVUN
lxjecalMfGd3CjBd8bFQA81dk5AHZ4R13utfwTm1yQN7ASrgrkODih/S8Uxp1rsrz/45JzlZQ0I3
spEW36dTrxaQ03H/F2q4lBPMj10iHj+zVOgCM9L0h0sQi/MjQX9rufxEic6ik3hT5wTwlQZ0zynV
3JdUU1sTxrqZWs/2zJpYDQXJMloFJdo6DAi9ku4oaJ5Pk17RPtq0BPORU+NRyIN7sIn/sV/87oBU
0xJfJLFlodUWuqiZqdyOUFwiw8zYjQkJilVMhgNYJAA1dvOcV2kl7U3LQbVCUfJ06yhLfyJyHCWg
Ynr6zsFzVzK8/jo52CMqD4Ipz4snwBc8Bk17uuTaAx8MIITqaOCoAJkVn89MidKT6SEOITYByYUM
rjmOSnUAuENAoS291crrhiii2b87veKG0idbPCtFiFeZrydaDNnSx+KejcQTDA6hMlr2VLObPCY7
wl1b7SJU57lptJhdfqy+j+abHbCWvRIi0vmAvKBcpVBRMC3YLpsCL3wuD8ofKuSjbA7j3QdclxRE
ItxYWoZCcDF0j3DPYdS9n4OJs74kqan1x/U5EKacaZutKOS6LnVc4ZI3Cpll36tYnZLDhLBV7Zo4
Lf/EMrCXux8+ozHZfDzakFwnoKzkIOBCLmtsQIcphtRczpynck2GE3U0+dp/9Eod0/+nI1he0lst
qMCUkDU3tdBqMDDplaUrLQmUNHuzl1fklTmm5zREo1Ct3ygfYIeShTIYLZiEbjqclFYyl7kLkX70
ouH0WRWFRGqSS9kcbCjuAipOl5IvFBzYUCHfrtStMwJZRm5xYHgDfevWvQqAysYGk0A87IHp3kyn
dxRBQmh/Y0jpKd2HCVkayxEqNDRQ/wxQJFsntJF24NzlZAUezbEQ9wqaJO5YPUkLBqRXIJ5bQ3kd
80BZ+avZcDpPOzeRyqw84uvyeYGPX7QWQrEOQeqDNiIaOtOwe5DdCG46zMWE0mP8iZJZYmCvXhfc
uNAkzwKvbGnJvrm9Pj7w4LKs1jpVvgeB6KUVOohjjPUd2RgucyCFPXGJPPczmUsVnFHEofby7OZY
Vwe2qSTy7XzHaWPL+3K9TbRP3IqZP5n/kK0qysPPBbmD/pWTHSIkrfs9mSBPt3xRkbKr2oTFRm91
uM/QDHPyztY2MEV+hLoxzPvhIEsvjamjj/pcyv4n7Fz7XTn9J/1egjeTE3IjwJkWrSQ/vuEFGPap
57ZzVaftZpA9MHwmA1SFupWbJVn9tXo5HJkcsPbVhr8+yYXIcE0tEySeuz3Nbb/S/wvYgPA46O4m
Z77orJoZF5HIEO4iZ3dZvAG9QVT+3vQgOz8XPPtBlDHL3/sFIPwBxqKPOgKLV5Pf427FvPtw/CLN
L3VVuLifUwTWIIHWF8tBskbXQAv0lbZGG8vHQ5bUzGZDCIIM4x3OVmT26urzr+QArhbTrwJkbrsq
g71PSLjSM3q/aRozz+2vkuGnorKnTTaXCM4mIv+oi29lUotICWvrxzOTCdEBXmCYDxGrwUVwmUBV
y4gF/K++WYCplFbvwoZKIg0GbD+DNfBnNVcEW++/MsrwYJxR8WO1hdIK5QHHE9MxQnJGIOGov+WF
oVkFiub3Shr1djpwrhCk+jWGT2pMJPpz59RiDvqQSaZwdw1izzzoZbjYZKuD/FzH+lRLCyTXxKf3
90aPPzG3Kq5Z+KgtnYu/nZFwHHl4W5JoaeDRIIef8LJozKQ0yrnkGsN46zsNpiSghF4R38tUDbzq
JEZx3Leoa2x34fr6oNTaGDzeBFWTWq9G19FzNSPzyQIgQL5zhuRh2wpJPyaE77LnaucU+iVJVd4o
h2iY8AioxYbzDSTJ06/8a/MK72q4V835YEuZbuAOAjBRbRCObcrQjl0cwe4IHi9rfkVF7Mj0jbXb
VFcReRuAg4qnPU9rH0IxzbPVbkoc29Yqt+hqJ40ug2qdBGId2GZmnFXgse/wZunOdaK+CvR5rKHp
tdWp4z45XSacEhw4fvywq/csHjJNoS715/ACK+WoFqtPXjXHEgmJSAxOc1ONe0AX4kRtZFKjTE0X
3jnV2tAWU5gNPH803tBc1xbCEQzpbfzFgQzuyMeaYUd+If1R52HH/GoEzGevXDGnUXjHDyrjcO+3
lkD6jxA0ixM2V0F0mhKj/X9ch5CAm6x5xM1uSg/HsVUtvPvJyIWA1oGD6Cpx0DYP7/ujt3Kikzuh
a1BAgCrpjRmFKpIhKHxbjvUH1g5sdM5H3CeLE3j+r90eFz84ZJaSSSbA9LP5K69M5YfhlF2WurQj
o2xvcEAtjlZa9MWlmP0FdXHkbl36p/R95QPrQmTj9Mjvt8j4UP1qQBtPcTLJG+Is8Vf07NJsunWx
eYZm5QbN18MkIZEdYgGIsqUfbKLyVm8cWzySmkiwAKJZYFDq8paWB9SQhVvQ0opoItm5iEANTiXl
shlpMMq++et90dCInBRX+eMMW1VBvv+7ZHVZ14r4yELwRGNY7+NM/lE9aMEO5ZAL162OAhhtSRVx
lJdY2A+d5OeLAYp1rCF7J+7fBMd+gZEcltJsu11KsRgBZvflwfz8KHv3NabbQuGjpD00dqnDF6vk
4hkdP4gzkRvXoVlV4fiAeLHvGwixB9uSjwCzxgylXbYKim2X6tMldhK8fnUcAPjvDrPwSaybSIEm
qe+aWRm2TpdBM5X5Y+hOGF3ciIXhr6kq4uuYQlXuyyA0+cW1BOEaJebXm723mIPv4VNXSDf1Fxag
REc6g9ydEbzNQJ76RBCQxqTtZ2+GIIi8pbVTTtc8O7irKgPhDfcC75CVKnWo7YJ8sLXTGa5aD9Bs
HjrPOxfjnrEXk1w6fB4yjb3XwfPCtmqiKS+2nvPdw6K7Xvpvw4W1ngS+GKj3VF6aHEeTP6G+8Zti
d/3Q6P7t79qyaXGCCJchBgnkctz6+NauyC9WHAvA4S+eHT4ZsCQmxADV10bMJM+axV/+k1+u8GYh
opuFHADHDXj+lFGTsm+sw8KwPeyLfgV8H3fpXhSNsbQ+Nd4F/c5wL3hejPjlbZkFENYIOrSeZq6/
osVUDFEEGId200MGC8jioMWIxMUMvEo6QA96YlGJcH41HjLt2C8IfD0FJ9ny1tQhExDISgpRAMBO
gCGMxYLdsDIyHlXDtr8hG5oQ8bsmwmG6wBIZLrupFSqRNfcaqfHQcjrRy9/pGugWJi6cSYmHLO2j
sDd9VOUqY2Q/KJ17yKFVOEiKuZOtGrqg6wzKC3wYhq4B1reDryb8CqiBRYgTox1yhFrBujyHMVHW
oMwg7RHSw2CTSFM5yQia0YZEFT6LJdbzcveOYpemp/7w2gmuF1Zbdp3i2nK3H7Eb3aUmAr43DwXb
J0QieMHuKU4uUzHR8bKGUhU2w+Tc5wYMbD+Tb/jMYlCSXjSJVH9yCxh9HvW7sQZomwxCE4xmU60f
3cb1N039aL2hRJtPDLZPz7oECxta3deTERRxsedURfmuo+N6/sKHoOQE3+f18Q0P5sBn2JvuG7xo
D7bz6Aa/155/aw4xs8NJUNdN+wwiJILZaC4N21R9XXXJTOtvEPxYSZOy1LQghbwHuU6SdrGH8DLd
2zImyUo8cuhcHpaYmFIYw1ynJtQE+8ReDX3nAJiclb9A/3oRhvMtqD756BJJpsRNfxbDA+XFkzjK
W5pw0kkq+uEpWimqthZsRjrNXnRYpRT6lyRkI5a5vnlrid67Z/Skr2D3QrSBFKsOPOAJVeVnJdCB
HONp2Om6kqGZbbLtLKwR6C9QJ1MH1lzGoTQFTvMoCHUnef/vadbCbAF/cyddrN+rw70t2zuO8bna
geDGuNdiHWFIg21/8Eze2yBTOLhpWEVhR7Jy0QZVsYRKon3M6hNhEKZSgDrN+JHfLNKvcT65lTnl
QQESNIBOrx5i4EqJKURWTRVLSqOdpXpTB5q70dF6ZoUT0UC3GJcTJrlULMh8BIjJHc4Y+5/VR9J0
XOttM6B9BOjnNYIn1S3eF0QOcJ3DY0nxJZxUped/c5EXPWVqGZI4XIjtATthMLwSC22EWxwVdu9Z
Es1A5xPKt0o3QKkgr6r4V8k4N9w7YEK99H3IbiJVFQ6+Xm9XuJBR3b8LLU8VyFbsK80yEmOswhSE
lCi2/IVFNAPwXiFSsa6pCRvAmy2pjAfF7jacmOmDhSub6Sxb28dfvydAiMQ2zZ17rm4pygDZTmni
U7Rl6z9QtFm8EmDNC4Pi+afQ5UIo5DG90KYnqxRZaAFNX1VDz0J6473xtpVzRg01zgzbvTLfRGIN
M6mQo2fML2ga34LerLkd2fWnbuJCR2TgH8EUZ79R44gkhgoKxDg1pWMeN5n/ae2KcziGpspimber
fmTB6MCLiTlrYKHjx0p+knombYZzH21I3H3BUTq5b2SnhQbMMTLzR2xwGTnamzxw/ordge0wMQn5
eSMTkmwqd9CbOUJItgKCfsjXJ2eCPl/XjqZ8uCw/T3YG9zjlK/DQEXGsgokVNaOQJgHoFthRM+Mw
w2whsleAUbGpDWCj5BbzGjk1P1aydvO86ic1MImns6kyV1iKWA+WDuK471fmapU0pM9LotD9/jMz
9PaCqKmHSFEr0rlzzjcv25+LKvyeRZYLswYB6zr4u9GArB3bVXFOu1CsOCN4aMCao1TTeru76yO3
xUXPf7WvtTRP97f88TR0gohlSwQPH0TkQt9qjUWYhRKSx5cYwEC/iuyvgyByq6KdzSV1hV3IMj/D
S9eTNrNVSDefh5+feIDj74VczFQyqU164Cg7xCzlbSpjzUvfdLhhRU587oDuYHUgE+KRSRpk/sp7
tGfHNbV5NEg3s5X8K+L/iu9OoIXs2fZKrskQC8x8I7mbccVAMzZvUFA0Wwhu02rCuIiGhczVKA+u
tz6dxjGa69BDcdQq6xwnVl8r/LN3xdsnUjivGS0Y23Ds+chFBwVugiSqrXo2Klz1MS7151JvYz6g
icmqdiNhK9fVpoUSsngekDmijNsZzFgW0l7dGrWE9hXC/ERNP2YDUfl9lih0f6tT8+zEYq72VbQs
Ulx6yInjigD2Iw1EHMp0W01zAFCWkQD/BgEbBSjcCiev5fBi670y88qWaUQYQs0QUGReohAHuIjb
MO0vOH64wkKgD2uc5bdyQRCAlyO59tvIfQpuOl0VmMMtkf4H3+8Zl/sC13NyPOPzEn3nG4I8518m
XagZNH0tS/n36Ezgoxy5/CWtahYIQ5LvXPiFiKJJT0CAFwGH0luUC6tKDxyGtej6egGEinwjLBEX
4+2qM7lvMIDOKxe1/lstoKiOVqp43vvridFG+uG7eLP+0nl+iAjyDAQPQjwJQVHgXYIFrF5eOcmg
T0XiX0OIqky7QC+KO2A/mKFfgmaCembtyGoaEUBxuMwjCs9zgDh5A9uKJPN1/n1HEIrUWOEjbga8
L40krBEDZ4jLczUYWBogUAEBj2h8sd6WvK29MUGygFS4wmT8taVwqZCLHRZ+kd9t/HgJ78gRU5yk
xkXWomq7+9TI8kKg5nvKVBjOsG330lmf7YxRgpLrCgm+32oRCuOTX4zWZOXlCD0Cr5u/nBQHJKU2
1vbwu83Om4yXkctND2q1nMBTS9JCVLDY/YWjzIYtb/7QndqzW6De12TfWFsrgIAuU2ragYGPN1f6
MnoQbmJ++Aw39DU5ic1sEfsXHpoQ/UKFIoJo9zZ/acgH/FdygRkiSjxkZ2rfwt/SijIFbqzFcIhz
nrBYwbqTUwlheKNgKWxZUp7FqWCqZmp7kqzhC3I1QIOfLA8vwZNvP8q8Ousx5kQ0SwawEpo//M7V
7GDcd5WfHwniGEBKxKP+Ch/ioZLqbMt4MUXATHMl3fMDAOepHnstPr3DdbalvXJGaHyY09OFPiI3
7SxMI70Qv21x3aHdOSc/yYvmW21xU2RlH/PWNwkvuM491BaLRUacGElANCoCcAxsjxt9PuhqXeVN
vJDkcxiluQU4j5x7+XjQ65xGCyQjU1qlHMmTkwPH4b6knU6+sLpg+VyZpFte7M7VUmEdGvstwCQD
Q7sMB7ObE/Gm+0+NYOFjB5VqTXRx5wo8HcJqvHUqXWt3I7TMz53x6ckz96PHz7arvjU6+mun7Ca5
oaeqCkSvrICWRXNvh8SCM46UM0dOd5yFXIg0MywL5Mz+YRbkdzvuXtlCYnl9zvoFkyK09G5pmEdj
7jMfQVXocYARJwRNIdv2YBBo7NefAKTAom7G6CAj2cbMgEPcNLKn0xRYVg1dGtlkXuRyqCqlWwat
esZofPkPT81ZqW7rACRtZXhfgEdUKw15a8bqmJygqCpD+0yHfLge+N9Kc2B0W1FEspxc4jSfpP2n
QKf7xaGyBcVbNeXKkPFM8a7lOb7s4LDcRGN8Q1zhx12nndKaQxNjjdjIBxrjUF/QJuwh5OvL+KsC
8tNsM94bdabfTwpHz58MdAVddFkqOYcgYGJpjOKoO2a2WGt2u28xtgMPqgxNtfyTCXYKdxSV+x2Z
z5cRUzsYk4h2oR0ZD5a+9ARaWX2/rDKIHed6Vvu2HexyOXqD2WRxKO8LtlEHHQkkyOwIdXGbeWyZ
hRE7xNcndRbhtMPbGB9Ah9h9SUL5Xr9KtXeYKmUzePX0FHw82js1G/CpnmYMu8OSyLMuYmuMpTEP
PX6dXlNU/AN2CcawGOOiK6vzL0vLnffPj5AvaHqHJMqU6Sn6+e/KudUvAh1f3bA2SdoUbeFeVC0O
JGKLcmFWW5busj+FsQiQbkXmVZEG2LCbmTAmP7DWlwwBbh5U5SMR9Z29itA5Fzd948Hwou8NJU7r
IUmdwon5ntQA7Td2F9fQGKvgrbCMUkNGMELbBBQ0dN6LV+4j4qN8OGNxPrHB+3ApVmAZqz1EP5fM
1xLf9eVYQUv7hzT+gQ/LBK63fhX4qfYTUIuhaEk9Wi3zutsqg263JVA3pYl9+8ZqpjIFTZsUV/3m
EKyN4hvhb+mO92E0BPziAncqWzKU4qYU/mcZHMeswHZXPbjXNAEq33OAFNqbrjMPRNnRuYfjgIvb
s4Z8jrsTL1wq1A2lck5G5lJTO9OxVsPO+RiVgOg6OXnrCh8eMTlK9lIhlMsFHu+Vy1WZgQGOWNAQ
31PzrN0jxgL1pDMDx+G9c1bAejm86X41cNsFtvl/AIF/dicbT4OOUS2BjJuWHN+tiHus/0QWYn+g
ebXdDuuMr9/kYdf7XstKue3CdAUL4ZX/wMBJq3vZvCyKHBHI0I5lSbkpeIO3eLmVu34s++3X5lbd
DszYpSjS5pCnsN4knhvRlXUyF10aBQ8HzP7C14p9mfep7CFhoGY4DTuwAYxoyW4UbNdgCMcaQMVU
X+RwTKLDcrEMh5GC34nOnH0X+ZD9hHRCvrskkoqaBg/GUmRifXk37Na0vRr/7SPquci7SUvu2b1x
wm9ydwanNVqWppu9puwidMRaDE4ukIupi/e/daXFx06M8TZ/1UO+xaRYJDq4YCjYqbeccwHtkj4X
0mOjq50zLacS54LQF0+SKvukv+ye/uYFITSLcr6HfYk6oGq57dz7CvRQdpu0PB+tjndvyfCzJaF9
qo0y2GbC3ZgHt/Ad1B2amEHYTSQcsMxwZfm7wbmC7CmCx0PaOIFbLPKCZpCnfozabw6TftRgVdAv
9B0PmiOUXuVQI4oEsxdUPsHwKlk7z4+yumF4MaG8ISkflkZ3a4IG5kPGytUNjGfFjMV4rdI+S4H7
5S+3MNfJbfVsn5cZQonEF7j7JBd1eZYGBAx2Ed2wDxP1eOiBLAC08IgPKOn/Qx03jTMXi1n46Nfn
pvxLY/TeHXalS7IjsSgXK1WDuT2H52f6AjUsIy8xlNtUcNdIpNs7sJdmiJ41C7rR4zdsmde7q6qD
VW2tNjFpg2b/ICrrO8uLMw0hZ3wtzoUGyuTqZbYYjyTE/Ns+iK+WQQ4h5X0ktj3YOU6A8rxLjgZO
m563bCXy2WaR6U2UwixekxPyYX6KaDTzJm1v0gMYM1zz0yXOMJaslJvtelNP6OKY1TMBeOuJ/GEN
Sq/hIORJlb2+GAE6gWVIWqIGUYpd2bbEGVLb4IbZiK4tyvUqU7uO/9vxIVG9QYLcRgvRFMr1yGgA
m0CKugkFkLigB+YAAP5RpyBWBL0x8q8vSg6wSRT5i9kMH6Xr7/pSufysM0opwEYFMiuaD/k3j8HO
9YlOHt+0upXMOTKVmNX8Dh9Eph8FD/wj/GXAYvOuMAbh7QAwO9XEQ1VEzPLp5ARnOXcJX+c/nCMJ
lBtcjptrj3nrM+TBQTYCLfkhz43lOctS43lzs1rKirgh5eV2ncVhSvx9V7RMVPQstIAE/MNyZdjD
5xBKA9jb4IuY1VLKfygy0zt3HWytFGmJBqDiPsvEkT7v5KFRbdQq88Vwjyfr6tYv6O4MJWu44BLq
OLDofQDcBrYgchgKdWCSzZ1MyOlIPtcIjvaTj4Aa15JTmftPh2E31K6970sLvXDjl2B6pmuQmwZQ
OdPnGywyTXM3d0Roz5+OrF7Z0yhLVF02wUq6JaLV6yJ6SIZkeg2i8w2pSOlvAD8ag/MclNt/Ii7O
uKnM/8DGkhfNuWuvlZ8FwobTP+7sh4vJVCiJKWVu/JsmrXzqMt63Eo5lhFkpmKQCp/y1j0Ngvnqb
Qpp+YcWgycrb/k5VqClQ3Z8s32gOyT/zU+2c1KQyNZbNftJ2NGV0CjM9ApJ07hCjVs98dd2cVBK+
KrlkD2xOUjhCVwLgIpOIYm3ypfiJ7NEIhrk3xmZeWCNDj+16c8w1TiI1Juzm1aXhjmzh/hjX2gdy
+K2BSeuXCDrlMZGKCTF+0PAg3JDp8UBjRWWe2HAHgKJmRPGwObKtu1ZEE6rwW6E3vcQV4V0dPwAh
GBx0WBiU7aJKw6/VeM1Y40CVL7C2AsAncnBasXF/nkbzNpP2TJJg9xvQztHI4DFzB7Sl8VcSMXVq
qYr4zU1JMGCuiMaXWcA0BCDsvhXoMYTjH+sMdwhz6LWJY5rXYIwwbRoWH/Cv1cvRok5UjPG7LOvT
tnsYyCEG20+ieq5F6OAvb9BJ/HEMip2/zXNjkUrtnVKrXTUSXD35NNhQwVUx4kQyPUWx+LsGKVKl
+PZ2DoSbIxb0x2xwAcVOBaImwqLohqeZCWqo1zEvUPSMLS/oApLLkNg97J9clt8BVQm+edR8VKPU
BoBRTiwBXsw10GrGYDyaa6sXVWxkgegkDgyCQl5O555/2gJSP3lKuUiFII5LWBNWuSyzXc2BtEGa
wTX7MIo6aZPRHth5cUw2Clsw/AxAJBUbUXnWY+MqiP3FM1D6TlCLPPke1/TvNYeLEay5jv73O4QP
7RAh1gJkrn3NIXZk8hB3RXprutRUHk3AxegD5uaQOZVR58j0FnuHy6nmvsqhee1isTjJ9rMrSpSV
XQ47+t5uSHYa3Ap3fc6XYJbCrmNvhV7AXPOSZq1Fm+MlebQcatWUMXcZ8olXAZUdjdx4wI8DU12K
wokYMTYdzssQqe3TV9txKJpmo8jSMPoUyJ73YYfZcgXYeIcCdff6aXz1SjkJaFkT80XuGx8YtTQr
3ijNkvJOcysClq/UbqknOKY0DAvGMvjD6u+D+VeQ8Vl4huHo6w2Bg4jLoH8u3WetMfxqQaINhhbm
kaw/TdPxGuFTnCnh7tqxzw/fv5bfbSp4xIaNYIUhfaJB42n12pWqdEzypYYnBzalJLPSPoY/J9C9
IK+JEg19qMYi1uYKGNnAKBj1QDha/NtgeWMy7WDa1Ny68iVfivuWDG9bpLGakuenfZ+zT3I3/i7A
4xQVNZx+6Aog5McMfENuUjvA8gDJQ5H8EIc+TR9iChEdOXHHm5rZ4FX/C6bKtWQJ3zbWalpkQmxU
xwj8odNE9fVYL8kVUZs3bDDCH8p6Mr0xG9wCSfy5sOOx0NPQF19PfTSJPTy7vRCeB6yimYz9xpBD
tWX245EGHG4QFVXkXZVc8D8yF3Qpy9M3dgdWgxti3BwcOsbwclVnVHjHIet53Kj1YoUc4KmO+xs1
czE+ic+gmBvAJT+XANiSegKbUhhd2fxXZEN1JtEoRN6QEM3Js0aSUEe2ztJrAJUyfIQG4HkkW5DF
iS6CmH00YUjluL93d2etX7FwU3ZYTfInalqZYy+ALI0g+H6OK0qwH3xwkQMTZ1vEsr42ohRvKn5B
+DX3+79vrTBArD5GWnMMbYZmfSdR3nFgctwRU0kun7345kbaKSmr/qe77ek919AnZOMsuy/ypIXO
PMqmAGtMaxTWlUR2g6GlLL1AmWZ1e4yxuCay1BmoeMDXBgocbZe3cmy0FRui3t/SOgrsPpeWM7MQ
hZoo7Cga9CQGCMw4DujU8/5CDDueHcPk4hhauHbsTPymRRxJynZTFRxcfoMK9/aycmKWYvOjQUcm
5nmAqd8fLa6e/kJ0eY4BPZ2x1LSnSb/ts5bmQ6JrLdAsCEoQrkLeWp95Kb++c5grO/RBv3Pc+08K
zhbHtskls6o/ls3SA/ytmAV+SLBsO+tR93OWqjD5QbyZl4eJw4e+CucrNbhlay1Ynq7cFc8BgVdw
ez/go5k74hR1SolGCz6YQTlPU893BuSZv0l2jmJW/GNI9CXwnx6hpZJhaXa4wG2mmQi9Gf5kEUNk
z5LT87jeQVUmfTsCfO6FlgBcYRSxh8QA5KgzqbcFt+wF9TPLJSaCm6XizAmSbdiByLyC7AmMe/3i
fNroVB1nUCrLxP7UzgDwEeaXqn796C/z2aTaB1yrHWrkhQ7WrUUH+gsUImaV6tYay8i+oYzhLsx/
t5EA3r+9/AAdvQ0q5t0ZR+grhKrG1BJY98mgamYghoYMU3wrDg1K9wEXXWY0Aa4IJgezhuHDFN40
FLbZrZc3667SaeWRwQPTDWwdKPsGb+Cadm6IiE8dYUUmHjvQ7mNHr44Ylj2hLkR75JzxWCBNNu3O
RqA8caivgPs/ic9973rJa2JVvGwm4i4PH3oYcsQl976dwC1NkqgE4+E75Wi7vvdiCdqNThcdRkhr
f9wGebH3rcg31lnhWzPSa425JYFqwTxzKdJIezwWHcgHJa4LxfEyoA73Ece4NbxSjLTzcatZ2Shq
BUWGMqHrOlyOiaKihueZHK/5aV82Ppp1P3zSygSwDwL1jDceV86wJmclCrOHBxDdrNmxGXfdh9nN
TofO2NS4afdJQA8270NZyfuRFedaHkFZTL+MYJGA1PzQ2mZUU3WN5Ia6UAvfcGVpmkDwLBb8DAmz
kMjQfoow6LGUbchrWstlcOdzapdBY0Akel8yT+oy8Ej9cyUchvdX6Kfc6dzWchUvn5LjvYCU+kxK
yxT764aWT45JmeCamZ8gBTucDmwvTcAZUmSXkK8DIT+cUdoel4ZmkkcS2Bg3c/Sc48YHNvrU6RHy
fTqqHIE0lHP/pwmqrVQZeEaVIWRJEtRJ0sutGLF03x5sWHV+REcPldKljP6kLKnY0jr0lsfj9S4X
JtOgUHmlw8WEnmAAu1jqWM13N8C1/rTbZqs6+nTqDGPmXWY6u5jZqa7OI7ZV2dNGJG9xV6U+PjTA
IuDd+cHy4u85dvnjYX8HioCXcZ7prbSPcAweRYl4xBrRwcT1mm83+FZeHiXIrJdf8gz3Fc1KSCD2
iimhhrqieIKAcz2z0y/rJp0Kx5sYlF46srPtKY5o3Esvs3Gl/LxV5sKXfB90FPQR8cTOy9S1lHjm
dlkMnSKoZL8J/872p/YauqiCufE2suzBfjL+nuKRziHuWIno0wPFfNro43D4zMQH4kWvJDI+9LvG
ngpOWU8SWH/9oM286hrIse6bD8KYFpKzGvFXn7pEzqsrsQEDfDrWsHDoCJGkWnsGrAEcfxScYU6g
fmRWpSOlyeT3plSTemY5u22Xd/hnQZNJI3mQHG48evK9sxxnR1He+uSGAOWCciCkhMtonxr/H77a
iCmFca+p5JXCbLp7OA1uyPGGpgy1cly7VTKTUJWq9b9K73njLbyK8ntsphS/WHVf2B48xK+8TOh8
D3/vGShOxqLY32cICwuwra2+tBzeZpqPP7W7Fr4N2J2NZdZ3BSEQqGLLQ4IcJrCulBoTo+IOpDAC
cEhuAp8bk+iyUOjzrpi/F6BU5HZHoXeSLfDdzJsLlldEItW2rRiQSDOIEBS3r0SYsHdLo2CI4exS
Jnwt8lvKX36XO64RAImIUIim/uP5UIIGkbLFJuBYMe98j0F4cQrUNlfqNyTfghicv6GfxIRQiPEC
3344FYgAJ1fp8CCng+gEpRnwLeCODrNx7jeNgdz8DIA+bJgBcXxFw1dYqvweCex1Eig3gJ/7UllX
HpLlUZBRmYJcY7rByqEhPBxmPM1SLjLOXLyApwXeS3j0moHCN7CjDTIo+xVKw+HhdtKsqYqrNnla
RNK/KvM05DsYFm6DGQthaavcjmbemPW/q6PHA5BMvCbnf7f5s59md9v8aMt6hLalip9PMiUcXgMZ
c4Cc8tDjygTZKQceckELq3rZDGKqhe5CbkoEThpX3jdzHrOr+Lmt7QYor1mlcA08of5NxgW4o08i
kicOLnTlbObJ4ITsfkap6dakkVYP+rjdOSPcNXU/Vtjbb7dMhBe6S2gQ0J+l5H01kvyw0a7vBYS3
hxBPLTf4ocecJVDggr9J0AXRySmTjn0TBMR/c3o/1EukUm2GfdmYCNui/F4Hc4GAq5KwZdXMIiMB
jC1m/tgg3s6v0ossfosi54w7wtgZ68tYYjNFKVlzUphmpkc/p5tJKR2WHGpllOyUoFfG0ipMEUrh
Oj0fezPXmkeeF2gIDh0nwkOMW70E1/o2Dg+EolkilyhuieXUlnMOgYhN/IkXgn1kNJndgRUddBuK
2YtfqW98afwtG2KVk43vy+x8i3UgIuWqsIejKqTtbAWqiNjrEZxQFEtdDan4dLAEgH3zMkfgmqfH
+Giz897XBtw3DP0DaBepCQDO/yZwAeJzsHB9NgxMMCyLg8284Cn99MsBZb242gXSrW/cnC3xkIdN
QCwBGFPTRcIzeXn+aa9qLqRAH7SMJOMKOocHPhu9VXMFz0PgvuifEprAM3wId1IKe5lGuuZjpRsX
i0blu8gXsUrL8C0Zn0KoSViuKGFD93It78zq+HJ4Oes/JRj58aKXrma7MLLg8PcbvQblkpkWaQKV
In+8YuCXu56mfPPL4L0ugedaLHk1ZJWoN+lqkB9cdekm+8ZVGzbgyGaDd4FLHamzZQp3wCuYDfrn
wrce0f8kdWQr5yixOn4E/T2P28M5j3VaFG8OHlw85fP1u2wMwrczIVmJ1HJqCxuXGeJBNSuS/MdY
A1cmiF7Wsby82Jpoms7ABkKYIQDxe4efpBdPmtFG1yWgAypSIU7ipFzvifI6T7kJT6E6CWcadi98
qmDo1dMH2H0qraNZ6MfDRoF8VdVVTWo0TNL9Or2FYSy22d1SXzApKjZy22//AcO1iYYZnugGqN/w
bVfPsDWp/lSIqe9wgEn8mGsXlfwxbNYXsX9WU59W1g6mhUr+ezT40Fd0xheiGqcGw81g0UY4V67y
Khvu75xmU+oiliyeq+TRPAt6VjyNhMUTwLRi9nBealUxZMDO/LfzYXxRtSPz4d62Gc2FuBbggUer
DffI77lYhsIJoDmxz3opjjovDg6+ZeYDPMBb/4J0Ordrncg+JfwQLDo3U9oIxgLrwwn2HvR+kiN8
7yobfsn76hTqonmihmocBTJMcEKbAOxxiJH/vrZ7hHV8tBycaa+1YsmaHxJorqbXLYwyY8/bK579
eYHeBrg/sJBf7dtJZtfHd1zgUieQNSCTiQtXYaxjYqt5r7uqY1+pRWaQhDGWMZZ48frB9QfCSPJe
/z+/A+ubnjyupPGzFazJwkKodIThMHBnA4tl7cuJSfJlA7hltkoZyPRpKD2L291WsdoYkHXXuQ1s
vXm3QBRgp+qcpGu7CO8dBwZPL1XXz7STh2LEicIJxNmSxkEK46CDoj4hE1ztM4AsLSg//bEMnpG+
uEgA3ujCwV4y9EVORFZVPo0hxwYJ9sFmUWKZWL3QtNEKA0t8kj/kzLL/34Wg/iZ2AJPm7IPtieu3
DAo5L9u0dOgq6dndRHq2RaOwS1FQUUzNg6CkDVKPoxqn+vDOy4soJ0ABBA6iaZWyr3ZudyXnoZd+
kKFA2aIVQS0z5ahqG5HOO2g00Ji77IGHf8pxA45cHz5g1Vrs0XUepzJp5enydBcatXGNJWDumV4i
RLnpkJs6u1EQDHCDoTH0xlc5v69Hw4bsKVuz6+cNplIzHuyPq6PmGrZ82GKT14kDl5g3HtXhhmuF
yynKQwHqzdxwv15/nj+dRJ0oXqY2bqD9kIEO8GUZXaq7M6sCqXTQzoiKK+OPazGackK/cFV9Tyy2
rHo+a6wFDGf5RGxrq+xq2ptIrk117o+wnnmKpFYXzc7zJXGMhhi3dycm0MVill4LMfJNWmSSaowG
zF9JqDVX5ZEGZVue9C1WEeWAPPE4t6sXav3AEtqXcucYNUoxRRicsU+eA1RCu/PC6Te/RktX1PmC
KhTjSQWWRgf0dyDorX3FmVc0l3mEfVt1YzYG2lqwVaaYzgPGTct83t2OqX63hEljzWAAyXD/sXlO
luAG1EBSzhfkxpbaF5GVeTWz2GQD9eBNeW9FCVVZvEi1O1UaPW/5priuxOeSrNuRelbww2EriZIY
8lvquHGSoijly0Mhmm4Ug87PdL4Enj2hqQCmfrSdj4HqiOybOaLj9AMHKeMDzbg8l7Gq/WUFXRIH
2q5qdsLgQyrkx4h1TJU5/BQYHJNzSoWZpTc+7khq0EtirYZaI/GcOcHQ8FYpQOnovFIFJFEyYUjJ
KNbD9fonuNguJC/V/lnlVPNGq7EgkC3QA0I+1Hi44yo6XPHdIgPa98ftp8UK50CqRpvbjEfyYQu6
XBTRIPxrcRyePPbzpmgHJRdhRFJ6nySFVC5mCXxp9hC8s7q7iF8TlQl5ERKTcjD0LL5ryu53MIws
FA3FLWFjUwBdeYitVtZdekzUSGwYoWI+wT1/ynP8elVxHHHzBjItRjdrAgbKq4Y5HX1HSwdDGBv3
vbydM34wMn7ruJSa4IjR+nAVBz/jrqJsnevQb/wsj3cSe8cefDFQzxLl0zo8tz8ZkgVTtMCdvg2U
fm2ykK+JjQZLFJwMB39+2ttKd4nVuyOh/kraO9DmcxWiv4RLeysY+gL3mnWFPwqNMqYGtFCO7A8r
djlZs9OslTHQLEsxwQalVgHz0aDIAWUVs0zJ46J9wxZBQyXEYr81tI4OJUrHTsHJjELdRkbC9++5
7jcejMF3w4szpfs0KkXtpVmskt3XjL2SUqZgHZBgOALVY9prLmn+1gDDzdgfDjYTzfkslNzU5o4r
qSCdq77dXn4pVBo1EDrePsC7Fa+8TGN8kAIMjtJPHygxP6L2dmfmBXM+gB42xjXPDZseBrB3pV+L
T48dN7X6ONqer/SmQrSQrKCxpnmsg7WTZoK1R4Xxi4Fyj+dImwLXA5vxqCkEkm2yDSDv9bl2CSSj
ryZr7/fWj6gB4R+8crXNfIg+pE0uv013gNJCckjJ/v8cDAmczjfljP5e3BqkblpRmUltdR8zsSWX
4ZffXbY4cY+ZHzNXz4AzY70KNbNZxr/74XX+BeZShrMtvwmlO+LpMnitr2wPy8p98Fyd3N/g6CPg
8KjBgvrCBgIA+hIqOBDvusWMD23sxVCn82RpkoS08VA8KSQke2i5FSBJXa4k87+uoAxIY5O0VblU
BxBCLztM5zilbFQY169aj2THCShgOY4ZpAw2767aXNIqGamdKiwI93cRQLmQ+57/6UCiAsO/lv/e
0tFWsFz0bjfUDaiMwtPm3zAa2tO7mMhHBIm3Rl3JJSffk/qlOEoCjP5R9qbLDxPUEWQJs8cbhA4q
M6vSPbxEaZedA+G6iln4u4d5Qq0H23nRWVxQaOdtWZ5hQJiO1vsIXZpNC+gxdC/bCataFqOPDrr/
6xXrTwN1h3ZlnieQVFmkwOJXgS+tQLXmZG05/ZGujhePn+F5ZUqOGN5DM9aUwRmW9MSU+C6EzI3D
JmeUgGUMZ99gfkANKK69AKf+3m/qOGgidjoeF50m+ttaXMewgPCwBX/7H/J4qsN7HDJNiRr6JLOX
7xk/rtI+qPJ8BPPX74w7u2vzjgzD5DpzmGioegBkUfMz6ozVcfrt4QvmTMLRjO7QJdxLiljF2rsx
7clC564ZoZWNSSBV320BAE34d9yGfltUcnno7dN2XrlczoEXw1+9iDmaskDs98OssInLZG36KDba
N2hnmeGCMfHmsOB2KshsEGSJT1JAQJOPc4VcrRLX/N8+4uiTYR1weq78a0J07vKI4qTcAsdfFeYv
+4F/izHsgrDtY9CyiqhYwDYTAtj+jTKtsAZxRUa0SicA++a4a0JrAkMyX90aeTaaJv52+xH+QmkP
Awnd4HJs/H2VFxwyujS5jSJW6ds/pmcyYIErpcBA+E59A2odonENjdVma9eaOlEmZyX5XIR37+ox
xsbq3j+PWtshuxKL0Gjsu1qWdr1WiaTlmk1cu302iYWzbHvwOXcjzXuFetw6lLlr+aO7puvFpMiM
ia+ie5aYCll6iOXxABa6Ef12T384Vg8OHKms1vtISPMBIGM/XjRroAMFObk152jGeTK7/vQhGGH9
4d9VDb9/vV4G1XeqGqQmh+LjN+hA+8PiJaf6VlQAVgQE+sEq7apwBV/daqdkXyuB1cdHjR1XIXru
3e9XBwJvSBm64opRIeXpKB97yWR9ew1in02gS0Z2rJAAmqgRmVwpOAOOCVJVJNHNBaR11C8bn5bB
HWX7KOfRy7iR/PVn83zgyM5N0sxONME2G4s9gkyAeHkOxDyCunh5DWmjc34Xh9qgG6Gxdztx3Imk
8Gp7P+YTOdiGPXEsRuCRWT0x4Ju65HOm2oJi8Lm2RMSke0GZ0dqCm85arpaxAGVEbOBS/Xge8rYK
Jen76fWWeWFu44jphYdIfPWm4PTJFJuRWm7rakT27vT7qnNsjPrK+l4mtXTUKZX8oWyziOGb9RIf
x4Sj2K2CIMlSfWmdu+cxUZXovpzBqci3FB9CvWrJofe1mFCPPIboFan4Bk7Zz/bg71nYGVBRfpmG
GkaMQyD3BwmgfGOUUYvRopKJQV7DIses+ac6JkHAC7KvfFQ4ujwKeteG8gVjGkXR3Yf2s6DOTAM9
Le7mkq3ec7vS3V4ntOJ9YupE7A3qjITvj9JiDa2oXkfsbnr+tqEVStc61CEi9wRL5vGEEKxUoG7K
7mJgwX5H32hK/oNMqiEbB0zQG0W31zp4i1qwJmlzGIHFAeZ1BVoV/ZtFR4znXLuEMEckBC71pRQI
RJEcpXOLmE/QqPKcpsI1FkV78Wp7qLTky/9lqgE/eot0Hv+35njI5HW5yHuJik6vdGRtBr+yQM0o
dQcfJd83h6rjVeo+iWJGrzZnZjSnHqGugAFmB4iHYfn5GJ1KwbLusgLNkJsTRL2U5PB57UD/Un/N
1SlM9VNxct+Kwy7dqtCvpSGGsfUAV/SoXrG28pBbfoegpK07RiWQ1GHLDOn+yj+hX9kOfgYy1IxO
CwUQ+TjfMXXJECnkONm9ZdNK0tiQFyD+OH/xx/wkRJ7sI+Ffui/5yxDBJyS0ZaaUwKfRlT+HAujP
4M8GyYijt4FzSPbWCr6ty9rgxzh0dL3UxQXQu7VfPeAB/gc3qTpO4k5WWQuFBN/JW/0agm8KEyJE
FRidNBINAlNkp7iT1v6V10u1SiwauW8SJv8wlXuE7yq06vbSKvyTtwYJwFTdM1kMZNIyOcCkkb9Y
7VoBw3Ca1ClP5YEs7ABkLiFulH8yPn8M1EHipPfy5tkwGIvZUi53q9pTuQIaIkMiZc1piRRNYILp
ZH58eBoLDsclA0UkbOvy9no7ID2oEd6xfeAyvHOjGVGlqfibjcu/6fVNnq0qmfbazxdfQk1r9CDx
RnHhBVbHoi7EbArhZd2B4F2Vnj0AEywegJKlNSFZP1x0k6qTfLr6xTpa9hHsULRWij/797kEjHgY
Ea6e2DXE1VL7TpAfWyMZ0oZRoQmnJNOxBVMj2CW6Zt8mYiC8WZDdZfsDrTHUmew+68WdGj/cXc7z
Cy+jgy/QWR+Pnoa1hOTbW9bVq422pGQ4Ut74gXByYQH1TQJRsgg7fOhuqrYZYuD4LDM17ue83Ivf
zBrtY3Rtu3JiaPlrUzeEpmXW9tawi9xIdWRW7vMb2erm8Ul7bA2Kva1WBvcCEs1OQkR1/jGAWxgC
ud63pUzQ8f1CqjibZeYGwGDpiljTBq1bAUhheYoc9wAu7EzhleIFgfChgZ5FsWYYi5P40YKq7emm
Mei1Lr6pJJ9pjNI98yib9u4C7lkV4etkMUkjmAmXJTwtvHdf4sInpjo6ls5c4gL9BkyNCqNSDqLY
+Mqbkuijhal9IkuvFCssxYQfhp59MZKkAvvV+o5uW9bR8NScK+cROWc7Fzx0/ZQtBPtYA15NG6u8
OJpTvLeyv8DLVUPtX3+bPJ2RvwPTGZ7/92lyrWFV6ulCTCjwIcCmOdE8Fd7/KTm2W5Vv2Uw1d7D1
0wpT1DBGFkOxGrDtKN3oGXox0H9Gtm5ZBX0LkvVGtNng1kYPZWDWW5uI4nJH976wHQvOOrGZnTY3
tNJ74/Z729QkFWAigOnaAo5X+e7DrUC7nAFJjoy3W10yHMZ5Y2/RXvOExjZQv9+m2AqKCq9IcDgr
6DhLrmW2JuAjgq2kDpCYG3jom/Yyhf+ojVArQTzxVj6GJc9YxzBIM4CNr3FzKc+l81Ul5LIX2Muc
UC1yp17K6TXWGmzqzwkahjuiMoue53vH2eL1QXEqyMDNwN6IB79n5BEb5il6osLoZPlR+A/qrbhN
oJgE5HOVt75SnbBbfIEWNMBI6Y5EpN7IR6cgFadYl423++NQZ0/aVKyBdQMbkmPb1IBC14C+NNdh
TdG1hKC2Ju3JF2h8FW5kUSflAPQAXl0se4wOKRpNFFdugT6bPC7tYnLBW8PZ5iQM1JKg1h+nvXd3
iOgpsYZCb5jrI1KmQ8T+f6OR1NPLyrackaDq+c5aGUC5KniQFNK7QfyxvzwnU9xMFvJcTTe6SvlY
VGlyv3LhFyhucEYdmWaqgpAjtQXn18V7TR+AiC41hL3P5zjGTq27PFb8TSVqhzSwM56nGe15oXW3
SMyzwp4qmdd368kRYE1htaXgMzSrxkUAmrWRnsLLom2ltoKm6fcKpsZM/cjFL434bTrYKhVlAY0l
/JgcRgGBW87v+/NHIJgIPChCH4cdy3DggLUy1MM8DuIQcB6gcJ0j0VclEDuRpCjj/gFxZqk9PT9z
qj7GlFGvYrU8LgyD00QekdEEn8jNNUqZpUWDSh2aizr6PmeN/Q4+vnqBMcmMAKh4JSqbWaqbakRZ
WntMgYkNsI0pnorJPU+kHue+E/x4d6orAbPeqG+jVORmhSwYqM/NpSMK9JokBF6qyjitOL7GCgWo
7JBEWQC0JdGPo8T7JoIj280jK1zLdQTKChadRuzyTGwpW2+h9n6omAkcqOxootzWgDrmsCBwZShD
BYgNqOw1cuWvrpZX+OXwFuGHgw2Dp3eaxTaRQmkZi0BSQu1tbdEm9/yFTKyqAXZAg/tElL2jheN+
ot5cw2WF09KuXnz6x1bALafmyaVJZvbkxsn8iAD4OjuWJDQadtaHSOtkYqSyJaLgQVwGGXB7a3QN
MhuU09O//jgUu2J9PICmcu8n714hTHirhigCh8mtsnatruCIEDwGeo0rjSkUjlr752aPRljdd9QB
vIf7WZKXzt1vaFDztpyvx+agY0Qk6yepHDJ2Fnn2ByadMhxkCgENZWtce+jddjZoErTGnUPkfVCB
JkLTlF2hbyH3CCpDZEdH7vecR3IC81JSbMyjA9vPApT4eAM1GGO5ZI1+F0pXcmVHFvl3qeavxEci
Ut8K2TgXc/fKOskiXiAybASOOtC/nUuVYmlul3ALsjCh9ibYBJ/HiKLuLaXH9BUQ0jhcQqyuufCO
dyk6P6J2skS7KAJeEwT253D/JiCEjqMRMibDDec/ejOKifg75PN4RnSu9eiI5C++EweTu5h8li6a
XDhiz+VQC+a3w0dhXEFcmxtBUryJ/2rTRgqDlHJHJ8hJN60JuzMBzE1D8VtskMaQb/ZJj0DSXAN0
O39Xn1g2je2jUjotVVNWnepofTaQhphXtFiOR40wSccGuNc9eMhFy5FgCygTIDwjIqFYIlvS1x/A
ORfv4pQX46NIS/k1uH15kBv/IGldcEiU1UDOxtNW3EfZBptAcDXK7PzQWtQzIBvoK1vbaSmz6P2s
z7efFSVx1i+cQxIAQlppn5HVuBX3e3EIgGyS/V9elhmB1pMzEvLF2CbN/nafgZ1XoZ9c3UqRSU7X
ek2CpITBIettyXUC8paA0dsEo6QSac3lmQwAWUjB4HqIX5LnyCuyENL82CVtOTqrHaCoVLjXodjX
4El4+OybQMgB4xb9vFsVhZca60ZAZneEEw7S1ISZFKiE15klVaVx6gN2uqod4qIqwOFChp2vgxej
zUlWePV4aNNoHezRIKQVpPId1ExLHIXSPet0pCL3B5UbX4MIeLsRMY4xVDEb+q8XM1zwbb7qDozt
vn8DtQ9ydHGFShHWW0QF4F4D3SB1z6J4xfkMoj2dJPyaKqnD1hob+mi6l0FxHHvq6BhAPWD5npqK
pYS4LvIS25oR3kK+vwOa9En5h9aUPBpPX+zeS8qyruWK9kNfPT6qHk0vVje3WWH17lK+l69jN/H6
7EvZRECp8OXOylQ7mNOkbdfab5UJZa1Rim7fSpSvMaUDSPzn7t8GmpArlgnRVTGV3xNGrqj9ZjbH
ISNBmWJYPPcnXdeQmwZj4UohKbw0JMZwKLNIQzkqEPqTQnqmidP6j8lRrsoqhqyMUs6PetY4oASr
mDHoEYCzAsTc9kiXtMPTMPVX9XkJE0jUkBqVjH1d1m9qTQIj5kwllIold9UhP4wnCf42XCVahqfo
CcY2lLJkzNlTNVwFJgjGN4UPE2b/Mol7uMdY1prZDYWrNrKnwo9QUCkGzgVy8IPwXxa9AnsDjPPz
J4t1IKPxrDWDGY3oE21ytrfsaO0NCYRUihmORZvcc/bmM972n0Mb7wg0OaAHxC9UsHQK+sFMmcTa
IOm9ncLz0IhP1KTM86MO9Wvzx9Elyud68K27/gIvWTw0srF5lar6pg3RljIGmGbfGPkkcmyChjBs
fMEssfboehe7u2ky3XFyIzy8fV2CEJb3YfxEz/G0ka2TqArmr+/to/uo1pRhSz5KRPqUMxBixSew
k6ANeMM7ehWCbwTuNhePmRKSAZ+TKW62D1qyk5k+FHASC8Gnu27O5D2IYp3TI0Lp4WQ5rux8S4M6
nQZLxalGT3yWfyEPlHoS96Sjvc1+JZVgyxfBiLEj/tlMb5yfk+fgRjc+il7R+QfskZfdCCBJCIl+
cEAerpglXLs/O07JPzR0KwDjwly4TgpZbWjmLJ1EoO0TMoOo6LZLFxo9ruxCic8LvYy0sH449M+7
ikiDE/uqEfHHMU4bawUQOfSLCbETcga/l3soi7edJZJbs17NUtp67zbKl7SUkGH+U05ht9ZX+oJF
ZsrP3Z3UOkFYFu83oFq7OaAeEneyQSUdltxUFeKIwomgTe6jFmFYueZXD+NtRYHsr5BY8xR7zuw8
OulcB/ZHVICP0bVE7gX+9QlfS67aR4RGsMjzf4M2gYsGXSoK0DSFS/E3VLzDOmepqR7ophImplZr
dVPHBGbBfsRnRTXzXxfQ1jiXmdLr7CMCi8G/wOiFrUREclgu+2x5HVU+R5iqyalUrVb54jvGfyWV
+6BaoiByzB87qlfUmPJOY08f3PjmmNIvM/4kZrRXwtWcgBDD6SiXTPTfZO7/jpNvLh9+0+sKbwhy
WPDveeBIWOdLi0pIjcN41UJ9st0xmuIQtuzCmQZpgCmbsP8tWYlOcdbACtTF7crH+JPFdK4b/6DA
y9nPZbBeo4g0UweY35CLRPBvFEsTgKCWKtPorZJqutAn+i8pQ+xP0s/RpjPmrFc7VVWAoUn6BBRE
WGnIivBa61GeN49iaW1QsHqi+WF8EUpgDxYo8Lqbwrpq6jMBJVKHSb1K9gFRUAlXCjzk8kLywWJ4
7rero9iBB+HTPCBq2bLj/Lu7mtCpPVAlw7RHzZSSiDi3N1xzuxdbZGpPmYt1Pxg+JqKL7jV7L2Rf
mkF3x422xSx+m4y2CgXEnI8YAnQVL2b9hlWoJuH4w2nz8mQ1KCePBsEai7JlxY+A9Gp++Y5wO2KC
WxjvyKiYYyWTCscaXx7yQB3YSgI5n12ZyiM5GwvFh1jxvB70tjdUglqiSHvfzDRxBSIp/3rms7UH
sHhsKuTb4CCX4tRgKnrCnDD9849Xl0rL6EZRCyqq5enC4oPMPxkYRzUSXwYT6QkhqjgOi0tztQ8T
wImUBcE7BFTFmiJtx68t4Mp842nusFc31bGCfMPKlFFoZBvUnsJVCaX4Js/kRXngGfbc1bqEK0J4
CMIq632V4yHWZzSXD3oE+hI1gBQALQGeZwG21PcpTtFU4qSBS3EhCnY3dpjbmM3h+FjJqAwdJpxI
beDPS6yRHUsWxupQEzuAVlvV00qrOmmiXBZr+usCHVtPV/3jkPHKPACQd6gKevFHQKCXlyJUzekK
6678ytfcAzmkmJFXmJS5ovAefCJtm31ee0MDcTmPiWaoOtpF89nTkKWQWSILBlEi9xOk67gwMVjR
AjKVcjEjlg/jBvOzpbqMKHvZ9GOTLMswcVK1KBBuQytf323ROSV5DOUrxPo8GUHS0GGxUnmE/cgm
FxNdN4HFiU/GMh43etjgzl5xBGuyYmEoh4bXWwZF5N0pxnXOIfxzGzCyZO0SKiXz0I19WuLnX5Ii
0bBIdH/mjtQRpMUY3FdlL74GyqKZDINbC4t4V4KaJGsdyVAgt2aZ/RwB4pyKUFepAFeoRuNgmklx
MX5QK6fgYauKI3PocVj1dWoaeG7LQypsb3dn+Mq3GEz8XZIqNvenN53Djd34/cZYrAMtV7y15MPX
0nRMWsr8pBrJZ01qQNk3oWo25e8Ox9pb71Rtccd0GFR1DcUlHq60OgY5XDLT3ZwGXQd4fIBhojOc
g5dVbrxxl0VcdmPSHMySG0x4u19xNRgBkG0hAFZ0KLMli7D0S8WOK0RfdQcOafl/MH3q1tea7KkM
vFDw4kIuwSPWiyEFAjKKEcwArjJndnVnbJpk7thkC49sqmrIDhwqGUY0EPS7zcPwbpwCHjqxcvoZ
tWwtSonnMs+oMRjcxE+4wZ2+qtxbwttuEVVjYETLuHBLpNMN+rtdI+vX37QYPrYQNtu2G6MMZ6eJ
9AHSO5m9hpV1FGUDghBRKkvk3iFl50XYxF5URvJ216DZmTTVeDIaCD93Hv4CaxVS74YNiKjHK2gc
GJ4ozp7EVBaR+eJpyArgCGKiccLk/Jswj8f0tc0Iay17RSfcKNBSjZX9/YMIIzWV85yf9s2sfp/G
T1BBB/0CcM/M3dOTnMelvAu9PO7O/RpK5D4pxOYC3/CNYPj575p7ThmOCRzAavP5U3W6md9cBV1S
gHl8v7POvo5EKoZfk/34lF5JiFhBd3muDicO93rok84n4xPC23i+Hfle3k1HQ79ri4G+QGM0XlbZ
QNjjq+zsoq1n7YQJYqqsYexRAO6AjGjcHBERZ0Evwx0sFWJxIssc09Xn1Zt+EE6Ps1M4nx4Yn6Xh
dXzHssPMgSDPgQ9b2t5gvdVn7tptJSnLlTBvStzzFbOVfoIX/2EmXkTPRkuFCdFK9ASIFmXdzNHh
JFiXCmlxzynyN7QjTTSfLiDTroB4GS2hKdMh8nzzEXCP8DZSbOqLNuxwH4WYO/aX+2T9p0sT7qs+
Q/yeHeVePRDnsmIttJuSq/iqw24nw7hN/UPT/JR/smdg+RsfhDjHtgiOOLaXxF8rYn8H7LsenEic
gxFfq3ypixqwtn7LWvP/P39WQ8y8cq6VpJKy+f5L1Z9MOsLMBM3C6NpPo3fFDML3t2btpCZSLAWs
XUXsNin0sA9wNUC/BRsYUyma540tTPDupWoi94E/0PaYaNSqJeahIQ7TbozR7tSr0PB7/e5Ucv7T
pkSQQFGS/YEriwyo+PhDkGewwG5u6LIskRNE+HjUzmr4YL+O9DejQ67PmUqes1dCwdzmHMzBSRSK
sWivJfNoy5aZcKbjXwsLQm4wkdPgHMSLUlt3ubNlogM/z27ew2vOcByi3HCmcYZh5bBdK7Bdpymg
4BYrHWL6UeEe6cLe5d0IRjHinHKbKnj4H56kt2Klm3uSGvamCcejKOVZZps+zkBSwyDbYduD/+hf
/woSBLc1WG0yGMtPn4Gk3Pcw2reAf0VHLiQ2XVrUF6BkolkYni9jwGpii8s6UBCltIwzYbk94eMc
aAcL7pl8ESF/Qo+lpscCdadvu4FC8H6/qEhSLdnz7D6O33Tf/T9Qm+rxu7vTtmcUwYgisGcy8Pzv
/wuu1l/zQOxswNFUKcaYdPhBTCZI/27003JCWbTTnFR8aln+exjN6a3SjeW5FWCT9wjEXpLkEAQj
XZMHSRQYRl1/sNlI98eP4C9PuswYu3P4k0XJOxgb0k7ywmk2UJPxlOnA1a4a2UShkp5vJB76ozVD
FSUGftSUnspuPyAWWgOJp67OhyqOk7Fgm11EPnP2w3tRJHJ1ORATXqdGBGiL3zwSQZLLeiYoRQzi
2VXVsSzHPH3F8Gz4avLY2xM4e6shk6dLO0mkUJzwQjtlbm47ftY/n3/4zHrvT7YUF8qvTXSo/+Xv
R3MD7nqAuQzt4HQ/NdRrMNAusoGhvG8ng6JOnApBcAXq1mn6XC3l5QspB0MoGEPe8kn91mkKqpFj
DXl2tAX2z+KgfUV7x9/zbiToE3yLgKq+oLZlFZu6hUi7ntNTB9Yr+lNXc6bYS1SNQ85TB1REqk8Y
RXuq41fwJxN8YYNwaXtYq2FvwCMCJA9NDpV6qaGm+k9fEVVIidBelP9VxBuvwg+x0rDDaHQXZdYc
luNWpRB9TDHF9MWcpNANoUPGnlGhsWZk32Eh9CEqAsZsG3/oO35t88Tj/KY98D6cDsfX2DbAMwjD
Rj2r0bAUMYll+9aUGJ1mA8D6ZZuKuF6rT1nYKDoY9pfuG3T24hVJO0rD3zR6kszrSZY0tWiSe2dP
XNHr5Tchv3LIqZHnqUvDtwoRGpto1W1A0mdyobeLWYwfzIzMkYN62ocnW7oQAVpG+NP4QZbraLjy
4+mPDqEngwMuFCMz3ahjY4P5Es70XsedxCYUG5KMS3wf55eJKulLpDGBN0CNDGeXC2qEaCcdT35I
GeBHrDi+wECvBinu6xSjKK6dykqLCQwEmQGO+EZBMtl7o14dJDVLqRQNDyyaspvKXKXdnloaVhYr
KCA/xDTkUMj+/qzn/YsmHAvrP19PZTsRvBvwMJoWGg6EJ0e0N57R82OTEIcHtPa4Fn6Aa9yz2fyD
YDh7tstmpB0SJ/KZ3Iwxcxt6y1J+JiiEtK5lcV6savPNjc/dfaz8YV2tNZTRLnopvXLZGhag2pI0
ctDRCTv8KJYbguQDKuvJ1akBaGWWCxCJFlPLtXCfDROKIl23R64nyHAVi9K68HoXNtFE+XXeSiMe
ovzod0yMSPvwksc1aLNe2TJR2mGf8Gm2YXcz9KJeyE+e1buyFrqcesBgiVLX1uOZtJQDj85sfQSo
LSFpdQpB09ACbVTNXT8NQ/QHWYhTixOj92VG2RZOMPDmqFuHiEjQoTsMIBuBGuc/7NFNiUUZSv1e
KsoJKXM+GM1CWNSdJxPoUwn6Yb1OC/2pLQQbtKfRuWgykK2btcATEn4i+B2pi+IIgLwC3UREBsDw
hxvRBEgH5L76Bha+VgHH630Eb5iCZepJV9abf5TuW7o8XFYqoWUKpgj+mi/jacKzgoiSoDNBVDdD
/FCqZuOBImcIm8blKE4L79vYNCsUhUDvvh7NHe+qYJoXb05/CY5hw44FOA61tBIkfMHUqtojcOen
8X6/jMRqRrFJF6UL0t+SES/0dGCIRdGXT2y0ErTj4qTaSGNEck0EwSucNXakL7rcsR2E1I6lLOg6
ElkWQujtM/ZYKYQru5UBhA9qjbowBdUEl8gSyaeMHqwb5VsrGtHzmYQBbjJbefOBnFztJGx9IVeF
e8kc+iOytdv1tLfH8LMwXseVdBYVjR2A4Dp02mhnnpYYYcSP0KnPe/Cf4U4pZ9pPiubyrEoKeRbW
+IgpiJsriKS7PNa2BKUQqPaYQzjzfGy5/yyNc+BK3erranONmeROKd8Gg6TzekjnL7vshvcc7RKk
SW4OhUvA1llcjGfH3zEfx8WmNNhQhFzSv3sHSRFTEUDMExt1UgkesRLA+F583bvUha4LMZyrG2kj
2x3ps1EvdAe8SOTC5JRD/Uw2Q6AvZDjX1qLVlBD/lVj8sk8Ux5vBjLkMDV+LXr8UM1Hif7F/fAPf
XNlvmgDuKx+A8wy72TPs/geao/CtLrH7jPyLBT3kNib2cjNKXwJZVmqcvCgLUpyjnPSczLS5RucG
Dm+81co1H3hEHa2Nu7s6ipH5jmop0MCa4mZnrYtVJLQGSmrBQpAuqNF+1zUIMx2Jyl6V+sml+dqC
GPhgTOl6qN9Qh8Qq1jiZwJP8gI1fjlhBnjpMbhBSjRdR82tY8i+/7tlHyx1GCq18eS7zbZV8ef5K
qn492CGFuL8CHeFvbeVIyulwlhmPDaqmrVv0OupBAgid++9GvKG93sDo7grFSVPfneQeJqivMV6g
TBzhJrl8NGGMd1GU7d0jjjdIjuj6vZjjiXWdbSZpgLzSIP9ISN+zop+pbfvHMn9Djq6MPykZzJPR
Nh3SHwFXYhmtReBlKVL4qSjC39lKifyj+RRYORxfISg27NqK3uaLWLVy1aCHiBsaCKwaqvvVoNjv
nCEVekt2HoQ7ZGPS/2aXBULY0m/W5I6uTujcV51+iOO6C0dXcIHGM90QaAJ7MpuN88rHu+iqWUl6
ab2a8bdfmRSQivyPE7DmnN+4SP5Vi4I9wK21qYlWX45v2XrTQ4WPwRGEBgmZb29SNAe848wh6uSD
RCNTWP/x9wW7x8x7Yaf4ENmtttIBNoRj96ZCOOONvtm6fSHZGgczjnwcMQdWV/n2MMwTVL45HeYA
/YMgoIdP9clbRaB6hoyGAd6F+0ZM3KWDVuNCfmlXKuc8Ahy+RxvOGWIBz2bKwh2tEF6EAVE3Q7cl
K22gHmRkJYxMl2o6z1abhQOU9iIONk2uMEypC5yHkl4nIf6uJLoG+Cy3L/mpR3AH6akNJcdU3V/l
SwbRZDI5vuHmdmwpn0TmPoJAZw7mRsnmHwljsGJ0FSclTcOUMBgLBRTFf2O8XjeZPcCK8gfJf9yE
ZuM7IdDUv1R9matdodShxWzk0CHVoUPAxk4HRb2VXWwtBXlPFB9fS5aRPwa2ZB8tlIXbaRBOQ5gs
Ram3EonU6wKg8iVRJpa/lbnhJe4zUGc7pYzumyKZA+1hly0bLWDd2drTgDiaSYsA7tRpdkI/UD3R
TAClhwD5leZHCmHDx7i4x4H1TsmzdmaTLPrhdy5qkx+D4Ze/fd0bt9rEZm5JHHTaZAr6sxkD/fow
MsyweSTVi4U5tcJ0qVMxVd31zxQiOww6XweW8Lzo3XxXzDJpmOttwYpKdUW8SZ2gLIM2yJRG45n2
2081m+sjOhN1zX4g9/M4xLi6y+a28AuUiat4HPL4XLows/zgar5SxynVUpqn6gpl17FF9OF5kLzc
5yKKqnR7fLIwD6UBx8hGtZ2XEwtGtCGOtdao1HV2M+Ic6I4EgXZJ5UvPNI5sxJ8deav3415PP+CN
vbyORZahC3yaia06OFQ/HdUAfoOO+meNKwaDXYF/SiZJBPv+z795IgUnGiDmzs3MkrZccFglQMxD
cOdEf3GBiNcqbc886YmnCpssrV3Lu++c+LuwRUL6Yx1sTRqA06el7oBJLskyANZEGHYk/jemDtFa
oZO3+nGwFQzSFZExVlX7VzH0FHT4BVP2LFfnPWbx2gcCKQNEBS7/C2cBppEakaUypPx1ILiXXjRH
AkKPLZxpJ/0IYZYOLNUfVnqpoF+cpUW57ETYI482YsgA7ptuW0YBusSitf9hCprkzhJ9dLQJkLwd
rWuVtakjlvRw3cz+Z2J3smsAjX2WMo5wz2H6GoPL8l8eG+fjBOOkA8NAgcVNkgpHYcnrJaWqF+rl
P/jX+4T1/B1gBwITPcPHoVjk3ohKzVlsO40pQEcKT6YRlJIiKvGMK1j3XXPf7XdU7twyLmm914Bm
dbATXoiBqrIfvbrkUMrwsyVM8CnEEBLewNNUE+fy2G+OvxSyK1onSYgCaDqmj4NqNwNRnBKcOXFE
qtgde4KmwIYc0ULp5isCu7izPVqFfLmSaq7tcp44POEwAGTvoGEMwMGIr6RiYyJmTnD9bYvLQdeN
XH7RQVtEiFpAKL+xX6WVsfCk9KQopQ+MOMq/5n5R7sqcSXqLzT3xxqUtBSlAR8yPiJ6hTWE+002p
9CHrxpd6pT6w2KGcLDlh3M9GebZ9usUUWJJtYno5BaoKt/KcwR7Okg2m2AX6+27PEf1APK1LamNm
N5d3mFtMTE2OwndC2zd/bMhRkO+i6hUZj8PYsLjIaupDf40fv1Hx+5E5ga0yH1aoHcqXnfPfcfiv
EQU8ZBgKn/7gd5SffkntnNFB6ZZJZGlKTS8a2eYf7w18ADyNd7D47hJ3wd+iUSoCsQ3Rb/DJn1++
Lky21LdmiOyYUiPXFL7U26T1gkGrGosL9TRnBNrpbybzQ9UaMR1v/S/MbsJlnGKxS4EVaqTTiNAm
IAbCk0toTp2iKh8plqTPKLHE0pL5L4ftgAeOg8oNNZq2Td7lmhHf3vZ9cosAMxnWfJF13fcCi2xS
7UamOnQr+1T6d6lRioNklbIKpZPwUDYJlyeO7wweggYiMbCkJJB1BCsSQyyBu1LlEzjv+6GKwDRq
X0hkd7841k925gVpuyU/TSpsS5RPmiFuLqL/EoWzu7bN55taSyyjA+jiXo/2T6IEHrNRk8g9k2k/
v0bbpuj4LfAqmJOVqhJoOmHCqfEW0Fq3Dh17ADX2mjMvPdEaRa6NqsXbG9HuxrH00Riv3xvuN/3G
zzjtRSBZx/DKxO7A8EQGkWHsa6Vi16jCAyxm6k9yim0dj0KZrGdyS4w61+p3C2hhk6Gzp64+DMrr
UrAnRNEcemvBzWDDgWUqiFpqxrsLXSqufXvEN0bSiTmaLd4SufC8lVj8jJzLmiQvriPYErnd9y9i
yoF+JX4gVHPRrVJv3YbKVZvAmqSdIDqiiky0ogECZnHTJq6XacDwAcY+8ZqFKN7RvOWshdSHhD8E
h0GfoJgx58UWJPWSoNkbg8d4vTOh6gfs0zf4UMqI6bs6Qq9pY9ab+UC6DH/pM8jOzR355gBySLoU
rZUhdFrQAWbt3bY3YyL1Xjsc/0/xpK/mlvwi0FMctkm+mhYm7rcb01CqHNdXnWP7iVGZkpzZZH12
quiIwRngtRZnn0SvjdGirAN0HiXKSdUfYLlE25DyEHRd/V2hXOZrxLdNHArUihZMukPY1Wteqalc
XonjZarWxQ0HQkcUz2zFuJoKS2UisCnWFbBfrG9VtB6izzg7Pn4ENkZcDu0eon+oXEfKOpWVDN8i
TFfN9vgmAraK55HqMBGPnjZ5jzmEPrkL11fLStzb9adiy19HSJeBh4ev6Y3hs5y00D12wX+3FxZ7
1vANu5ghqiTW6ZwKelH02k/Dl0U5xCl4+mHQKk+NultQoiKxcQlB0FC2p0rtUoHnblWGSueaUJgg
+RmUEivDRlwCC6/IPmpwxjrnIbZYj11vyg/n3iHRFITDWG90glzyU33ukZGwyC60tztw6+4woVAY
6bemASdhTY2R7XZyIlpJtj0xRsaAg/es14E3TPxGPbQ+2QTkcGZCFm0ZKvUsSsiGFkaC7Xtn91yV
qQTUEDNdnwfj1QcSrgvQ4CdRIuqP+347dD7Eq1JLuC4llnX3Mq6tQ+SAfj3NfACqPnA5QL4YVDq2
UfbKvSzd4oxK9AxQI8sesrkvwuy9m5WPh37K9VbRySrchcN6coNiQR5U65MN9/NvrNlU4IpGaQya
vTBobTmDQ6BtuKKsZaNVIg/cA2IhVyFo9CRHklvUa/wmfE+e6v5ZFXiCnd6ruNs0P3Mis+MWG2nc
IjLNAzJrqJDehJWT6zmaa3/ZpsQKxiv+Rn9cFP2WBfq0RSlDGznCjAppT1TjFX96jwi8uEjaA4/7
wrIFonjGaHTVfNPOy3KaZPTUS+DkGn9N3e9SYvQ59vzW42tsE1GBqWwGAfIS+rW1DiwRiqmb8Eky
bybur8rCfLT/C19QlvigLVOPudGhXqxRzQxqj0qFyOwNlMQeT3+JgHT+Q+pM+Lw+hzqIadSt+F4/
oOtiMRcyglzORaZ6cuFelx9mOm+3c5orlVlyYaP4yWWcEn/CKRc4Cz8gteoWDK++ZcJuRKfP/uI7
XmymoiLZ4hPx7LUvfp/70nRl5hOkqLmrkHEHalz0phOrfedsw5HssQgogKG+ETLTQ3loO4HvenYu
zNTj4jciVQpkzrT/MlenLeqoZ6vmDtORxIKjy7b1+hyJhJkYAdAAi33N23X4P14STfthgXrD9PiR
0oGnnSHpLxIuU8C1n38qiJmROfqDXcelcHGoZg7Y6O/8liY5GNE9Ih6EyilDsf4XgxmX3ufZqWVz
wsj0lwtKB5P8H6ckhEDSV0WB8wtdsmMloPKCAuqcwmC00LbsZhP9V1mSOF0WqlL3ohRzKaQfAnJX
La5O7Pm/ehvuvuz6CEpZOSktdHEZZKT5wROMNztOCRaNKs7frg5coPFt/7pga3MGKORch90KI9cI
lKBRuACSFBhF8zZtxcFHLvQyRrbSRE5j3j/gnR6QOB8Tk1XkldYP2jRcIZJcsgbqZZx1hsuYRmuf
Z+OANyPBzBOGd3n/Fpk1BPcxm/2smND0jfqqkbh9Lzzcoo0zt+C7ZyrYgPj/xJmmsAeaRcuV/058
o83K5UeIiV0UdQMF7a4dilJymz+lvxyNPWunmHJr9+Z5jkvIurDf3fXd8abLnFUjUD0drvv2BSw0
tkooeJY11U4eiUOAzu/NUcZRNpk4Fc4LQZSMIxU5e6ZqT9M+AAFs62FHcgSKm5ctQoEyeiD4lLLH
GRUVVzofEhVDVq0kkw4mt5yFhF/C9R6FPj8eegtQj/e9Lo2HWyRBtOJnNfcD4ZqB1kAsA6HecC2d
/Slj2R9tXX0dPoSCujpSXY+0/NmaKoE6y4+hPfe6nloijiPUg+V/wxCiTX2D55veoVCiv9s4sbbV
6Fmptk1RjvPGX8wztgVOM6/egs8ekPTqI6PYcGleyqpdTfSn7egyK63R29vPfbOzjlNPmBjDBnWS
TIMU5u1nqwUsWz5NJWAucFcQrSAB3tsPzFctgLCz/SHtkgJEw5DogvpQeAsYTbVzFGqAjvKo7wJ7
PoUY7L3zg2IyLej13fUQ1ABtDso1sxF8tw879k+gVCgoxd4+Ael7s0pOhk5zb/yvcpFV3Ymd5H5T
LfD5yN9JQnJTXF7fCRdovEHjgt5w0S9903cDmydJDqKoVGtkhAplIQd+Z4Rkbg25Uy1RKLRqn9on
MyCGCVsAoOxkuar2zrZZV3fhDjG2ZAtDGsA0ZAV9+wCF5O+brP7QKgtOTXSQn+j4POWqsWL62wbk
ACDHwKM1vktInnkOQCML5J7rPVpUDRjxPuqc1Ylo5rhLGYHQ+xlxZFUUjCMnaOJGlFVkgptCYjVj
ZVIBwDY0fWxY92Lub9XtDVYW/oSpiugZJPA2A4KdcR9YI3eceQ2x0U+K840HDRd72Qrz8y+IWb6G
daZ0T9H2/Ce2HDYT+9tD88Uj9LFfajm/bNiohVZn7sbVKkMN2t5L393Ny5VxtsWGiP5DmyIvahiH
ugnbgGTUhIxp8rZsNbzRgEAYZ8OggoW/ngftSgFTSjS3G7imlqTY1G4++IXInQsjP4viPXBOb2k3
RavGPQb7zAOVLeHZ9cEZMloEBP6yhLXXXx5zjdVwiF+13+gQX+ctr8uRQjfU29DWf6VNUMWsSWKa
xXjyZQ8pkIpBlKu1WLXuG5TUXl110wg1+Z7FtL1F6S/oUceEs1qljsvZF1EroMiF0sVRSkIZBFaq
ewA2wXdB09Ioq6E6Kqq/INDSdMg/8X8Y1mC26j5ag+cdXHDYPtYE5ZZuhci/pcoTGJ8tLnjgzrwQ
/YG22iwfCbmWDT4D8k8nz5FQvtRyqYL8ffQMN7jgJR4XMOYxks5obNPtj62Vtxh6aM263MU5Od4R
QPup7tgtDkIUhB4Xv9dbsRdH6IQYCaDh3B8zunCDYyLJnZb0ldhm4DuKZcuIRethti+4nohxmJVI
gRvbmaAnhAL5E9HR5mRyfr7wCWLidyy4OrRxFvQ7gu6c/QetBPt98pRp6PpAci2+OcShz+40EP1K
VfHFVXtxeLG7StWhTorVc9Z0ffNwvEEx6CWQ/Hxwp1UEd1A1mw1PTia3TdxldWSemWT/XRUKgR5J
rz/bHygLueJZgM7hdm1wFZUkxPNYXx5A3NfM9iijenm8HohKZ9+/uvmW1lvHkY3DJ3C3mnmIjJD6
CRWw9ieAWyqMiAivBh1eFEpe1hX1LqFh0HEhI7q5mXGoDlMlVk1gBGRCkYflgPsGQ/978NVUsE6i
vVmFK980OKvrVCEFJOh+tSQ/lC6PGGdjnnjwzerAMVdu+P4awHBqwZF1G0wQ9p1YMn4HRcWu3iXB
mMclLiv7kfFdFf9cHLmRvSZQ4jDIu6K61TLfQqi8OlVT0bvgpcwfpCyRcf9RFfrcjsa8m6VGULIw
aHFHTCmKNLM/nlJulU62zwj+GCk3m7Puk2s1jfFL9RQR0FRU3w3dEiYJKiHikOc1djNwxnyccjif
L33sbphhtiRDmZxD6PlUZDJrezKXjrtkd4G4FI4o6nzggERL15o2h+H4jijV7GB/2GS2FA3o8Cav
SJvALOkwLZcz/ufh0ZaCES3oOkyPt12WxKJaVGUTLMqIKN5a3FlZ11jyg1QV/WIYjxXaRpdhsQhq
gL2Yhz3k8Lx5/K5KLg/YpB3WceTTLEne/FUZQ1VoGnt6G2fSEL4CLRuAT2KwDjGvx8Hj/SblOiy/
72VoJ+9ptLwPmxPxcWdPtcGuMuwJuRwUr1c1E52e4PzSu1qzjOUgVfPvxB/qukkqY/kZipbyj4wV
QrEzPHPvfHmtodxJLpY2+2wyIHDpzTksDp2GZQ3O6NlZfhJRJLNySpT5aYvYZfNcpXkQhS/3YfdK
W3vw1qju03wAMiQfr7BqOva4fTuxPIMsFGDOPgOjORWBe1VQf+HrqV7uE640ArG60z/UgoGq7m0w
xCmZ3Kxb7/FK9Eumx53DV9j4po8TgMx4+QocJ/VZdcBqbCYOlo09DHXYBaybawIguI9cOBfPeHcK
7Bf2A4QzyHrbpoK2bamZb5G6oQC8xM7xy4l6vw3/6oGd8qiEYID4epEvmh5nQQJeRSPDzi6mk3xB
f1hjH3GiRMDi/EJmjXGp+18qPugKTr2lJLIdf5hKezmag0+EtyExwTAV338OvL2vGo9zCd66Icsc
RSwNnAMKtvR9wgAnMBIwBmNn6UDOHhBGvDbuSejCUkBaExaz3rasXcA/2rbVgkHANRkeRolHyKbj
hKXnQ4goIhQEq6f2BrTrlk23YTxCmf2nV+8OOq0iZNEcyR0Bx5rVMeoGXGnz46n5+XqVkAu9gj7w
yl+RFNjD858JftlDFEW6d5o9KdSE0j80LqTIJPrf/RnrmX/lxvJN6tv+WV1VeIqxW/RY+knfpdwS
r/W1i4bF+Y+ANLuuMWfP8pNU/CpNHJyCxJskgfDA3106f3FRpnmsYy3VZ09iNaAEq4pKrZlzjKb4
K8frYxDAvqcj2K0VjqQ/9UcpG2fb+k/EjyHgQC78fCcFeopeeZpujKbfxOKQHGijTMvZCLtkaujq
HEskfa099Wnmgy/1wnk8e8OHSnUhlMZYUQoeq/Z/L1MvVPb0Z3lLkWh6mBgHUlJ4SlWXNlTId2sp
zF1tSj04DyJW5VRbwApiQ7qNn4G5yyg25Jx2d+cDk1rT3MGLRbtQX30BQJZeTzGl8MYoEl8FhWb1
lz+24M4SiY9ufaGp2JJigKHeaphvpjmB+Uv72Dks2Tq8yQ4qickTkepl5TxRLNrs9J8sgsOxzVnF
WMwmye74t9QGSxPG9GINtu1xSvYR4hwcF5hPFl4LKI0oFJAKt5NUpvF1vJK9GJpL6zS0kbSMQza+
7eRlBZKbQGzSkKwNFG75WMUOEx3ej1daLRWM+yG9UxJZxXFskXnzrQsFutc9y/Pnf02dcX5xWOiJ
MiwI5vX5qm85L+1exYTbebTHBI1jAU+vjcOsO6HTlE7la7fT8e5X3K7DJshiTOFEm+VJlQbW0oNb
UN4pqHw1TSyFTP0VegiIjlVst0sS9jBaIkkxaUun5N5N/+HUIJ3kSIzbrhPLmdbbkTKYsSHHq8fb
eaHwfHLiDYCmF7PzVU+SsyELyEbu6GKZtcbycGNcxNTFeNTAv1OCl/33/liIQLQLWOAktgWiIugd
4HMn6Dpk4QoWudeIAx4LsGQHrane/VVQ4w8gBnW7623U7/7oYSHC1BxxL/VjtKa0WnkbT/TrIXp0
y019VVYgv7MRZJHdOyzcf+9X9XctSYbFyL22Yc9V5xNQcZzYO0+z3e0ab8O14DfmvhH4a++HT/C6
+s8ineLwnJQHk0+fcexjujJY7vmXZszWQNr2IWJDkytMzd8X4Zg9v3fsFeLY2EFSUeteAqxPwVrF
qYBwOAVWYqozNBom42WsaE3pb8kIWxUgHlz9BvHWc47CgFzpSl0Osis0Z4iSrgGUQZZYxKeIJhuh
j8qIEy0qdnQSvnjVYtUYvHe1DStT6qWQ/caqI5XTZjwmnK+Rvb3bLXlZbOukI1HEhZKT8zzPNgAP
nQ4ISRyMLdh3CVNGZsUuFOgwNKru3bpNEza86bBpsMH3DxNnnBnMCrJhPpiY9vMns+eQyMg36n5w
7HzC00Naeeo9F/w+4QlYrXGbT7Lz+zLO44eBTCKsLT7/QyKpGRDswiAu9MT5++4yGu6kbVOP8b9e
rhu7esUXTYzSIlgX4NgWWR/3WRbci5JGcgudOVrE7WJ3ntmI+OSTL5brHvQB401Dsptearv9qIbf
WhYxfEgdWKBEp9f2nZOC/b/yujV2TflDHhfKyfQRVkPSh2Cg3xawO0plg1ln7kW+P0SCYUFmhfU6
z15FzPpFQAocrgP/7tp49W9JjgZPLbzsnj8BKhS0r0Ab/dfOC8MwL1bcA3vuBqECnI83ZTxn5REw
lWkK8mB1BcMNoy+h3KMvBAneh1Iol4/eg13g9Ld0JAztEhAJs5d2zw1ccUTURnBj9gdupoOfx/Kf
U3NkZEmNwFVyuQ4OFFv+Tzj5W7bZiBpaHvXFkZ7geLGeYHeQKNMoDN+9tCxR5ZqIatJzG90rULV7
1EM3H7CwmIvWFi4o5zPMfWTeyMYManTlUWjdQCfTgqzzW5ipYLjXG5r8IUmBtG3AxOViY6RpL/k/
qAWY3B52uh3bcrC10j0xCgNlmcpn5vwVGo2SS5zcpJVbdFjnvpZFPRE74VN3BtD4GiAo5MQlbGRJ
C9misB4qWYXI1uT6blN3b0xQsdUJzYw4bdBR0cybrdQjN5AlZcHE3yk4Xvi6Y6ovCkFOd0whT4Hj
Lfe9n/jw6pAV/5BMQ6HALNuoLJfjKsNWM2hqmV9oC776Z1nF/mduXdhWjTelHKtCQijtnjA9AHMc
qNEZFtIzvFvGo+TwRipabWKgUhEdzBtODit7m7pSRIF682qRrolF/9xiV5a3fglKpr1+dKDiHW+7
XY9LZMFxPkedFlr2Rk4rZiAsbYPZYD4Q8HxayNgxequrmakgLYFK0HSYueR/rUX9RybqNq2RkRGF
rJpC3zRdTaojMcxw4ziPDPs7sPRbPbfYguJdoxDDXH1VM49959ycjeMPgq9ABFUhsJjbAELeiN7e
MWtOThEj5vCjRTlY76WsyFxxSfA7n0vt2OdGv6Jh2qA+dM7790cOUWkwKmdWWBQRSGLDrgeaKqGz
AMuL19ihYUC4gHTjZ9ymiplWOW//BxBuyTnvGzcaavwYY01L2qFmx7hxnudOFFUIFrYtbpoQk4cG
Ig6X1/QeILFugE5qHUgg7AHBbsDYcBseRQsypoZMEPn7uRsQrA37Kle0O5dO5G0rKt0awbl4AIIF
TQRzZ99WyJOubbH8LMv88yWDXo6gotP9Bfk3a0i7fVh6WKPvZiSsDtGTnvttdiiAMLOF5oSF+oWB
nFOQ8Ozs4yTqNwNFJkOyTTwCRNJAKylvgRcjp6K35PNfqxMlSmXcQCPCzz+scPwDZpYDogxpx0yY
tLJbXRd4pCQLotrsCX7zi2K8V6yK8YWhcsGAeQvg7EWPU8qiOlsisBQWIXdiZTpR9QZgMVWIRcNa
nWTakhrJxhtsnetRZkCL2fASfU2h0L/o2+Ql0GRnu0rOGKguH7j1ueM2SB5CnRyf321p4MtxUAx7
Oz+sI6GVXbnUyvVh3nPW/rzZFR6qF/Zxh2AR0wzKlA0LksZsfHEBetxil9YHHA/glp2K6a2TXYqX
bMHM2TCY0MFiCfW2OW9mZZqXEp4h0h6oA7gpy4idxg6g7cuyMoZ8h9PHpkrrR9ulD976PcDt4/gw
T4r0rkbZSmlqsmik50DKAjDVtXYuYSL+Y7Lb2ahduh4kccBR5w9JLWK7iJ/K66o5SNpvHkjOHAOI
1sq/xLxhSDydFNF1F/j1E0rpFQupDHjVE8s9iV0O2EwFFkHKHL/plhceSFpRo5SJfGzfJBYC8j6v
m5M9d6KRhC6sqDU0OOIA+/GcqiNi5xfloi3HfCBscWgl+uVYRnFFBcawAWQLybtm+Ebk5TnhzX47
7+VbnQ2x2IR6zvlSGke2EKZWBcVsQCn1xNvCa/tVAj9BMlLF1akFbCe7f0GAY3XlQM4Gfp8MYvyG
9Mj7CHI0KXnO1URno1rAc1tImzAozXaJGmZNTGgoX4+Q2SqmU+8Su14tCUMpEmKNimlNuw12Tsjm
JuH+LUGH+zTbQaFkt1ePghKQHjmzubzDpF7q+TXP5uj7B9t9qykVxEmsCHG0tAm8KvzGGGnE7g1B
HuWznmJ0Fq/L7i0YQSEyt8DNRmdpk2vxAd/SlrY62HziCXbRNZvR5hhpwvYzBFA64BmU4EPn/ygN
7xe+lltWNdBLDVFprxS8ogtRlg33N6OXg+U044y8irB00LKfBARBpO9tkWcm59te93djSeNn4uJu
CSCma5dLX6kYRQJqdXlh252tucdPxJcsVf8/yceuvv1h8c5q/3oE3R7/l8JoUkLIBd+YD9YI0Fjo
JT5NzijxBEMPH5NWJKy9AArzyfPWN56d0sh4T+sLJ5zsbJSgL2AvSPIwYD74JZHbqsofkfSPzv7T
uOi/qVSxU7DdJC2ooJFT7ydXb28cuZHrkZ8Y4Z+R8EyZxRmYy0dWIDzXHj3iEl0n9pCoMebQoRU9
NPDV/ekFY05XWXQ5iQIC0wEdsCloolbOttTDYnkzAWByLmbmX4W0zBXK8ORmnkv5E5TuVrxZoSm9
frspS72XPkKuxDUdH7CfPekTvkah3TDaDfBL3tRuRxTiXO+/jf/9Na+0DdHzU9qB+UfhY0QB8d9h
ofXJStIyT1wmr4IdMQfWk3qrVT0hk+FmnXoSj8yMMRX4Ouq4awYw7lC9wwISiokSLbRjGq4jg8Qr
WqsHdP3AviJIsmnlGz3b9ThAIm2zVxeEvs062jAEw3DDbtXIlwQz/msj0/GmnWBEwZ0Q0zdNypTc
4FR289Y09xmYtPwJlqp0mbFwbvr5DLKd7itvDGeYa3O36d66ul6Y/dP/55MarxqCaENo2WQXPNuB
2I12+USxVBApWFmTMM36mhPoNQz5X7cKu6HhdkHvwfwzfwtaOA1YQ3BmipaGa1WWCfGbQshXaDV9
f67/+rCGge/Vi+gpH47OydBcBD7hTyNYWM6LLzK3NtJrAgSqy7U3e6f4I7gL0qTuHionDRGhlJ6Y
wzNHvDHkEVezUJ1rywrqLK+wEZSVsfz+LvDenCHGsmMydKcR0KK52KuiQmRh2SFhuZUGWrUHOZkL
hVGGysqpndCucvIrUE08XZm3/E/SMxI6U7QdqK6jcY4yTJyH8N0a0XJ+5m5aTwm7Xfb+LBBqcLs3
gsYhU0WGnjdn0Jw1CNxdUHwuLWn2w0L0Re+QaJDezU2F2d06D2vnJYlGZ7ndYhgWab0dUMXSUUDn
sdfSHfso3OdchmzFA2S+Wp3RSLFZPGFki8Y7lKl+Iy3KfTASxM90WncV/cSx6Mw4IhIpY3WnM15m
/0HAj3XhZjbPxspmY2PhaT7iG1a1coKUOEeSSraOVLbQSwUNIw1eTGyQtvEUXG/yX5uX/MiHjTtQ
NREiipqVeBSWGt7w62yFhoUimcaC/yCpxaQVOPZSmxy3Li0YYJei0WBrnGTcIcIA4pgcwWIFz7aV
tVtJSCpxwy5E6MZlYNWrGRDQa+7eAReRe93wqgEpqM66Z7ftDTuMr5H+lkA/+YOzOin4wHvmEJea
bJb0qYUxq6atW9Az9hoveONCGSWpvvRfhlf+s12paOBFlejOas6aW1fJIzKlO779znvUVPPaLo+/
4bA7SOa8dZuTeRjeX3rPwXRveJFFFKwjuSeTEkDsEgEPIoDNRg6ULMia+5rxuELYM5kb0XwTSQON
pNklw7mVPElpWEI5Nm19KzJ+u6C/q+KhXcHIZ44ZiRGrMtYrHTwbK6pgWVKvW68JhOIn3VnpA7YQ
eI0N6OUgtLaUgmnNcPcCDEcAsTCM9rwdMntTx7ZdUG1xre7i2w/9LrQoOow5Y4BtVCs1Lp6pAXDh
IBDR5H3LQ3oz9NBl7CXEpyCDdJG6hfivsLgZdo7V7z9IdUvLmdbYuwgkYLoIeZb+tjcRVMELAchX
sz/idubavSsl4AuFz7LyB7yRPyzsGEwVbakLYMRZyxDtYux6bk3V5aSVyVAbGxyqugG/d6FrICXK
nT/BwyZCoBQvMk+y/cpY4f0mWJ9K/CaXrFNpj2l2q+Oop3K48vXxrOE2nK5OcACc/tzwKkVFRnMM
1JVd4DJUP2AZOC6fjQEk/dAvhxH0YLVnoLlReEKeOZXVlNY8UWZOBrg4sQmSecOIUn19lJKgJUkH
Sp8ZTYldDIUvIiu3qllm9TW+saxBfQVvVp0XwcuPrT9UJmlusUM1lh9pQgeZpLzwH9w02zr1OLLC
1oYSsPyd/XUJD73osSMY0govmK5oiy2OeNg8NDQPpBAloy7toK6OKPzEOZfpalWGsgobaClSs2Ht
NMsmDaJCGzkn8RyO3Ep8HU17XmO2yTuKf6+BvcdlP9TH+eherdflWbsDn7D48UFdkhnMS77WbVyF
7AWtZ+4yLSaSdsenGaYaM8U1kUailOfovtRa+fRsd/WT3qN1xOEIOlxoSSn0YBRUzf2S+RcfjY/b
zzwQza3Xw0e5zF9Jjf8MtdIvpkPu+iizdyDIyZv1Hl72BMqMREyhaEdtphwEU5RgcL/isTYqY/Rq
U/FgzhuabsvTsp5HMG3qOB9+zPnuO1Ej030VG+tS2FuRx86qKX8BSola8feB9WR2MZww9yqe6fWF
LHei29aTP1tlZsnS5jJ7Re2uHwSFjpCm2lrv8PmSnbX/VOXKzJJuPZkU4SdtuvfxNrAJVnDSVEA7
Lssicu1bMOpDyZ4wYfdI5VZP0fEL8BDLQ9DPq761YlOsAXPG3wezo+oAQuQnx/sq75dc/Nh+cZI8
UwZ5YYbuik1exV+rnPyvXQ9LnXOyMlXzF0C8bdZkVzkPUz7InqPy/TmEB6aLJ1UwzeHlBiFaPyoe
nIwpmA8aqslZB59rJ0gHgw2hxpymnXR+uoyT+D/E5F4UXtNEOavE/TzD0kpA2MPaz7WNQeqQ2aJm
E1BGPiZCtVTunD8opZV9B4Et8ZkLAtNP5KdID8A9EfPT6BvJnYtCuS4IoT6h8S09puTWx0RX4tPq
uHQbPRY9AmvMtzJZ7lv4NiuOieAik5Xu9VlQKub0jnWp7ah3MJ9pmTbyqwBO0FGFCIdDVey1SlsF
HxLhmpIqrYtYLrT8kflnK2Md0+iWzodM8Hkp1MODgnNAwAsxUbaTlibuOYUOW96dzJ1OfW2m3nCz
7vdUdQwxpNjxAMbaWFAmLOWgJzT2+SU02uGYYQaLjglNFStMHHq4Ud3Jr0Hcuic70fH7MBC9BAbx
JPPJiJ2r5pi396uewOhjtthZzB8hf9KE3CK1/1dv+T8xlXORJmwmBNdFqYGvGcIc8nD0YJ/fVTEY
0QN4F6iTByswCX5YQ2ArGiLfltDm8B1Wq88R6HiZ50b7C5H12pw8TebE3o1PHvJlA/DzN6t/pN/T
iKtYdIzByg02LhrSzT4UIuwQpzxnyU0rpDWdwbLiwUBe+Slxj7Avzed2psCnhcJ4WdT+TyEp32zz
rcTTLAvLNNjcXUvj7z3C0znuc+fmFL9fVL/fm+SmLx8k+MWn4Oy0cyrCFt8OvMh9XjbKlFSt9Gz7
O9Dudy69W6JtP3ic7ThtkYUthNhm29aQgm+dSOEqtL8zhjWJtaJovTJmrl1FOYNb7wKUvykVlvam
dn/lDiauUWgP4mRaCXtNEtWts+Br3ZXpXFFux+a+92b54KeTTeDQwfaxS9jhF2BNhxC6bMCRAOLw
cRqPjfUUQCL/cBfOu6+rGcu/4M21misPEj18+IsS48NTepF2IqIEPkRZUa7P3wnZHB+aXgNYkOkI
MQ9Ech5cqGjKITBOt5/Ha2ykcveLz5AvJdtxZT7EjmY5QRI8k6Dr3WisENpkr79OtiHtMpvHlC75
Ft6gY8C3IZO5nZNEjTvrKHfjfMp3IkCm6OVJXiUkLmitqmOXiJMCkoNKYsmB+ipDzzuQzx0+zevO
Lc9SsX1cm55h8z7RqQELKrWGFoyVKC7cMYmZ+9K5shJss8kKJFYdN7tB0FZC0D9kENJi58v0mvY4
Q4590qqpzl8sOioqgt6nKAY1U1MI/q+PzY/Nh0pOrMG3Fpb5fhYoZxiMU/fEXcxOmP7bA052BOHM
Dl4ZpOgvbaROZyY6pC2ph4L91HOyJUYQRwGunyc9OPPX5+WUXtEswZxm3BdDzHXN6rB1KtwhRAo3
gcO3i9+rsR2YG4g47kD418O37i8nVPDXhr2yEZRm3zaoos+gNWJkMTtQZ1Rl15Z0rmKwgRKdeWZH
qaaH7Vw8nPcfxn7II3O2+IshMit0b7GgfbhrBiCc0q/VHFUuYgg/Zhpe7sP9efYkuvDbRaO4lOf0
q41zGxoaibDMnHNkvi1hFazkL+FJZ+5M/1XWZc60U5tXKmzbnxDBPRWtHpO6EnQE1LpD3LBVbyDf
455JfQIkeIhMt9rvCUFVOTNnNIZwmoBz/NKzWll9xgbgZearnKMg9aiuSjfqokQSvlpKeN0EAe15
FVs7EIhg5SIoC1HK93mSS1nKUyubhTbnenVv70dzC31sG7G3PV/AcwTHRCP0H2CBjyyg/+vc08Vc
ah9M8THjajV2c1ms+GJPCMje6yveEIwMpWSjGDwo45zM/hzmwrreSK+VZv9dvbcFvV3R/zncr66u
1U75i/ZcGz1k7rH9h9D82tMPhqGQ++7FQkdUNgeTfsDF5m5nA6OcXh8Wlfdasdn84fXxkPns+nLH
HHuA74DNsU33/MIUxspDo3P7ndhGo1FQsOkkhU+hVgmHc9JLQ0AOci5i3tIPRXXQ3oZJNcXt8aNR
miEiaAcZ77YWOw5/4x3Y1KBNVQB7HqXM2fpEI3n4DwrDBsBtqxQvTKrn6JZVS37fGYDaAdYv2my2
fX8ty3qFmn/ymnXto1guWzuN2kvWCOcSNu5Iw63TWmNBs10d9DrF3NWX1/4/xqDxCgjH50S6P+yt
mQMpX3avg62Xq2gMEHKe0axmVQ8OXR5TVwcBA6pkE3LSsUxibnMyUHPcA9FzoviPsvbK6piSHBiB
qXJYy3v/8Y31qKYVHpxh4yXjYrzZrZXAE4gwBlW38WpqcUTyPCPlQ2ziNkEdEKgM/DNs0kcvHK6L
zKu5cnD/WpHmkW+CQP6XVWsoJSKlAty8yG0oa9MgPzNSRIjqCZN3zC9DhHGjqP8WNSO/Jdw0NRwj
iosyQXwRs9HCDziYh5ASlCF2fzRZyancUVCei/rM5y5GGjiT0LQYF3WEKomaJm1/QPZnnzS+ZlgG
oG2tF+CHTDwIFE8eKpdPEc/7mf8P9bjODlVRw2//pbsALIy+BYEiyXlanrf9OeZqgVYOC+rof+tA
vjJ0Xv6pU5aqlSf1cEFw9lbeXyOdF4ndT7IcyuW33Ym7OwqLnlDT0bRUXT2Pez//UYYMeXqNxd+S
v9SuFQtICravOFn1R0iSAhjzkDmRPxQMcZ+0afTSLnJIU5MUhUYAmw88U0qjlYfHq73k7jnJk1dj
LmiU8fmjBIAE1nPb38c/3qUbfq4hFxlbuhz/X1zqsYLWrayE+iuPUqdlg+VVgrPDIeknAoY1aqX0
vZEmkFf1AZsaI1iSE3ZP/0lrmRm2jUnoDMNiEP8fnK9qzAb/9nSWqKRScCGpd4ySfLpOIGMmPbZD
1scS4m6sJQBbhX6NmBsU6voMm9QcKVchDjMu7jKmrodpttb4odzggPPdtjZVIey1iaDl5YFlWBpW
hJV8aMgRR0+xjE2E+sIL6vDFVeSJuIVhYMIiNNUNH+g31fc24k73FSAh4gVhrvDlCktjnswRVCB5
5dqkGs+EK6LP5xHq4JDKyCSVzNIy296f8cF3hPnPRvXYS5zbqmPHCaZL1v48ijv2cWLtPepgYu1e
8j/wSVLwrx2D91sPiZpEEVJrFcNfEOVou4CVCM8g1DYb5CTTW4ZWLrk5ylZJeSa0/VB/Fkvw6rtO
MvfInMDvA1oecVZVWH5DlhzxN6ExNmh4ooarF3yorEcgduGzcFseNx1aUWo9DNuZHEcYk8ntcTmb
f+qq8S0fsR2ikA1KMKw2zrVqPojF2QjK59zKUMl88HSR3bEdIwnIOs32Bf7CIF47OG16ezTsso38
+xv8o3QbJI61T+Bh8P0yHZqXmwwneMQYUbBtDZyE0pg+9HP/MJJdSJB5hzDKCZiHiSjvJCzodY7W
EFGfPnbuOhcS1zEcNT4K9JLMyVuS7whp5mXmbk33OgX8MI6aT3n3pWGZuzBtnLILpgGFg/ATV/qc
s0bFpy0T60snBR4Mq09Jlcb3i0x9wBUX0ZLcXw18Y3jbpNZPzBJJtmMN9KbIKLvWaLPlWC3InADW
yxVOlx1+nqdJLtvTycm+0RzB1OP21se0pd51mMofTm0lGaCnUxr/ewX9CmWgbx1Rvc0/pkbor+ae
N0Lyb+aGa02bbXCJnPs0b2X2K05xQLw0qWbJeCvVWPUN9JnuiEL4Io4wz/AmgsBSSOyN38yRwkPH
nSaB5v+2+UkbW7vPqJTrWm3kKTW5a2hyHc8mWd5kq9mTxXC0MYCeqWIRC+gz25R0Ruy1YuUmc9uM
0Hlqj24NBqRqyRQmFbBYaKOffaeJLcwKbDuHZ8Bgl9dE+yPFfLNVfccpJUolTBQuOrfx7qREv+87
S//7FY3LoOy8lZR99UGQCfueX9gdQ7B2kZhvjl1pxVubf+WmnNU9iq5pPhzrLyIQYnGqzhEhzYE4
GnxDCL7NbVk1pA8h/OQTu+cdVYMLJhzzBKsoU6ZE2ntQQPXsf2PYp5EtoKPLDT1HUHhbjeMQBDTD
WGLVcTZRmp7FIEKd4FJFm+D3SmXuRYW3DQGwtP7FFdMDUWkVePiR29gbf3ydRgvrVTxm+SaeHPnw
5x1ZdtUR7+nBv+SmYwRxmBrLku+vXCLq0toDW1/WErszsBJfal8hzEfkA68frn0uaV4SWSQTcaJx
ZzoVpYfhKmU508YaLHwgQNDv9Pkw0g7BTXLs1C7Cifra7J5wry71+OURXoTJ4ldqI/lWAJQwfPue
t8Q2CDHJyGc0CpjY8vskH56BG7R8CUXohFo9G1pq780sEQMG99ICh7Wb2WISkGhk0MnK90eYcwsb
DVxCJaShpY0pgL5ZbiuFKSG+jvgjOI1RNdfIHof839d/u6TnSwjaMoDxJZdGxvwOyzNBfQVa6qph
K5nMsJiPvr/seJOlq5tit50QD5njU/QftzSBGMKAu8twS8Lrt8fD7gs53/FSE1DpW0jw2ac40gxj
0mmq+iUlnfQ4m/tqKI9RqBtPuvdPiHo3DyPQEfYQe3gqm2jKW+dR8bej08f9UP/iM9Duo9ygbz51
scdFaUnEulPnGjK/NoU3J5yeW+yu7GYyMwzGRwgfPpwxpc9FWX1gnhK1j/SWWjJeS19JDfGmb6z8
xIBT0cgbcd3ALQMPQnj/NCh/yii19//gVhRJTJaGEjKLREynpqGP4nt8/69PuSo1R+oyzP/ZBzG3
aDDMbRQ7G5LqPX/xvRYps2/4DTr8DvJyLEA1uLX1oUwTRUfe3FaIfNmgvnpSk6XPNkKl+niAvvPM
TghtOgJcvPr2PYEulEMFXZ7jyFQ7s4NxjwfN6rwCDSP68yOStSadw31gJJHDHEjEpn0kLSWUdbkR
rYyMCbmYLi5NDDWGrGK7fT1+GVK6hJXGovA+7sGVWy5qEs9cjjLQpwUXCeoHUSN6UWXzVeoeyr2B
HAS+pjGsoq0/d9+HLI8ZgatBserwf1zkz5YyyCf+I/Hekjwuqt0n8qg7yvDpYYAlc0s2RrRGcMtB
USZJTUy0stzL35jWsYT/aYEZCB0qVfc3JuEeqwt0L/WTL9+YGF6E9IhtGTJm+JEnDdENXWEGkZ7f
uhISRmG49uf7yVXVoSYOXEJu8FOrN6ZqtWyuB0KERkxFE3FUSqIjK3bYhE7R43zbVt+YuhrAvBYr
jtJq2kGGkH4zmoUI3+7IfIO/4SmOCqQQHHXHxaGb4UhUAdIRBn5U6ZFjDnHyu/0fLeQe0nE7bxbH
fxte0fZskdVXtI1Z7111NIWH1rBkiNMZjn5UcDgPbBDUc52UuwCnb91IHYiRIdatYli9Z+u0XT9x
mElgwdx8+YWHTLx4vL+faVhGPQqb8HYIosBHGqpNFNt3/hXWYo01/zSrNzPU+itrwOBJnJlW6XBI
XYZJmtvAPssPd4r4ZzHBzNpvRIeDF82v02zTyaLxW1Exh64cbvRQecMebMYV2R+ASpy+QMbwaWGy
UQ2BJKONCUI5jaV6u/WZWTctGEulWCFs7uNDzDSzkynjoFOHKejK0uV75aE4d6MJ6elHSqUDdDv0
sm2bsS02yL3IZPlppxdk9fzR+JoDgGHVTqOZHk6i8mRs8jwu3g++nmpZWjTL2Fnx1mpMm30rrIeA
2PRDmXWz/2g/WDIzqAGl2HiucFZB2JqWBjAxf4/wW2awV58aZvYPuv/+FzScqrSZs98osAFiruhM
zaqMkrgp8f67CMPnvTYI+J6RIFlYb2W3cqYmypWZZ7ExBn7qIOvgYgCuALIt1AtJjiqDNm0vHgwo
g0AsumDqjObCxy0Ot9fy7B8+dyopP5+RbqM0N8VmN7W6ZOLiWZzEauqvB4w5815e5l0taS8fvMjy
T0n3+7jb8cf4/Lp/SW37kD2VOyyX2Dm3Z/psYeojauiGCwSPxWcuYSbh9hAzfTGHxdeAI5BHzpWS
zvquGDgrjJxDSVXPgB4+dUiasxfBSQXtdr+FO4cKUUCjKFHEtqS+HXYujwEyBcr/yxgbCJTpQly3
aanTxdatJuwfQiMXrgH76XtF6OE9z82n/fNzn06PaJmovKTzFTt02XtpNxlW/GVg7JpLZ+HJvJi8
zJ2swXpEdvcpsXc2TyusyH0MsHszmtkNFPK08p/uNkVwNMr9chkwmRtU9UaPkCQzvzpzyHGIPu3O
lIPaA1yStUXr9IKlSUH45lbta+QPSHQ71exJlh9fasts00AXTagPILH+6/i+voD5fztW2+G8QjxH
LpNwFAsoMpIqukz+8FxLGN1OgCXry/XuQ0EosTaezuaYk/8kvFfrOqKDMv5ZFvDNugmkK8e51lH1
SlRRY4+eKXjZTeQfRjpEfJctAeCmGeTzAqAvu+sFNMSP11VVsWR4DT5Aps6qysVarM6iEfYSD5Nm
7sM5ax0fyAQQFG/oTxBYiiDB8Ex80sa2zb70036TTg8Nu1PuTp6NZsaFMgy3OhFLv3TnhQQTFt8F
A3PEcdULPkuhQoUVj3d/dnJDOkK3mOQp+AwYrED8TeRz4pAKUNigt0JDV9sM3rV3FxORhNNFJX4h
TfeHIUf+N2YlG9PRQQzmGw+J8LOvjVQC+B1zadA/Zb7BU1YkLh5VAemA9L+1LFx9AcGPpxHl6pHl
tXhnzOzVuTHc4wx6OTgsWVre/IzDGET+IELp2/EHy+S/uhTEOSTGMFFR5SYbOPxN2H12NGY8tIV2
CI9grab06LskxN1Fi67SaVOA3ZXWkR6oxtyvWaF8v2ZgbD03HL0AGmvU00oGZwEWBSZHMUz9wRQ1
bngb3KS0XFgDU+7el0OSUThhZsVBvtx0XDqa2pIN3hJhk4DYytHULMqqfzFOKXQZHyuDccgOnTf4
+Y1VGDySMYnT2Ez5f1FWC3nkPOR0fS6guj9qqoeDjAG/CHYwC6xds6fg2vEulaKyrBNKn21oZtrg
mV6dqN2GQ6/TGllbq23x2KHZcxvxA5YE5f6ShZHY4o3rC/UucJPdYp+ykTtMDYLq+trJRcPQQlBz
ZaMOJPt02AvBXURrD1jG2JVfk9Vyu9onRyTmzSty9Q83mcpDn3RfpL7FWImjVSD2JpA1AHRUDG6J
Ii5Hg2CrJpBJ+Jo6SzPavKUzicGu/u1W5SkV0lyhrKYfFsDdws0ZXGFlEPFwDgiDW8DhTmlXGcZz
TkPmGRgBdI0urGJFruT5o889n06eN/SCr3Fpm/NI9HoaS4/AUp3b4ksEMkMwyqWun8WghCX3QxDU
7hqRp8rDbKErCvXXS1V957u11oN/o2FloC7amTpijSyrLppjAGawSa9jsws7wVuXIwcZsRRnq72W
bU1SlFXjtknKuArdZdBV2T7ljqAYvl72lh08RrccyhwDobWktm36Ip9VfiQtjbVwl+/2CuxSJKey
5VNIdKbpxTuPjamkZ+vS3p9RmLZpC11BXT4yRN+PdtiNIvSfaLSRPZC9S19b+WtWqfkz2pqHSvcX
0xWOw0B8yT97Yz1c9FEZEQ0gM+bOEPUfbIBfJH+AJgfGlILwwnHgkTu/6RIX65zW4a//ciVk8F2t
inlKMeEh6KlL2lFyYoPs1xSueWNchBxD/+9nO8ybmYi7JjNzJLdDbT0yYjAa5mUh+GgRTNH7AvA9
nBZ2zYOeMQRSih10gXVS6ZJ9nU2wVdTNZCvRbNvxX9V1OGdm1tKtY8+NLZoQqVBtTxRLy/tipSBv
HuTAItNBa1cdHeEpRAwMSOyvZIvAFpQzYgsYovi8wNDIAtQV1ghbGaIH9SF6sY4phI+1RXhvWWMa
hopeU4TE7aayawO0cPZhrcWct85lgqYsvQAk7gbWImXuYz6OTCBj0n94yqgSCdbhHXyPXjtavtrJ
svmHaZBCyxwSMCTXxRhKKwau7fNS0/h/tAr5WhxF1RBvmdviYXbVMPyW7TYfqKwBNJx02fkh1BXy
Yzmmn25/CeF7GeTRSl/WqBOcIikTsuIHORloX/zUCYwKrvlR1u7i94qlf3wFmZ9p9Q0+I6q2Cc10
Rs5y7fSI6JTsBenW0hW20oIa8LV+hrvrEIf/JUbG1rYmDHm3G3zcwcc2pyLxFJoZRwPfjqwO7p45
fgclZROpjlzD51bVtNbXHdgaODHFQRk8rh/22SsHzLIfryhTn+8aurmZGataN+xnINAR0z0DLZua
+RphqhFVwWB31/PW+BaFM56xIfGQ1nxhVg+OYp8w1h6t++wVLXgQFRqK8vY2OXdWvyD4eURooq2b
W15Tu+1JO77CNNuelL+8W/A5l8jlmCT6hWjBBLTIy4WbHsGdRZuqQU/Udndk1xcfktMDf1xykOE2
4F+VqksjjhcO4ZaZ+NTT6lwPcLwbCHSSuUKuk2mlnvFRcBiXsVk4T0Fw47WMIVd58J2vPncIt/fY
xsH3kh4OWFUX9JKg3IWLmnvDlhr4TQK/MDXS64JOIg5A/0lXK6/agjbGT2LxEJ0ly+C5s9+U4Tpu
LClDBGlrUsKzmsjvUpjPXYDMIFxu1i2bMfz50koEAQC+Y7zIC07qynVvIQz0+c8kHHe5NOX2QB8O
KifodMgHKj3Cg3892qEEhNl96ftkSZ04le61Qi+MdqJ6mBOqaFN98cXe2SSJh51RzocvafLowXWP
v/nj/wSjbvW57GYC32L2FeJGyy/17zCMg5b5M0DZPyWu4iEl8FBG5XaGR0weDFngC9ktCkfQcLte
ZQ0PRJh/Xa7wEFvTAora/S6ANl+CMO5bg4a1cRVRK0gzq70AA9TZ7V2KM/62qJ3II3FyCU3H0SrC
OvN5ApfWoQVIix9ByYNBH+AhVKizs1qw361ojQ5FCf8Oqg8OIitaVy2wGkfk6L8unh4BaX+7185l
5vrRd0HBQukjZS737xsqEj4Z9n941rvubLRgWyYelBhneBpSm2HZlq6fG3rO7zJgXm5tgFy+ilBA
tMrz96GoJSDBgVUsO5HfLYVsKCvwwQPi6v28TjwP6SB5wUZ5gG8zVTi4bBg54KEH2fYQVoCtucbv
CabwIjal/Pyc0KdWct8gMihJrcI4XG8I8063OXymtFUuJB29BuJr1ZlXqwdGh8mfR35MICa1Zr6m
SqQE2pzF7Gd4w92K8buLNlar3og2AuXWPX6AJzt7nqt5NgB54HyST7UozolCrIuHHigOBDX5Tx3R
OePeFa9J3CaCzPsHuwgsc4Qt1KRGUcQd93Yn8fezBCVLy9FoT/k/VZoyFws2Zh15hoAUwhIJjRTj
8KntbOkFDI7qWZUOf/hw7ldWR2SwaFQ+XQ7gdqHO3C5LeN2I0OwsoHXcRAFVcnVD2eglUZuwrvts
arYgFCjjEFv9jnpcBT64QCpn/6MiwBc0GxtwAhM+RwHwIE3oPdQs2btnoUkZ7wd9LwO8oOjB3I7g
jGiUHnMxA8pZlB/+atGhVK5cNzRkArgvAH9AqvBmJlI3Fhx9sgOAAQse2ttSt/juLm2DS4JL9sOS
CnOZxaget3IvZrRN3B39qQER+xWZQIL7YPuNg72Y6D724WB6N+zutgG6qy/DwRAh7JSlqOZrymeg
nmw+xLkBKt9e5FlWRU1ihQHBcAL5UD66ajd1YY1NvfOE19tW+T27QxjUQYqagYOmdi91wkYA3SZb
65GcAsji8SYUcs5yLnEgrNmNKI/KSrgnKoTbyPzEbMJ+A26fLKep4QcuNyJBXV+O+nxQ8+yJFW9f
C3T1PILiss8wzolUUtstAI56uN87w4AzawQEiOH91uOnysmjUlvntNGiViDLvzsHt0SbrD9l90bU
WLUFzeNOdaFMrH4tgDBmDefnNDhWGZm+Bx4y/YFfdDoMLIULylKNFqki7S5qZ2mqqyJgHVo3VToW
njvJpdcfU5wuhM3jSuRCGCsTasCG7lg+qH447UY3EhRK3XIiT9BDZtFQmYgedqKjIP7nLMekUWKc
NtARKY2CECDraDN4ojBNH1Vl3zKm1/ncHG/HlYMChkz7pPqKYINmd3YrdPKY2t5pqJsdIaNd3fD7
wcms+KkFJSd0zywuXCBXJoArrDlliMo5E93fNgR1RFJsRgMyJhpA3+RVPAm83/wxxNNZHOBkEpXu
do/kioMi3gxjIKhMA+H/3Vlt49e67kSknBYp5r+DcdLo83bx/1sweZHSX1VLco4Mn63ar1XZX4d/
XwtgHCRlJVOp+NMFeEM8JaoyRplAzpVRC3q7gBKMB9lU901RHzCHKdMVazDc0fFo1pnAJW9uPGD6
oxgjxzFvs7vA9YZniZETnjaBJKsvIj+TXBk96pnFU53KCioR98zCMQ9zbpUDGCnYY6C9jM/bjPHu
s8oqYXCdwHmg5kSLT7NzWdUBWGZ9jDxMapIL0S3QRWCXtKSjkRvwMOC3trEto6OjdxZBKnGIzVQe
VpmMBx8nwNXD/Vz+/tSpAr1W1iFhdFIhfjE3J8j7J4C88ztRDtFLhlnUitjqbHhvJeWbE8ES1Qys
D+l2pLC4+7INVmRAJUKfr874BayXmEsuF+DfM+kdC3qvjqKACLMbaj/wd5S9al9szO+dvFyhuVXK
gwmZlu7LAlrIdyfGBHT5v1UQOF3C0wzGA2cwu6YrAY9NYmCFhZuKwjaCZeo2sQu4YNwCesht0ATd
yMvHXfqMXUYAmfa2bsuWjU/VaRVDaLNd7tIBOqXa6A7XMmr6rfDOdwEMoVOEnZ3KOYfQyoBBN2FB
lHrbOL2Q097/PKOFJVCI2+6+woqjuAwsR/tC9ArdMZX9hTY/3YqNXlQmqQvoVDvLFvf5zOOmcPVe
6ZU5uBVUqgM1MhOSPbssQq8p4xRz/Y0UNornOfUL3ZOEg1A+vIQIF6RVCK1vATXmiJRRo+TkjCy4
Ri3WQ+HLMPe7fSf/hA0lCZjFaBCuvHxXYnh16/0NHNfSrmqqIIfnfype5WuFQ471JzkNoBUzlbF3
S2DuuBdfwyLO4Qng0/G/5RuK3ZYCWboi/seDoJE4/8n6Md/O6WRveb0oEp+NRdp82K5/g6/dCf91
bPGiZTbcwTGCv92+i4dV4+in5y65LmYyITq7EctDoKLlU+l2ZDr/FZW5IU+s9JTxiiWkwiPnPTyC
yQHAeY9Cm73I9WdqKGS60e6whfqD+LPRf3MAYbdADzIJVvATr+3/eMHq6CwEZGKNVhmehAa+4t96
N/KK3Ewz+1ra3xmeWldSiOy7oaSZT7/gU4Lx+84dxKkD8ltBefvyGdAFA3e4saVmVbVABHKR8w0k
1Gf+6iLYWB6E/ns1lTnn/EDdMk8WQTCU9DgufrD/UiTpotOyyzU7eAVGmdDMmWur8+P6zlDfRyww
rOKp00QKDFDSfun4eU3HA5kWa0FPDy8Las+poYjRXtUyuatwS+o0Qyy0xYe+84Ca6heGHg4EOoon
DHomYCy1O0okA293Tacxn0HY9SN8gPW60YbPMjhfwAlHepiMnrO4DD0E9PDMFu8SrpAJrUSCXrN/
rOlIIsKHBbNA8dK5qraEdcCK/dbW8VMByQJ8dTqIbjw/a1imgDWL2KAbAE6fk/UYlLc/ZSgvnOyA
NGszP5H2sb6YDWYfqKme6swodp7lUXajR1ez/nVTDDWb/diGbvraBJMhpDpH4DBIm9lS89WvRvio
hb1qWSFhCk0XrmITyAAbftUDv7jpXkYMS2amAMCTdW56WPFeVpupd4sTArXTAMJb3MmR8NLJyD/l
BJvmEebXwnpzgRcBW15ZFMp9h2a257keC6YlyFQbtuRmJtsTwOQosjRGeY4/4cmN3tauzEKxhPbE
FVUxr2ifNQx2d/J3MuqS8zHkoHZFQOpsXMuTNZJW/I+MC7Y2apqnRAHsjSBOZ7UEGRPy/zyqTOhu
SylrlM6/m4NQrUlhBKMevfm2JoGu7QCw4732YK5dijzqgMMdnnc3GmL56149uMOy+vqq14AR04In
3gktmv4dnNk9DH2E/RzYbn1RVi/m+u7GMaYjm4z59PAIraAXJ/0uI6/Hiy8L/4zjqJgDoEVOCLEa
T1txLVj2sTjU9kA4KttsJ7kZgBHwXtRmETvmwLzfHG72Q7xNOLnW6Q3ZLFsW0InjRbKKFMZug0e7
14wkSXQC5BDt+SxMV6C6WOXkZ9pZRCMwm1P/6e/YJAgSZwr+qG0jWHj7WisM8fljHXCkSsKE3O8m
EvVho6XRgn+tYFGiDB2JKCQDUCIQ4m8BHNDoMbBA5uH2+J0U7Nm08C9TqUW5zA1dxYjyUb6kxBJI
a0XhdlZ2o6dVRJUTAb8TGkbGLbPvYLktyn22+Uf+bHX3FGKQ87hyv78gfude9T57K7lP1+3H17Mh
YWOTAUoeT7ZGWCjB+M+n/NLYbcbuKrIoYGGg+MeH++xC+kBusRIHADtLTMfEj+m3m/F3Bw6eTRfi
RPfC5CvJ9UItseNI0RPwN58BivlkhxYww7GkxsbKw+gpTH7sgE43cW36Krh1mTPcb55GOEKjHEEa
0sTheBlFn5KVcfQnfRcUqF7vzQIcVxkUpfIvMtj7qPIPbHfaDoONityIbI+pyjp3uS4AskZ+lzPt
bspjqLvlpPeyp/ZW/Ah39cFFffm4ZTAJjYAeok2Q7ACRSf4tyGWna44z/wGMjP4+GeNuPEe43hhZ
6E6DqgNMEXAgV2VlnHeyq5jvV6+4orR3TiCnawppjVN90ooG5svlXXSrVQR+b7gSTWvSCuBJ1Swe
nNUTnffNxLPak3Z/3iooE7D9Tb3IJjspaG/X4X3K0XubT36WP+ls4EMxh0l1YpgKBq1vySFWdoey
Vvn/fCPnsxIrCNOTu6Tf64J6+u6hY+4vkj/H6wHNh+PLZ5bj8DOnp76cksrabjqk63RqUe+pVOBY
toE4DUkSK52yESJL6XjN/XSu1Rw3XqD1s8e4W9bPpSd5Es5scbvlOtWLW4uQX0fJpGszS23f9LbK
0DHeWjpmZ0I/FYX1htBfkqo/uVgzMMy9ccQN8Rq2k9dzUU2Ahq0jRZkP7whxy36/kCfJhMNhKZUj
/AuKQmuKn8pfN8TEixvuy7cCxJJo63BdyDIFQyys7Jz2sPEGcdIRLKQfuTHtvhJsXrbk+9QVTGih
K0xqvI9SdOewuEGabhdacBzETYhlE7LRcj/e6buFXOg1/sbX6wiJHcKOhjIIv0Wds+JEyWEUWe6m
fF9r1AgFMAlXkKti2JhsyqsqQsneG780x/kZ6YCe21Qb+NTOQ3iZKmr+uxQYrKBO6mkkBRpsaEJp
H4/7pWQk2beuxGDa7upkZLaYbnLe3WWzevROfVDzQ+29WeXdRe4we9uooT+ol9ungEi9baayDDON
XS9UwZh2Y5RVzFepulIFpsNvmgSVNH7UmO3ASsr7ddS4gPFyoSQkSUE04PdodGXar6YcVJS6WKs3
yc3A8o1sM1pLtVDu9QmyzbirBhjfLiXfzaEYSlGqIRgY9o7psbX/kF8qgLAiGmeJACihpC4cK5x2
C5w5dEb6CefHX3FiuZ9Ni9m1yr9a98fMtmVMpUnLuk2wpWT0/fNwzL3RwSTO+NoPtCrWS/HSTb0t
uq5uVPJ7f4vEKrLBOeDkuPnE8lZ/+j4/rB07v5lhEIi4W5/FpNOUus4TvGdmlfj3+nNXsqNxQjGw
QT0KHY8Un3jUbpu/L5DYBpPl6BVt5FaZ6UwWbqVILfj5t/ykI+2V0aVbzm6vwjaDalmuvflzWrZX
RHT+S25Rz0/rsn6540FF6r3vdf06BzvNbO/8auzJHTGHm5zrVUwBlJxCFkgrBJnSyUroTLjJfzve
QsFxab1be1qteAcPkc2+HI+B6uYEbDBGYT5ORbyEFshR89pRjMFljmabmUCudn4AA6OEAse4lw+8
MdJcmxtkjM8UDITpzdnfEztqV+1xT86zCYaaqmq8Jde3ZidMDbvhUUS40TxjnRT0Z9k3FUCXMgMr
roeeFBVvHjI/bTW5x0V3WWRLCoAyLeoEuakUILEnEuXCjG4K9Dmn4OT4OQS2OKD/mFacI9HS+PnF
4sxaoGTXfOVSrSI7OaNl+6V+rKVITcwpYnwhlSLvPOCNPlqmM0hd9V0LqdHNkVjFKA+/1cmR8GPC
miKbbSvin5h4FSJwx15NTwS4iKm3EBuiWYKoLZE8IZWCC9hmm5mC2znaSH+A6LfX79SdK2r4E3rj
kFkSvRylA3D63QI42cDijbTRxLpZmtsJw2YoyV3tKpCuAtuk1qJHUqAxCJgmDlwSqXdFDG4/1o/3
+YQy7tZmC0QY+EYII/HdXoznuhuBX3Yt3BedgpXWj6SHflgwVj7e8t/sNHdx2WbCnExGJj7prlO4
7kpdaPD+hNH9t9ZGczT9tAL5QI/yvQDIYU4NYAasnUCA8T3bkE082VJa95gAM1ZwQWN87cy8WEOK
JurR5Yg75V83gEPC8AXEpXJekNwPgphZqrE2jBhKT2CyEPe17n90Pz4ga+6lT6+hW0eXA5tjUAd2
nlE75TWEzwhtbyJrGNw3QPAFTKKb3rbPaM4tqUrkh6ETUNC4k/0Cuo3XlERitnUhph9QRs3z/0KZ
rvfqVABhRF6KBTdRPXABT9wTvcbbNAZdDXKUxy2I+wjPCr6Tkj98ZR/xeWo/YGhDfXraVgSaCfd8
+W7xHKo4LU9lhRFQN12oonUS1xvFciFOTWybrnrv9u+qj1e3ZdhpnEOS2VVVVfsxNSCyuybkvjBd
ajSa3ybGLv1e/4DM7uw+HWiQGSMxg6KrmFujbuHj7x3w26fEmFcZyN9a14vgCwSBnP2UqIb8WYzD
I6UNfI8/YUM+NvI+jIDu4iCLmxjeulFtousZ7S2khCKny3ONmeFPjQcIWT8UeZAgjiUc4aF6LD99
Zblqm9pA47Ffen1VtVfeH2zSfbOddgjB9eVUkVgPdQF4iP9c0/qOZWBv4sd3FZzIfhBS0mk8+X9p
oVBY2hMkW5QlgVR4xM3JUA1Kh+b92xObxK5KOS5utbNCvhrnYoPK9Q1bjIbb4w3UkIsv44naWj79
uqlJZ1l+Bs3pJpimNrlxFhqy1ujsW/WoITHfhcI++tgWrjxykuG85gRM0tKej0OP10UG5LAS8stL
mSah34prZfIpAjHBG0MbVRS+xhtYdo2xjJ5Dq0nVLqluKem3YEjQnkYGXn8+Ok9pr3Y/91iJfJQc
Wjqo+KfzDyN8/SQHItinybhO8U80bpda5hKGIT0aGo/7Lr7Fym7ACVX0PcpjPrgGVpKic0FVBNwG
Y2ROAniRk804bU7xCTdpfP/eeVwHO5na3PXGl9vRgIxgg0pUEZ8sWvLghUTGzBbP8D22Tn3JOAwz
xEhgJIKoMnpmIRNgfsQjJ1P3aXw2PlEtLUDSnKtFWIrmM9IONVH4WMroITWtCIn1wq7HTeX5ivi6
Rn7p359LIHUFLdIuCdvtYBipoNNQLKYWqKHcEK8eH0j6WIo8DK0SVmpa+H4pqETwx350ZU91/Vfb
yyOjhDPURNa4g2c8L0K4GOg+pyJHKrNrpvy+6hq+wT2grcgzr2+3jTRT/lsYmE+c+abZqLnn9v+c
zFRczfWq96R5wwRiX6cZ8trPGhdbbPpKL8ScaxUJpSadlpDXH/gFL/CJiNQg6gDZZEW7hcaDVNrG
8MsRF0oFg5+cDTWG6MXuR37Zj0jxfPcj1M9rZ+5P5mIsSY9cFTDVgicp/hm182jWRRTccyFN8fEE
Zw2qVZMQT5zjJu+C+UeDRLrvTmqY5Bim8zGMeTQOE86fwD6i0QA4avGZ5uC06KSEGkml3GGN047k
0aS4GNCZmwp0coE9n1MZsr7kC/c2nt8fGBgsmWiRIybvHSg6pZwwZ1D8IhMDzAInDvfaQRw1CSc0
uT0R+b5Ikh3gq1de3bk8gxI5uhVOzJQer/0DhC+1l9s9+jXbueVYIqsc5EuqLMpC0B+1udCZn6CD
xfQGoQYb9P+/MLXjgg0cpOnzgQkcllqPrD+EHoIOv7bakqFfyqcYQGu3COX3Hs+msdmH0VR3LGRK
2z9Tbq+OWGGAzOoGI+6CzYp1Qy7Rt2oNQ16dHssVTvAHIqdr0XBzSUZES0GbDbwSVJwDKHYd3cdv
MKArDU3pETYyJaBTn6z1DNoODaXjQ8QkT0vUaGordpK4cN50avZti9caTiLk6zAOE/qkbLpknq2B
bllHSf0ddtfe3E5TzskQ3IWXcOPoxgJA/prLRCLxNcdmafgHyTz9UuNI2iYGdm/M18BwZAZIkAPC
XIBY9rtG0Pw+1MNCqL1ri43lSTrwRzVFjp46lpQg+JsgOMIoqERmCFUATw31A0WKcflrrIyvdfP8
Qafhf1hpBWlnS+x1wMTognkDcdQ39wHI0x6ibZCYDbHzqifhBW8Fqqjv4E+VvZFsWJJIYJytiFG1
yt9hVbVKzY8dpZwg4Fto3UZXJHoVlJYja5YfWHV7EkvUeDLvGUl8k9TMbMU6/jgWMWCNn97ZlyVG
bz4f9AobwPWnZWwGDeTBTjROES2JIV9RuTlRPYI2iD2a6zdyxpDVYgOBrys7eZgjRcDlNKFZzgn6
zXK7a1iVDnAlKBuP5xiwwvzatBE0l/srXrjGNwmwZnuuVQo6su+YA2CcXSg2QPqzPX3nxqUj8eRF
jsMrmB52OqfXhv+dahRNgAkp1+j0Rl/sfyCYwnd3GvayJQBjVw8SuV2daI/Mrto4lhon0NHGGV0y
+VIcvdZs/HNs76Rm3lRU4/xFfSBQvgfdsOabcGVblR1mYTUQT2CDHgNE99t4LAcrJ+dqgyRperru
eRGGXuZkKtfz31vP/w2kXd8IRZumU6spHtL2QTh5IPkFQR51rFnEyeJmC3tO4NjR876JT+7UqIRY
sMlxQo2S7X/GXGqgkwo+oHU22ZQX7bAixIDKFYpbA+YUQWes65j4LAlcuVDzncT2znU6er0xZKpb
j24SpVSLEsFnaSSJXyfYgDVuyYAM8UYEJUJLcy5f1xGtpXMq8QAvuWhOXNKgEoa6N23EF37YLfsr
FFvryfONRKV8NwwQq9DuTB04dGP1MdE8aB7JT8IWkPNRtZT3byOENT25J1uy8m57s5Kuc6cUmxIJ
rbvjEGciHKC9TtqGMctlm3vMuPnYDuHHG1ANInKgPEfa15/KfBuZ4R9u2H3h7UER70FIopF1jZCN
kySOt5XN0yXhkjmRAjzVjNIgtwmEui1PIf/UddFCpRkqHzHiwJ+nXe1lRD6slf3yvRIrJkUVls2F
OASgMk2v3lebXj4XLic40YeedXrW68tlTRhBTLlP9jzIB2yCNMMbqaXhJrn9gSKhWox/rNXM6Nh8
Rdy3TZdsUV6LycQU1IDwA8wR5EE7aC5JddmHN4eJqiSN3s0xdmN8QKXAGZxemg7WKcSBKldh6ujy
I8hMVYUX1g30Ojq50SyjBNQJT12OeFmo9evlR77hoz8c3l3YAQmH3DHcTVkNh2bdbgbpB42t8JHf
crZq9eAKUFrdkAu3Erv+3A/25rzOLqy1DuyCa0qc6hm30+WxRTpjXLpoG2w5q9BMYdIAbSxFLzvr
txZHZdHLXMt3gx2/Ldms+xXHxOhRNLysOB5ofnbcRviwqwg8iOYr6ESVSwuT57Q8uV2ZELVZm9aH
Btvfn/ZqihoqB5gvnSznleYnwux0lWYBYhp6VBFZQ3stISPr1XYJoFBLKqK6mgqbnlDuwjeqdROV
AzQQnT6SL+BKEbqGQUHm90tR+GkaKx9Wsi4vu7juGklMj1INCLhlRBR/4PNkvljQSrtjrkhoZc2N
MmPvh+3DumXTcuCPoN8weXOIshwweo7iOpG4EkCgOaM+HIl8EQKjE3EQZcXi1q7pQrFZ51LcOLvo
0Jr08ERo7QLswcFZYgQGZaIlgqDQ3jyVoOLIyVO27GOELSWAWhciCWrGkK6JocqYF7HGjcZmOrR/
sEbgE3FNOcpbID9Thkrm/SBlhhqK0UoS/taYo7fQHnnKQubcAN1K4i7sL9dz/tCQJmcGBISzTbz1
LHW5TGMZ3/BKK4M1Z9xdRl3gWDw45YyfTGVm/2y+aKY14b6pmfesJCr2cbHlxa9jIN3Qwtnmhnk8
uBtTZ4SZCfl2q6o4aFE5QUjngWFzMsNP/juVNj3smi43xIl4KMKYVS2NtpK/jIwLD1JIph5FhG+1
pIUF4pWCUUC/2skAykUbLMsuF0WaR2pzDGZIHsWN+mtxNNGbBckulmZRFMw9Q5RvdgymkmsHwKUj
rlSHugpSxAoWyvaIFazxQwMGnbsgYMw4ENjyPhNJqhFVr4KVZacmolh6uAJ5hDGMro5s6wY5Owmj
Qv7+/2HZp04Z0FnplIIkaXzHjlqJozTErG0QXP0+M30WxQ9V/e+PNRqId9ToVAXc+x7TnLfscE7w
3bH66MaJ090MzWgPCy1uVcfTyA698BaCla9GrSHTkgpk/wBZYJDorX4aRaGKO1MA1RcVh1QPnxoQ
dkmm/D1i983uvZbaP6a0GUzqQiE2rsj+jFnjzNlGOpPHOHS92I18wsSyftHvYMqXTmefbh0KP4BP
25JE9GoijwmRbA+Dd/0AGxjxsZXvD31p51Y3r05kLMdkjgk8U5T/7Uiuturf1RVIlWOj/uFd66SE
MAty8QIEloF81CYzsBO9WHsvrZuMBfmVj2bejmCIwtTKhTTBA8jVfOO5H/QJI/Omj/wOHpvYkiCy
zltZ5UDiZc3K7I1MLE8o8WqUp5wU65EBUpDv4F3eGALkPhdfzXOd4tLrFZxQDiO9RBnDwIrY3J31
/16JPBzljFU1LebO3Iob4PmMhfMnE/gmMsHFRdilBiTOEbK08LfB2nFwdLESEdUgwwPJddm4zD81
K6uw+eS8nA9b7Np5WQ2d4o2F+I55nPIT6zHP9lWnoTB7oeVRxTfay0PwDMdC22zG1QSkqfzI7b9i
iU7lNFACknSqeuf5+FMnicegTbh4C0Y1YgLMqoaW5xcHdwUt1Bg7kdXUQF6UHj/2KNIrW0lWbbo7
ImOPVWPFYECOCJa9V2bTesd4l01qe3klN593qb9qclTbNMrd4+qa8VqYSPWTXju0IRl/ZD456Xv3
QtakKETSLgXluAQGtY6aYMovt9lD4qPN/K22Xp8V2H7f5Nj3c1ntE4vYvvquiIh7YLBIs2KHePD3
9N0cEMI5Lx7gT/PNrDAF0jMo5qJYFDwEvEvwJkYpATd67w3pMRR5b2ZOfvGeqaD1tJD8GFDTicKt
1/jo3Ukfh8/vzzrU8DGy8F2SUpdapenUEJCOfveC7u18I+pRreb22nZ3XRB47d/oOuInBLeDzN+/
NXGAFnRhslLhta8LITkgJqbHpFfmmFr29OuZ9rlX8kcF9hS1qxFUS7Lvv0MY1FzOaR7JMw05wYwS
Mei/knjQZQhj28VIfJ7zvOehQhSG4n8nAwlULRXSni706DAv2dXMWjjuXqTJDH3E/EWWbHFFysf1
8yFROu6oiJFWOTEeoMhZQN5XKHDRWp16yP2WkBLfkeadOK0UEKuDGu+kuE+lDEjfh1noTXmh4Ed3
fVjlMoM0mI7w2pmyvG8srmRGUMW/ya7RXOHStvFq7u4blvZovlEbNEKR5yPUyM91blQllEnBWY7D
Mti1FKbwfuZzyHvQ5pNRRMwMBD+7Iz/V7r6uppReqojtBBRs9p8ABJviK5/vLA8zGNwlZtxmwfUk
IWBypN59FzjX5dJJ3Qj8NSNQDFWhfpq9GRINFV8BKIieywpAqkELBlSferDlMl/c+dohC7h+K9Pr
QDhwT+Kh2j7jpM312d00Luh36ZSPOFPE6xqv6VniLBrvDx1tNFsJwVKEdEhupGAJMTB/M8+w1Il+
5zCceK6towRwg8nEom9xQgrFq/fnCflI/vT0nJyn5i6laazPTxRou1b8PPfDCE+d0hpVVOzO1nNn
TlLxI1Ij8i1ZaO4z0sThtZjuBlN7YSZVpaFRweW8HcfQvxstUj4N6/KSlF6vpZ3xRGWfnhl0FGm/
/kq2ia5yFmTXPRhIvjueej3mZdq+Tf3ualXjBEQQEf1uLXyuqH2bp70MNtdB8mbfbzqsFM1qKenu
CVgnhlCxiS4h9nT/md6eX8ICFs/si/AnXZ1GDv+duJXyB46fXyTg0VOIxZLR4mpYJDYDTZ7bYldM
jHl6kW5qg/z8F2YDMw65eW+DQ+4DheVHWOy7xYG37nPocr9imD0cyYYdpW1pjnvB/cUHKhqNPHXV
rqdeI4tr46DGn5iEtysQh6uy50h6jZpybh9I2u6mWacFgVKgJt9MAjfuDW7geJl0EGyQCdgRjOmF
61Uvcfk19uT9XLd1rz9I8to/FWWFRJ55IFPjk5RrgvQdena9N2uipj7JyPgeBJFMYClGgcuBJB+k
iY4647p/maZowhYm64jxaipgpv4T2LtNAVkVKU8H00P2Y1VSbRmRpLJn+zlg9kY6uOYZrK1Li4U1
7GkR888C29MVjVqxQuID3BkP2k2gT5iE/T9PYcDcJg/GVLZLnCIysndHaLk61d6bWvqFWBtDsri/
AMZTwUay7o5mkM8Xng8XAncifpvyU+xbx/182laaen8hV2tkg9TdDaG0Pk/SMph9wc8UQWgqJ7V2
GQnVvFRImzb22uNIsLh9gPbW6OTGB2Dr5evApXFJF21vO0f08nqgVCtn8sgBNi8NfPGMuLZhGhIc
QRUQwViiA4F+QRp2GcZLevy9D1SMXu0EUslwwm8BECEA7Tz/ezZL/9Ly2oVENX4OR4+f5QzZ3GlW
WGbip6ci1ZK821lSrFa8P9HyzQtly7d8Y22ihzcnIS6iuO0sUxv60E62Ntbst+3PwoopjGFslgB5
JvgO+P1wVwBVlCAOvJcX3DqIroE0vQVWxJbnMJ59beVEYl3CHL23vi3nanMYI1HAZ//HkrI1u46/
ox1V9dHma34W+dj7MbnoJ89hCV1zLk2uw4v5GN+Vz0igtz0qKNBgAsO3WA/GuwExQBQmM070LEe2
Bc3bbgvTyoIq02y3UaOSzXESiBxagdk2TISAR9j153jsBph6SYhTDfxtI+pzo77AY+vqRpGymoBe
b9x36bLTMeMV6dtPFx0taxxMOUlQUhmRaVfXx8wr/a6R2NE9fuUzidEB4SD5bIpueIhd8Db8SKhU
QQPG5YDJUzAwockRUuxI7EsJpwwWDpZzbza6qqmstpVnqysiCVjylaNdLaJcaZQmHSxQCpVuNxpz
A3ckll1TKPoOLO27CnfrVKK8UJYJlZbzY+HkV93iOk0buv0pVP6EdV16GJTuPplHYqR7SEzfsIfU
/WgG26Ar6J1BF6B9JLqn94wUgypxyjN3EZ1KLlbxBOS1mrZJz9Hd7HWBxcHv5/B/h58/DEFVGFpn
cAeDAqAv4tV9ZfEtMv/UoLKG2MOePLa3nmw+PHv3xRSpRpjHRPWVLNrazJ70wj1TgHP209T773h5
Y78tqPri+tonb7Q1Br+iw6nlYcJNbIgEULUXig+h6JO6RQ9TJOFwTxB3ksQRh49Zk3BbCgGKkFO/
YM3TSejP+2AU7jkLIoGokqtB3UMmt3fAtKBQ8rGRQq/FunvHRbZVvB+SBtMumzK31AKU7Hz4bjiV
Ys4XgnAIZK+coEJFqhx85jjvfsdkK+CTvP8UdlCRu6PGRpCb6krvwoZUw3Uz9O9XACkNaOweLbos
U6CpCErQcqCPtdRmJH1IDfQgrQ8FA9AWDvOvMGd+SRpWrNc0IprUdPLbEYvBv8eWckgamUA+dHbv
sVMWqEeRWOyEV+eXXbi2pEGgSDpiQ6jGtYBzJ1FMi7F+67I0JIP30Rd0fJqkbJ1whjjDG4Kivp3P
iQCp2UaU7P/gBUqiA65S28zNgy/jRwfZjCMFOoy4ijg+reseYqWgWuknH1FYF9XS9TSB+RvFasJC
FSk6pis4Y1LaccFe0V4UF7mPzPxpH+l9snGx8lA/Vy6TSiXlEBFc6VGMR0dDn0TSe/519Qze7vMm
0mTtpvj8ItejWk8XOwoxaZADOnY3Jbmxms6QIfAKmis9J/cXD3DxTAGSLvGb5vfPk2LR+6vG/s+H
aetxgYwyH/BZgvtgq20UfmIh+rJs9PqgoJB1aYlxOwjUtpoICCUkTL1fje50RRovWqIQOS7kiE5r
4r5HkXH+9ryLca6P7yXArMp2yfW5KZko6yU+xCCjTEK9B9x7l8yf0fUNn1hK00lvIM+NbvF1HeXU
P5gG/dUF2khN16aZX7sfQ3epWuN8jSstIryZr9d/woBjTGYXLN0NUaziEQaBwZauV7hvOWVeQLlJ
rkedYHQCpCt0H9waGIp/YVTYuvgiTpcQurjAy6B9zVa6hcgO9jWSADwwDQ5YDBLBQDzy8xO1eD+E
iyaS3Rg4T+YIhGD1L/6Bjf95eINayq9c6x0LYEGhnldA86wMyDBjDCVWpoWGJzEWTzINz5kWwf9K
1s7ANNK5V1xd8lZIZlZRH0glMuyLMG3xTMGDuDw4wZLYpwsiPJqkoUHJy+qklR2lrAcczFqiiptR
o22Vhf5h5GRzes74tPt0cZVgEONvGxHZycpge4UAq7jC9qtxruNDe5ashYhzd1v6WfUshtBsP05Y
/l1ntA3CVqDkas3PrA20jZpJ3bceDKN5sBUuhUGJZZX84H8Ms59NrdfEGU0hDz/W4gAMc07w7UDT
XIX1rDvoECeR5Da2wAT2alLKi6sJcnV1f3AvqAtR19yxhAwt3fMgCx7ih+dz7Ijk5Mgal9Jewfps
p10pnUWPtm1rxKKAFACjtO52WaNQV4z19mjzLTNLVozbE0A61vg6CdDaQjaATFQiy3vogHftbgIL
YM/VjfCx9L5i9ShT5KKDv0ltXU2mC4AyOrBPqdPkS0FEUZbmrumGlXmIgOz9bGaf89LO0gNxRZsd
ccUtYc8lP2sGtG4nhkbp0p2zueUqI9YsB3xS5RGOZ0b7/5rPX0UrHcUr6411WQJ3uGLcq3/5+Jb5
xIcODZdxKQbWaM8Hes/uHu5IcPLMhdqUc0TdOJauNKacEVvOb2jZFuxnr3bk2MkS63H3LC0TmtqH
w1MvhN4SWyYNYMOP4OwMAjrxtQkXOjstwj417HW5kJXl9t7oUTDvZeHQ7B0R8fncKqyVbGV6FLcQ
r4OteJgDFS7kKg49pxqRIaPiM1iuCMdf2cswfeKrKAgSzlAcj7QE8SqpI3jCH9tguEyjpkATRkaD
zuSNFihvs8/5VV5heokAN+F+HKsXWxu6kK8dqCU+CcPPHiZdObWs5upHr4gr7PMR7hdCWLOt5Ifm
bp7qcjlpUP0eratRyORbjiTYtAohzkaS56WrD+Q+aGrVjj7anMZ77NpQy3wzxstl1EoTYNXz3inr
jh4o63PHXWAGV2m5Yl6Zwr+T6JFxF9ROxswLTG6fWdPIelO81QGnu3w14nNh+yi/yS8pg5YTyZcT
QErQU+GOD2hjjUdjVTRlT+ZiOs0OBQy0nKO1E1unsiUSjR1ZIM+lMOoRyQcUhCDTN4HdPUKgmDj5
T0rUAUFT0Ljv7hXdaTwQtaSRLFegGP7oYCFsWmC+lrV3770HU9sV3uiH8KbnVaL2OjYTf1HTGwWD
lTnxURUR+yCW+LYUBWotrpGj1R1odNfy4PmwZVCnp8b/Aj6vOSsoxjy0rqx5JaJWGvNG5KDJcuTx
+aE68R5jI8SM1ZGBFGu8j2zK3fIKsahaMMpITHsr4sJqwrqGflpzLcGeDbwsXjYwDJ1lRwY9Bcdt
9mSLpMpqvmBqm9GaUp7Xqcz2AsDUBLJCX6m9r9O1u1ZMnSKgV+5uOaCzNTRMzUZU/9MIcyjs+Dvq
FupHT2Lq7GeP+pEzN5JmqKJpN96t6Ei51TOJPZn0+XM1KiSFtPAMLQN4LijwQKILIA5L5EEkTuge
RjAd6E80v8jvIT4fA17FigaYTrnIKPxQB8h9ECVGfw+IQG5nefyWOtj66UmSeCu8ypjDVZKvPzzI
PfBMVjO0Bn1tXrffYyCZ/FKAeQ4V4D8gLuWrxolsVRxZmBBB7OW8CJBoG03kU69YRLu0ltWLzlej
6gQF4bNy3k9kmbpXl0hGC8AawR5L+TtqpGvdc071ytA5dF6M4rRw039kK5BfDKVnmfsJKg83R293
hDzYV0PiVVx8SOumPGH2Ui7kQ6kcYA72FIPF7H1Nwqo725U7z8d5znqdjFPZtkyJ5Ir1hGn7Sh1d
oEeY5Y/GMtqYvD9y21LwaiFHoHe+oToXD3bJOIOasDuYvsYCUCtjt5LVNYJitmVVFdtNc6KjX1gi
cfzIA9/KttlepsBAhXq4NZAHkWpqWowqCI1lfmy9zHHMW5WFPVnj7nRBFoXA2KwNFihbEmw7iBGp
GpPAOh3GfnIRaglN8uJcaxQoYysBxkcndUSumrPrnmbCyvjVmptinBLRjgnebP2fI0fuzKVjphQE
KvyxEByGQj9yq8TJl7st3QGyrRT9GnSPM1bwg99PzDiN6DdpbKS5BUxO118PlwuRsaPkbeHFdJoO
Dp4LJ6xTe1JCWr7IN7D94jY+XJIvt5v72tYf3xmCEMZkiSwMujuB4tDFgn0bULk+dWxByv3WCX/V
VPx/UviSUwzFrpjS18Q1HaLqfKB7mB2/zUokhfb+TrAWsgAQVXZ6U4VwOs01W3Xl3vYkhdixtNC2
CiJBTwP2OzwP5+gHgF54YemA8tvb+VLNJ4fdDqKXDaJvhiN+2lYMt3ugTKkrd55tzBE8xjJQJcT+
LWCE6B0ePLDTILSt+2T9uxkJNDTVvLMvECcyUE8Ll0tTzKm6tBhk2qP4LaxoFgCa14G3dQGDFDgh
DgCK6R0zWnscHn0yebiQOdRk2wYfCHNBxeHoiNOZ6ti4ddddx8hVYF4MPTq0c/gdJiw2KiMFqdRG
iwLSFqvf9wnZZjMtZwUGRG/RQE2Xw+In7zlFNQOrdfTqMYVM/Pz+qLHk/OyQp1rdd8a87A+F8ygv
dOfHM+sD0nRDD6Pg09sb/zyfRytv8WXuI31HA97Mh+UqQeAyMTyJgLwPJaF7+RQ4kP322+ojLfLA
EGxQSKiHLI29XO12FY6w7iLDBdjsCSP4XnA4L8Bsx3/88gEZc/neqFHnSEBe9cGJl5FmvIabk8sK
AjjcPGNRbxwObeG/7Uz/T/6Hhh7uF4zkmW3pF29lMmGooIyee0SY67vKdgB3UycVnRtTvDQwnmpb
yzeghS/Z1SVOO4amluuXaKAvtdJzrVqF0ITYTJc01TEh2HKJFUKnusGJovphTqigrUvSVyNNBTsG
qKhinBcbuCcsnKSZmBhL2iB4yBVlX2ybdDhJSXy5Orti3bTKy8s9uuob9R/8bbGuaTOgIpEFGAH2
ej+ea5lkgkfgK84HzBF7o9CZa1Hwl9bxSTAEdVVDhc1RPDoBBFgTtljvVqCutdLN+Thb/dGZ41Ce
vGnxkEX7htvG9aCRxf1mD2C7Q7pIkiTr7JzQ/x7V5vssu6Jtw/ehwxGSmbxpgDGZmzWeoUpWfuZx
qbkaB9+4TBRAsZAGdfZkgh13PDeR/LHo3e7eVQHPuBAvDGZ3Eb4i7aq4yOavzyqpXbKd4vRWxkOn
0KAMQ3jS48o5YxyIPzZqZTvWSl5YInBFUeBmRLhc84lIyeuaBH2iDdiE7pu8mBjy0IV/68CGvDwg
KT+2oFCNo3vAsK4zsCT6g3n/y1vTpJI08RszHZWGLYlnRE3sjhhjBmqR6uqjKJuVpXk4hnhin0/J
E687+C8zFJjyLh6wPKBmtI/umqoKA0AtiZ6xUumNMOF5MCErQ6qn8cGkaDkxzIVsI6uo7tXkmudY
vsoRCPkSyXIZ1HQiOYwnNcAW2jNU+/FJq0Oi8i93gu/Jyxb18G9apPce/nbH5TQ5hYQbgHF33FdG
ikiWlCySnOsezfj/+/wnKPE3rQLb0rsRs4B08tiqgRC7DlZvUksl1adB9e2Hky2g6a3tqAt0iP4o
dPSGFrqjSN9/woBiPtGpSsScsNa8uEvqLbxzv7XX/er6t9svNCcK4esWRej1ouQVWYznHsVFApgA
+CG5xT4If1ExSBbM2kRNbwr7pWhV8TFhy/QxcNEB+ar/xDbRmp/ieV9sep7PkIbePzh5wY/R4OPu
lASKfPXonCD4tl3YD0YVr0vadjsavSfZcxhJrsIMeZyQZ6mnR/7kNYXbsYRm1Q45GHQXgMls7Ubq
WilE+PYhMXCxu/wYLRYjA+NlfU+vjX+diNU/YYB3pgRyGDVWPJvF11uhf5l6OAlXYFxMtNVnnwWB
6des74H5F9nGsSZr1qw6hpiJGhGcY78TWMblZU2Hb1c9xy5w/CeeTkXBVf+Ag3WVqwD5AdwN5n4O
NEMwLvoQocOS+H78yWDfjVNKWj5VqsO3LfOSenizL+PwTgzcRL8I1CgpZJaSLUKlVupQDZtgkPuz
U2WxKvp8REZI0TBlElvOdKz1MxnSKXFvg7/Gm7AzyvBATIPDM98rrJu9uFKpc7ahg6ZqRKFdsB65
a8kwD28m80PO0kx3wDlqpHbcnDUEc/snTe8ZbkOjJ+DM1O7JZgyJd1RGzbHFU3+kgmfgl28zJuSH
y9c59DLwn1/ersLi3QcW8Hgwo4/8vsjk0hNB3k9dyFZchiQLBmPXnVFXZo67W3YIZCVhTFFIDT3/
Y7DWeQgK4JjyYfQ7lThBquO1QGl5v0sCJ85ckGeE8tvrH8F1bf8iflvd4eUBEziKY5ecvw8gJtei
NKy+4hWUsJhRZtFQbIxmrreYYXmwoQLGHjzcYqguFGOXV8A/8wg7+GOFAZk/a+pv3QmJF/4lmh5r
U7/g9FXpeiLtYbxcrXWbm7RiNfDOJ0mM3ewIZe6qJtM4DiLta+HK5UOwkMnIKr3qn6E4Lp4UDeVr
inMyiwkDFZlPqhuqdG6cf5EOsQlKuYnZjFrlvhJ6N1fJE3MNH5ThjXu/p+GiftSs+AL7qRV+uquh
L6cRDOfjZBGsmEL4uVIS+hEBpBbfap6iAlm8aW6buYl8tI68dJry5GXMbJHxJ7TKj5su+Tym4ocP
fRDikBRWdl1DpQHFj5nIe99nEf5I7iB/F0+6OLbuowVl/7bJH8kgXlHwTW2fFvFsvNk7KceKEYfu
9lXBPw80qcHq0C4/hE8sD/cLmdMyP4d6/8305J9zl4T4M5runb0hyLjJ6j19PYlTVJNMB0aYN5+W
8b8HnQ0ob0XMK3CwlqOwYou46XO+k+nyT7MOTcSOPrWsLx8uc73w+EG/9G4kcT2GdwqKx89rUxRD
XV2SeGhT+17S9SuPd5IYfcYDkJywd5F3VFkc1EG/ZsyArjfpRJA4urWIrAMXUGrHM4tMw8HlZFkz
wCTUlerM2uLeFmOsF+h5phFEXV6MedJuu/krINCa1s4QB+vuqQiiDSgbbGBlcKF8VZMupOxmUCvE
7OldioJopwbcP5q0KGQlj+suimOIlS0DABq4RjlHghfR9qsNCPdyx8ThYtGCy+h82JQ+AUAXVbC0
+Q2d27nt8hcZGHG5GXBVEwCSe7eoX8yEu3FhzFT7e0NWjpYP9UlRBW3hzGD8+JS5iTbezq8PY0Cd
3h1bSYlQZ+5iyQFHQBRKVaFtRRLV0w9IHyCYNN6JYaa9SxZ7vPf7ObP804Uyx2n8VZQMW6YB7cgv
zYulRTLAbtSgSYU1zNTxfavQfmmpnymd1Vx7dO5JjzGOX/CWJFzRoGcrQNosHkhj11fSButbYZgR
3jBJWWH8YYHCbH3PNSgCXiHsbz6NsCx4o2nf/HGPs53PiPyUocIF8/qap3vAZ43s6276kxegsO5z
Ws7RMh5KU5RA/Bl652DSDOhM5GjCvdFoyxJOOzzw7j31gjAOJ5StiYXVWo00qheqmiRRkwxW43hM
v68OqesuQTM9p1Dzu5Pdlc1DJm661PcAJI9JG5Ab1MY1dfSZkQ6D8wArjP9ZNcLTIA0e83To1zXI
L2ClejjbJ+G1tHd0WqDDRe85eQyxZCIBxSq5n217+1MvTTqnmNuettdsFyItJkB3r39Ob4772Dfm
+nSYYzj++gdwR/XTaNi0zdRET1jnLSFLdvYwr8yCwbIpm0/i4oeaRzPuqRjj9XCXKMFLEIyD4YhE
YlsSfc/AW1nvMf+ZRbdrsll4gBorIAMfJBySLdZaXcpeGeXTmoLOxKWpnFWyHH3Uj/M908PjIQmZ
VB0imiZ1+Nn2CR+lLQ3d/aFs+VvEhmpCl/oWIWwBJ+xRIMqO2UM4D3lV7CbgnRUcog+SBGjnLTtF
tb6oh6n/VGzMqPzdxPVMc+JN14p4AgvZxlkM0PcwDUyFwFQSy1Cgo6h1LGQd0UGAzUOwS0H+wEdS
TXjkKXeowarh0KXj0SCMQZeMNjj5uMwIrKUpq38bDq8CDUrRA2j1w5vN5jLEKZbMW+dISKZdbEJa
ngt2PUZVZNA+9l9+ZXNhrpeQ9ns/IGxcU0Fv3e8JRayq1MpPBllWEIxQez+Ru8f07XKrTHG1EGYX
xidUkd5V2PqyeqR71BMdNvfx243oAKDiBCsIm92VQ0PHK7kZH7Ev/m+O4d30ga+0z+2yaClBEmxK
dkM8bnvYAM6cgoHzDFjMsFlMA4EGQ6QSgNSKJ3GWtiILylOwaYYUhMxPDNmaY8fJatIKJfRcn4Pi
5pdDO/OktUdecda1q1BrUevHqXfdt1KHHhMVIvk0ErFxvcVJOByQ7pyXJbtnHSSy705wLoQP8XdP
cjLwvSuvoPGGrOUjYo+CJjOJ8S8BQi8prLjBnKyAmVk3zxzTzwyjjOJDnXQBU/8sYw/Kh+DOhLra
iJq074c5gYiYdq0QglG0vD7Nm+gNHN6p9q0YgOAQC6Ky5Wcne7vtOfl+SMxhRVOMFJurLnNZhLKI
f3lAGlq3eNOvPDjIYPuzwnfmlGxVt+SGTw0h7ji99rJ7v/pIeIg7d3m9cn7YaVddvX7eRPH4SwWn
WFdCQYVt/oVRK8CPJ2yxBE8G/SscJcesYsgKnG7/kdI0+2jK4X6pejY0y061EIO4wdjy+R4Qh2T1
2R4z7r7taUY3VwuB20KAFrn6ZQh1jgnlbUpKkV0olpPZlqt3ihUQHtJ8U1Vob5m+EWBskvcr/oor
syqxysJ2pEE9XszTXWUwbPkUQOGDiku77DU7N93bpsZ/F38yHQTTeRZXZwEFdrIPkT3y8iuxhO5m
OA/+3XMefWAE1iv5gyeZdJYb2jNCUmpoJ4Fl/r68zZVl6apLXytbkDiJZTdr9MGpb3vjTUpFunH3
nvYsIL8TGOaMQykP4SISCRxdyuoALotKwRKfJorh9gc1HKJ283gQJIF6FKMJd6ib/3nUCGMKPeDV
nAlUXHBN2c9cg1+NZjlVSekp1ZfgwaPWpK1kUr68TPbRg/Jgm7JkvNP4T6SVUE7j8+5X7aW3GpAz
UtjAeVVMZ6o34+PlU49n5CzHeywMNOmnNgJ3jhyHAK757yJJuepep2YPKvO0E3ZeSny40FIr+AJI
AEag7o3RmUuKFBB94jga4AQfFM2ql1imvTzz47uE9mQyGMZqi8B70XVV5sZe+kmtvRlmMnPQis5P
xUxuziYCmcZ32B9V0gGipuC8Quaw8mcQGR6ZwrVOOOz9AD+x4+OxJeSyN7zP49LbwfCsrtLO5482
ndqDCVmm/VrlAYg01smDWh6Gzi2LEDwg25rF14y5sHizcYgmNpCA5Idwz6fV5BD65aj/SjSZvicB
Bp7gYVLaQtMFPbWa1oytkYupIe4ikKjDeS69lXJuST9agROYEXhOp5L1/f9IuPVpqSbJZBZcPuEv
J6zy205raijCa62I+KhHter42vUed9ihSncWfUK/LbSLRFHGR2pH/DG7Zrpu+gWzI2gaqvLjUOBf
ym93LAyP8m9jzrcukCthcH4Q0aH1ZgJ/jl0whlbM7bfT459YvGTsYDQkOubbOk0fbH64m2l7ZoS2
zp/wAbMG2Bfcd4dotjAwCm1nDhxgEC9nSKXFdks8yNrtaEveqREh5obaNNsLD+HEMw22gUCz3NlB
3ED/9xiglBZCc+mBd5A05xbez1NLPtd7Iukaz54v01z9oMJWNusvsNiUxLspXBEic0E4S5JhuP68
ySz4Ev8pnVFaLPLl6u+uwrtIlfMOMNWSJnrjmYJwWfdjCY3xwoQbw66KEFD/XNWaGX7+EL4HZ2IB
Mz0KQd9hUqUQ9EmJE5C7OCNsCbOWlElTsFQ3sxkwyzFHelhkrRXJ0aqr5z3FShxIhOculfaOkt08
288poQ5gL32bGRNv/9ScYJBLUCysIb+rPSpoTRgk9lXQg8cibUakhsBm43c/vG7dp9LWJUTvsqfq
Cq/G7xKaLoYi0vscyhLbrXQ0wZc5WZmCELW0we14lgb2KUDBGfeybBfObyovMqSvFOx4dIuvEyZ0
qeKLZrZ6crTgZtw3NaHbgCoFIaveDeq1nPyXG/PON5x+kiW/hAjJ3oYXAtXsSANnXm6DE0KVZCy8
Nqd2Nse+Ihj4S0Bts5Zq4ZngNXPUfNPKitvimEuFZg/DmVbyjIloPeoeD7222nY8MoSZThcc88m+
kd5Mqvn8LqZ46FK7UhuxzGdAiqr1n/VUe7iBNian8dTOcfYygQLnRBlUPenj2VfDaU37lF7AQFck
1JJrJlgG6oGduy4X7WfVell38dM0l1+UD6+Hmg86r/WHYkew32+aMt1h3E4de/H5ILDfEx/eCCOT
7Tyj9Pij4aF9u22cCtguHKJY6L5PNZLujCw33PTjFKKpg0anJCdypdIUN2uPgISKDeBJiqoCkhHh
OqRW5TZ55hUhv3Oc1hjAkSoKdWD61Oeun0L1yvAFtQ1Hi7NQrBgPn0zNGzmJyWVLpeR6AWaaBJQN
sRRAYQYxiS/ouYbvlFxzfKUr94SHDGfLtCcRpbbbBgWDfzyvXmzGKRtiG3o1DLH+yxadVEIpOPSi
A2DQHSNRu4VxSRO6QvrsKFZS9Mysu4Ck8QHjAwOiALtSApVFiIatCz1peIn86ezYGAzJazxm4qPA
KTKj46bPO/aVfrdWDcHRU3/8O22Q8zTx9lwRmisnvv/5rjwdAT0lEYp5vYf4tdJ8eyoC7MxDJ+7r
CVUyh5kWHZ4GFZZyce4mrf4VwERMOG+djdz+q4DxPXUsbSBbTTN+UUwqRYOALslbDwDK/cZdj/jo
yU4YO/TY32DuDJuJ8nVukORUHWM4kDTfuHvQU7Dpt6ILPFUPuADtOvlKdGuQgD/inoiRe8AB+58d
Gc47wWm2lLH57C+hBV7Ii8SAElz/QqQS1rAxYNxm1/MDJbSmjsxhpmFW3AzOtayGe1CFAJ1pghdr
azged32ukmuX4YJSoGA0Nyce1Rnwsrx/5Cs0H3Ousj2NB7H6Gciz07Hp0dWKoy5bWQLqcJdI/2/T
SkRaCrpYln7KgPaOsKfm73xpnU5zMRhwIWD5NLojRh0u3/6EnKtNR82I4TjDOwtj4/DW2lGO5W3c
+geCtr+h82rLzyzkWIZKK8YaSZhYxODx6CZFwlwDMbvfyWOs+oFDfRLXfq4a/KP/vyMegaTbPCck
hLsvasLKL1XgaLmRX5ZsHA+pSPR11Ak9X/QCWENrkNKBfYtk2BdnyG0v+hlovJPQjwi4gh/hA0jC
BQ+YxRtQcr76UuBwEJGDWQvTCWcHf6A75YQn2goMyWPLAAb1Il04+2mOmbMpXM/MsorcotR3vTwK
n6t0soEk2bHTr0Lq4U3xtSj3/7cSQXZOpQgG/e63qljJHQ8G+CxDscq0TWZE05s9tHjfq33A70t0
YAWys0qBQ2Z1LfFPF6PeDIuOaPV/6C5rvO7Ol5n1hX91BF6ZDeDQ7J+4N3KUsDyer46U68FClvGa
XteyXmRzCvrPYEo6pPPCZeF/oGjL5QQ3/v08boDIdwTe76p6oiXWFxjGJn8CzioakRMXmHFfrmcX
5WEF/7zUkFUzVjt31u3ODxupTzaloECMljsy3Jv2dArhlgLPdIHv/zlLVP4YRWAIXzYkEdjYcOpG
qB+gYfAGgNdujZIsoOYbeht6ouIjQElKgbsWcFtLrxk+hkAHPbS9bUtAvgTnK0sreAq0vfsPC63i
f/gVcuA6yniG/dg/oHs2b5WkieO+xmnH5lB4cjfV//SYOY+5tDv5IxInBEq9gRYHT6IGBxiUbEYb
Zqzg/MiYBe5TV3DTMBCCH/xJibiIWa36ink60LJiv1iCls53dJhh6PISJhmeHB+4SrmOFSAUlm4E
V6FVtqWnVCVGVXy4JID8GzNomeDMsxWccwWPATbWaISwS0ESKjz7USG6maI2SV2wFWfYxB08MKZl
Igsj82/la/TamxeurXo5GSgRdYkWzBtZhBhvc1lxz5jceLFt48beq1AiMoKOhlMRsPUUXin2VBAE
9e41LVkG2FiJQKo+fYxZ+rxICjctno9UgUJFqK7yVNHssmlaA0inuQvdIfApQgYOl+6thJyqnNMV
N/ZJpGe9R29F1IHB1gnD6brgA4sKhml14zHnBZxWqb2k9tETE+VibRDIkjMa6azzs/QjBinQHsv9
rQ4lzQEFMiKEwWp6zRJ75mE0T5X08QBbUPkk9YN3bqjfg5Na/wDjg8yM+akopgedOLCUxUdQoAvm
UgMwvSxvefRn2omYeSZLcDsW0kJKFhCduUAvkzPiKc3XX8n9rtKVQmSXmocTv1oqoqBMLaUChmCH
ObSj1TMODws54wYbArAcHOiYOwEAsvoqR3QbDfNXXEEG2D5Qb1hH1Jxem7VoiJObRqIUV4QqdT5Z
+eJBJ8Kr6Wm7+7AxK5kDi7z+Yr0/uwXa3vzcw/MVLP90VyjSR9QDNn59LSgih5BblTkqDLzI8rab
zxo6dx59Gm4HHWCFuj3CvED/xKLBpwPJ2qqdgl6ld7YcqkoZgffRTq+FUcurLalUc/bmAc7t41K7
qn/Gbq2iAT1qMB5E6EOzSDHNJtIt2t7wHJ32uhS+1/lKTTwusP7GCTG7OgWhRBZlLMNHOAgq0QUO
N0/RC+uXatjJZHV/Us7R59g95g+D2c213LW/lxiq2kykcbUmyVMLQiCVK7NoUDym2Y8IlWEDQVTB
HkQM7hQz0+Bs24ROtqW7ElRLqqIav0r7LrcC33Qg555R1tgwpRVeBGovGkzGW7K0PTw6AG+zrtbZ
EDmd9upWQI9mI5suAkBBCg+/GLWzn3v6E+Xwi3/BB0+kP8cSgLuRYBGCj+w3eAUNz3tv16l8sRe/
d9qjgPUInVpyCskxcEPifU1fp6tIkuPUPuVHr6cUlrO4D8kJpxN1DNAJOrbOlmIL/yRmb7wlpTEv
mPkYS6KybWLGCyARfWOCKclSpjR2odQMUIZd5FkUrtcU/LCz4ASD+qJEZxgjSPtzFkBu4huuOehD
1f+ISf6Zxbm19NaUO2blWQS0VV7T7SET1oniL3yMDDlEBmA1Zax8vVLKc+MKLZmr58uYCG3M49BA
IaqArF0mo8YB6J8GIMR4dWVIxbRAEFl62mqPo/BkkzjudthP8Tbgl01aICWGXhDKE6D7CGrT5+O+
E8E5riuDXZF9KteDEws4tyEk8dKJkvIbPcMPG5IL+fdKAuCfPXfApmR/BYycmJBYO+QrqPDiMmBC
JgdTyzYpySYuo+dUY0TXB/N+RZtYbFxHGhSG7G1GvOsyGB56je65aA975JRRP9kZ1g2j90r+y4n9
nLlbhCu98axr6rV2xa+Sy+5fs3elW6x9cPRK7qFyt3+T5RtCpchNi3I7jH4H52vulMfOsmPPPNw8
xZZLuFfrVoafKM/fAWpjqN64zz3te2BxCUceaZWbDoXqG85o121r+c2tzWXT5v7tGLtNIgpLoB/p
l7G+z+h8mZtucFxu24OxbeMMccZQJx1IWc44pFgoYp+bYxnTmhN6I02V8OTA51SO2caMt90/9MfF
AcB3+9DGFnjV1PuujsvTMRfcAymE58Jbe0/OAc1EESoMzmnDVMNq/bo/VPIiaf/X0FA4KkGmfv4s
zvMs30eBdlCVO3CY6iRExiWJ6Z48QUblNU3bbcbobXJuPbL4qnnBt0r94e03B6b4XTViiEIZLWXn
4yWMLlkG/UmFudaixnPRRKARuuhUO/I9oW/mBZ/SGhc2ZdV5s5nHrZDwjCCAjai0u+sGtS/kP/xa
+CXSHBPqdKL+gKdbeXgo2KQxSBbvpNtx5JD4dAbGZ5gVvdshLTQJwYxJ+xu/hNqQXIbUKc80nqvW
WoLbk2lzf8cErPkf/vOgOiJ5VpN/5MVoyYmQ/E3tNB7IYsfgma1q18cWPaKe1qSeKd9/vXAHfuHR
i6ay+0oB2CxBa6/hYRvBqFm3+ZaKtQwJZThWZk58Dum/PHbZMjSkjQEVrIyBU2hNBaRhhm2AnL8P
x/oOgM/w50j9Oswozq5FooUGxRLN4c8Td7G5AjViKE5y1WfwKlwpgSPFQD7msLBJESgoj3x7N2fw
UmbfA7VD4XBgDB4ZNEVv7eSQDK1XxyeHWBJ0XNQa9wU9JMG9KiZwu09pXjYIOljxoyqx4e4Ptfv5
hakCXFblnUzJJXiBL6MBUZvc7LMKZCbb9WWFjsrJxBSZ5knw6zKIKUeW9B88X1P+MMYZbSx3i7z9
it/gG/gfS1eosmI8FHG54Xa/fk336wzwWNn+95Ql/ZkSpXd7dkbbhPNk/n+Strv8b9uuxInXbDyv
jLe9E7AvCPmmnibjgQZQtWAai8caCIOiRJGXdRuI3S4pTi15RVsG6DZH6MkiXeT4FZu9dmcqtjRh
OP9td2UheoYmxb2OlSMFlQfxqc1aXF+C9jQZjwTdAqno00GMg1R/wRCIAL5oDvGA25FE4ez5pq+k
/UQZqU5qE2x0PFmhf1u7our9vTO9l7GrrLV3u9H6XraI63TnX3oJryTqWD8mZQeJnmbBgAWF/g0d
9SodbT/+O31zFebyTSKuVQWEDM1TVD7SQMo9CJXTNY5CB9+8tCPJ0gQyjEGQ4r3AyaIqT815nqhu
1NxcSV2Pa4kR2qUPoClsGZCLJRFSPMPO6CXaowvRpJEnamg1mHlVFJe3CAbaLDFmzud6Jv1CDl5F
tvYZNPsbXphOi32qWb9j8D2ZtV2PfM1lJUkEmiEOtLNGuk4fIYI9y1QRQC0zBmoe1PIKxmZu/kny
PXKoBtr+3KipLtXdllmoNzMLc1J0CtbAUy8URIgALU6mxFvSuAk6hmaZN0+L7FhdqEZ1Ni/3PQx7
livWEULpLoNJreLTiZJxMbxJWdGFaCpw+fn5f0zUEKJgxYktUjhZzriE6q9vgLCrL6ZhBfQ57sWu
isYRE7zDLcg0yTVttE9uGNboCPhC8P12Y2TAO0h/yXAJ+SKeGXokVP+7iBsaT8m9ajDylY1JEsxp
vhi8AgkQ8g4BCCNW4+Fvxzbyi6WWKgjZqsVlkQ06srYE4DgPInzgtPo8qoD+Qv8dmD6dmHHNDqDi
xG/bsUgkXYzgDTLfp3lrm4Q5IdBR60RBE6QyX0MRFZM/tflcy6TlpSqZIflBdkJ4g4gRdeGKUm7t
bsdT128N+OyZFhTtiS4UpiCz3CIse9FRpNhL1J+2BggtdbFep4MNq9LZJADdeuvhct3lenqMNU2B
YilOjuObXmJbEFqY2ADD6qe7g+3zrEhQ3mVQTIJetFxCZbD31mPbTfvQb4aDXWxJDlqpZIZZHKaW
6wrpEnfduv0ZLvWqUGWD5XjGZ0I/6teVHq9peHgijpNnSzXIOuSnRv90rWLve2D04L76lCuXgXJp
9obqDwVzbV6mazjep2vtzZBLKt6INCJws/CZrQ/NYWSnefk2CVnaVwjkeF5j5kgYaRiBrNcu32gC
+BJJ+FzpPGfWLNUqLGHNQ9CLqSIPypdq7YaQWkZZtni5B1GB+d2X5KLa4H0xxuBMTV9e4DdTu2YB
kC1N9AfnPgoUEpPM7DFKG0uomrmJOdBw7MCjOj4SBAQCq783AawIpouYAUiiLAFjjeYAQQiFNsfE
BhNtDJorebi03FiWhjX69IKvtX75KPCAz830TMICJRf2aIC6DYVcqYke+RjenBHOQA4Yct5F6C2J
XUrFB7L5otSCBOh3SXHx/BTVAPsd26oGSoDaQEzsTs76gK0TLqv+MqGqvhANSoHiD7vICkPSA8Tc
JZAZj4SpGdypUcgOoB7sbMnfiRlQmJTe9KHT5VFaEGANm2Ux5j+uuj5Uq9jc4BDPpJ2/WUVvgyOT
KXnKJMRRr7+zV+tcV1YEHxzOVplYl7uonwkdTfe1VXJfCdWRT0vGCe44x0elJhd5Udth5jzqMhN1
eI3Ub4B/A8gFxacdfGxbo7BVCXDP0b2ntN3Bf2cgQD0dw7WfgayJf9Pn6r5Z2jm7q+JzkcQw3/Q/
83DaXJyuDdUdAcfzHfVDeYQOku92BNYvRvKeNCyjpjfwIs+tJlVB81Wfy2CbcjGSGdQEmdXNyvK8
OK55V96QWMY856YVcIisu3IOG/Hno4pqnhMUDSA/D928XJYgOD+/VkVfgaFZUwwwH8mkgouReJlh
Y786aekg2BxZkWwrKdPvrYrIY7a7OxMHgp0QJ7D/qTY2VWBO0w9XEgHieCMJU+HIZii+OfhERW/g
D2BmGT8Qkl+L1yjm5stwIDRSOaA16rqtZg4RYGMPA7zoNU/IZ+IY4sqp7xoiCNNLyQ/K9cNYYs7H
sfo9WVmriDDQosuNN3ZKCv6XZxuEuh6DKP23bGs5Fu5TjjJRlREm49G1IjldbLtk3TSE1EO1kgPh
keK8RkC4J9h5lHqd3ia1G0te8IwQcPK67xqPExrZR0roflm2La5SwaFqy7mgWK4IQMeHT1WpMjUm
+f4Sud/i7Jl2YS3J8t7yJRBllEeE1xcwcmbGusceDSWffUmMYJibq1zUPpc5W9wLxs4EV1Wk1DNj
zPVaimhNA46tw9mqnZa9iHZKXdbu+Lcikv/rzRypqyNGXwFHqkBdX//wC0mE8D4iHPIRyWfZiXt+
iA+Mn4qUkphB24DggXZ6rkYFsJdwTYYYPpT9tRc7Uz+XrRCzD6E4jyI8Y6+VQlC+itXX9gII+JJ3
b99hRWg/sTlVWSJyUfU1sN1xkWhDmjsv59FOEHi9CHhpWkBtfp0eXlGK0IW4RTSVbKcMVPnzozAZ
erpfRSK+qJhcWGM3OKVPBqyL0x7Q7xFqCLhWJ9x6MeQ4ftWF7+FzvvT6NE2/LYJk5k5kMIsRamwD
ZT5zDm5b0g3VgOG3a2YyuwBMtpkPRkY6rJPv1SFUyMQsdnsTOtpBiusvRyVvq+aly6bzGDVWQfqH
Jutq8ivbTsrHSsgKiNjLLgJJ/J92TQ/RFNmUldGXbG9+l8zDJ21zhpLx/u6ArDfOvRF3vdXlcIH3
OKjORKtSZYg56Ni0NOtgMXWOe3r7kzHaoCLwjbUFvoR0qw0lqiDM1ZHjhbBe8qgZjGpCPbgY6Fa6
WmHvM5ncBdms5KOoCROiQwInrUBDxrUBafJywVGtwYRazYDK9yPKSfscKK2SVKVlavsj84pEmjQP
MHvBe4+ZM9Azm6wknLzxjc510npXLH4UhM9xMwNiytHoz5uNkXeD+4JDiUIbiogru3ABj/WsPasz
ffcJhh0sE8VXHI898NyjhotKtYX3r9xHJlHZiQs2oOstPltwbrIR7a6MhDz+AYgaRUx9YvQO911B
UtyHk+StSyuZ+5Smu6Tn7raV6dP24t6HRPkrqUtCNwfbYWYAXX1ktSbSI4BkulCVxXVis7f+YvHc
4bPo67TgpW8pyd0Mj0Bnk8haCEjgz8+j6apqyB6BEPnaH0rLJW7nKO6A0/yCuVGb2ai2ZNFOwFxd
XuCtaWrRNSqgsithK1ZNVmYwEYyP0i0QB7dAK5upJCZw0aVLNUtrFPo0gBIom6ISEj9nbFSK2gZZ
zpB3Yc10GoGlCAwsiiWsjttKJ9F2wKPnXj2FLFikY0mfbOEUp3202pJ73WkNaACkA+1NWgVoafLU
Xp8bKXCTmoJHeKngU7GuQCOkwUdGvKN+sOjPKjR3RdAzMfOMFieSjIiVaYWi7mhRQ+SRgNIAxCYg
ZdFRMhVhPfXOfCLopt/YPyKUmEKDJUMQHIbabBrNHpMWMfjADnrDipc7h/etwWuCvcvtpH8CN2xg
MU0vK/qji5GT0RvLLgRHzv1OjDVDm8O8NBoCvRPwrhs0DEDSCyXREC/y0+SlFbH3hQ0fRh6zDJak
Oj39ocojhE/+qUlOLvdIbwNR8E3hUZMlY6qjiTe/g54fkpa3ViPGZI/w1Wy8J7cEhyDiowKD1hSn
q1q1fthEjBWw9YJVcsFNsRabH5QfQIK3nCguli4aYv/jUvrsOQP8+UYOtUqKdHTsHqY12fvr7dDl
n4UM4U79VbVqV77t9+6smhLHQOkWPXsmV3OimQHYOUd1ErgF1bWSw4/fsUX7ZdQ5lSMCwCQgY0Gr
EW3Z5eHXjZnZr/nglUNdqo+TwVfWNzCH/vRP+uqhbzClsq+EP+uQN2i8WUSmWF8cBPH8ZEgigJkR
1uwIajpgPvNtCVU89gA28/pIYwKyVjAQ0mdkQUYZ+U5WVRtRetTrtxEuMzV9Gqo44AgiXBoziBHX
UlX4aBCLzhkQMg8a4R4VaMh4OvDxxj4+/2N19b/lgac4iPSAMn0w6RZl+J/Q+e2ikU5zKM/CvNBa
5zDQwsNuZbUHJzHxx+7r+b/N62GhXp3tqxBOi8f5OYlM9tIYBPVmpqR1Y54dqwoUwLwhDYtCPmZV
34rq8YCWZYkkgVaOkVkRfRhwRJttrQ7Lj+S8ZwFEwJuBfCZsq76FMsWXsiIQMR4jVgcS+JFnOmAE
Rz4Mvf2ox9m/sFiiQqUPeNitRJHdHHdiDdkPWwKWgLxY0wg0Izvvh5aCrGjjvUcFb0r6ToY73Td5
yOWIz6C3bPfjLxE2ewSdbyq+gleENMk0CJuZ5tA3TbRnOlB3zKwbhimQp21ajubkJKitUSJOAxXu
q+LOSHZu5/5WzXwYMB7NhTKD5uw5R+b/rPxgG61MLlbAc4wpSGNz+c9JQOkuDlI39Sl3CAyvBRka
g2PNC3GwRD1rj89a31VqE4A/DL/LpFsw5PKuVsSFKbIqXTJlaI1T8jy6m66FCmwq+ynqxtM7g7tU
JNH/UeKUh4N1j4xTjKcqddyOUmQJWcuOT/zifgvfkN9xhPlZrAo8Zg9Q9UmkvbBHpQPV5D6h2JRS
yltR4JrJy2IZD5dBuGwzUptCSfRDl7zF/beiDFutKKa0RF0owh8JZLAHCwG+FhIxHaJnHZwGU50u
JrEWLg1m2E7cFPv6S5SZWpObPjz4TrZu97LjGRNSJOJ6Y6xxpKj7J3zZ0emr5FCQ6cD4tev/WIhi
jCqdJMXOMQx/sAOilPF//wjaYWXoMEPTwJUBXG8+R70zLqi9IPo/jCVQDqMTux47PFsd758NJ3vt
zR/pkMSDn1NEyvr/4UfWFRKdp6fE0w3Gua0icTsamHn5ycCk9Nd9mzaefR2DmyiZqnpMX9UDlCeg
0bw+rhLj24MibuXuCJKd9SHnKijauRwqM00hC2JAPHy6HiqI+rfNpWFbrpQO+yWtTNtckeGJNc5r
mcI4bplklKuOmDuE/18l6GBt+uIds3CgXxg4Iq/Mxl40sE1OR5upyXVAhyOPQvJFsT06cFo6LW0Y
vUtYmardPA1P7EhK1hN0QGVwgaoRx9D/LCAEeggB2rK5fdSTUWyXVn3yRwXYe2HlW0CaHM/QY2QE
hNIIu4JJtrqwS7MTjMYuEly5YpAqN9ZWhaNfAtDBQJKB64HuvAoHvGUUfZNad/6zLN4rxLvL/hC/
/fSSzCJA/YcKUveA8A15VJUtZ/0J8TGotEc936Nx+GVTBPfjiU9Atb4QT+XztqIZOhTGBHugmS+N
ifbI9AX4qivBNYZVGfuC3dI0Lsy2+eEXwRfgiK4HmFM/Xqnyk8TZgS6o4KF0QcDm3ZdNnD797Brf
1oCeOQxdLGWMXu18Dt20UInepcCRR0m9t2pO3So7JGd2zSfYHty+kDr13lHEuwxy6PgdLfR91YiX
mlyAIc0JYDJW3AMiKMVPudqbUnWnxF8gbHXyTSYq/FyUdLzBcun68JfgnxoHhpla3u4953Ai2Tic
OEiKVX0nOaNv9GdiWOtDwyV1u398RGle5esrXaxN/d4fqL7WnfEL7ZFA8n1A3uwSXh70xJULDIbX
q4qYWa2xIi+fX+kOiKElp99C64EKRfMl/eB8/596qPCLQo+OMvTtxeZSI3m0PU3YUwuuWC5zRd5C
XvHMWDl5RwISA4rnegREuphazMMKcpp6VmEsSIL9SRjl6RDouN9uPhFOaZhn+yA4Oz3s+U2HAt2T
pdIDfuFc0otf2Hk3ow6t93uScimrrWUou86PmGZMMX+/JMVxwr400XfDY2gGGYfNMr50tBGnFOjL
5UjT1qtaaPBaPAexf/IS+CD6PoiImf+RHQJ1J/pqHBkMwVcSmdQH6oDP6Rpy9HziFrtSDOo9mZ73
JDN1VXXyCTdI182vNryEb/HrjWy48dF4R+OZvhLG+0pPSCxZMiFGtNR6pwRwEFyV1KejopX6xBU3
7bBkx5Bizzv5mOZtonBxUtUE7apvNaLSKiUUfzhF3at9GQPDQy4ruOxvxHyZJ3PypRRkWEG6IVts
FJLRB/z788vbU1Y2STh/jeYW10Xst2pV7imGKG/MH88x3nGsdkaZBuy8Y/Nr68tvxeLHaBTmu5RO
MVM9cjW55/pHODSt9s3+gFi4RJ83Y2xgNbPAKMU77OWOIaM9/0QHRzBeLmSVkhQMciwCVmNucLKu
Cuacn9nkkz7nREkBZc/voIpqo61W2720GFatyw71u5jk46F/Zmw+yFF2isY9TOkOLphnzG3XOIuw
b3laK5TxMwkB53QkcXzNx9UXpOw+o9/YvjKfF5S6tbRnREOSg8TwneiHWg4oazXYpq1fIrUxNvPf
MKZ+X1gB3sm41Z/nn4lkLWGqykGx0GW5hfPAk/rNGigH8jYEmvXRNHDc5YCevU9eItlceAaK69ll
LAzdJ+YcbSMDODjqItbiQrbPf2fX1b8JlR3KOUDVYSXoDR248+26I3icGkTWAhCC2KzyWCkBp7cc
0uaePU0BNKKQULoqdkk+U8BwvjgneVbz1ZJSbcurZ9qIuKkitT2E19Jo+yXFFg0okPPdevFxHY0C
Uaw1ws9PNSi3YGiCs+RhQ+YMAxon+HtzsMJSIPbEmCdL8KN0KfU9eYRmLyWfhRocLVif/fxz0AG5
AHXXQAQhDfI+h8zC06MCoKYxyNCf9iK7Ikx1S4GAleB2V0wQwB6U961FT+dghbuC/Z8DWsfchZll
msW5+Vn4NvwBTpkhQbsuc0ucpcOPimL1RyRpw0+XaHpukI0G+zElxFpjfAlaM7h/ef4drXy+3VIP
ZpQrcsNu4k6hlP8MhX6btm2taRVs1lL4O60W6kdaphGrpUlExwHOnl9p6TQyaW0J3ewVaFbnwQkI
szH0IlGVDGMIsG9y/rroK7Xb0n5fg3vMy7VqvRHYGlZIXEXReVcJWS/7UKDDoZ3ypbTC09SN41cX
inKP5c/Z6NZAWfUlwf3PwKb9c6dgA7UqwK+O2QWs/vbanAGAIe5lWtVCw0KY9k6d/3vJzQhrv0wT
ZplAXrFWNnJ8FO1HQZR62z0B3iifHT1pLm0WzF1nwrZn0RjPt1+s/QiEz4q2cwlAgqIwhfKsos/g
gpDR2Aj3lnidrbPbuRREh+XJuZ1pnV0nMtSE7MCixT9EzPZxnbOJuy3cB2aceK51FNdOnppOOnvo
kbH1ToLOg+Hf2tB4cnE4VcD6eQm835XI+wx8Du6u7o4LWlHdCE4Op/Qkm8lTnG5yGqrfD/EMBOJl
aLCKYS3nS/YCBRwwoQDx5ERZVrGLXcaiXb+nwWk8HZwVfEF8Us/5rGSHVPAH2tXMzZwXluYx86zY
ltSBNlxkN0rcROXSX8zduKDEqRcqwdlmXZUhfbncthJ9qRno4mO/fQ1EH7jRs55UHQXbkETIfR8P
r5mrhtVKdO46Q6Num/7vm2n9Zdpmikk79RIsZAJuVfKIe7v5xbtZUOIXIkNCtjFV6ccBZ9yUKRdg
qlcgIMxS+vbsIgM8pjH2362gR4T9a/qsbAo7OICies51uwTxwwvJTGlcKyrfWjYNyYI5v5P0tuGW
MDD4CjHzgRYZ0HMV9yAeoEMpX714uQoUwmte+6u+i/2jdqCOEIN8it/j4u2TcbN2xxxA5oQA2vsV
tLMY8gVjz8i5qWEQfl9e50UCMKsVsgNi6M/Jd3GyrKf7cY1TEV/VFDnL5Yn63CBYP1Ispu5TYsw7
1ZbKe4FMUSF4pk4AtcPIg3Z65wGXXbOjMgE2LKjc+92UIpvIK0rjKvgDitFuUg8Pn4/JLqdIkpK4
guU7L8VHin7muXkPUn1KFWjGCPuQiXioz+zO/mPF6bwgdbShDEyvmyi1Uz5V6wQgbT0lKXqHFb9d
Y6600bfzBzbTNV+wpJKKVw9OgUvm5dSD5+MCxMkvNsD187NSsyXrjCFIZI+Pl5dZTFFyj6yBFJUa
6/gP7x4MzXFLv8ugkd3O9zk7RY5ENe4OoeygX7Z7uPs1wUbmS6wTJavWL54uZN7YqGdGTilJTquR
majxd/4bAUgTvxrdVhtF+N+PqDvECgGg1COmFiDgKDgD4qB9jYnLXlyqjEV8cLARxd0/8faBevoz
BA6ajbGcbp9ChfieMtFwsLJde0GsNtmvLt3x+lwXyOnpCDOH8tThcEKjpgO0ez64hpyrkkqdzNjw
RmjwMg2ttEFIvMGlkHwnQNYm57WOyUZhjfb2oewXvbsquJJLiSeV9Eom8MOXeI9QfLkF7Ov+g8Iw
vLG71OEnIO5DwaRvlSAIUBxMAJPUswVKSyUdK90rm2VSXDdZzjno1FXgbn5dWc+IpUARe8nOzVvw
cJ9vSnkvhO/bxbDB4WK+Oa4ViOUt/7ja3m4p/17DM9tSmP53hXcIp08hymb49GdcLT7fYFGKwQMd
7FcLG27LSIKLBnHm1sfeH0S9G4Ptx7Og/lkPMfC5U/l3HZD3Sn2yJbjKLhwmXWvc611fcd9onT0t
j5NNFmNXYWyhOy72XI7w4X7goxRAC139CARRO5tnN9n1h472DSyvCZTrVUQJ4DsugPXgORJKviXu
VKzXts8+Lzk+kXI/DqXF6zLEMAekm1YFAv7l33NZMVu+WvdmIxBomqq4AihRHbtSr+LT+coHMBnJ
+H6EmfMjBPHdTMPLXvnLeu9ybpt8xqorhvN1e13fwTjFCdWyP5oakVOc/wYKTJsZQXvYXO/vTWsb
em/RlGJVtLfHpYk/juf0yecKJhFchbvH9twapN5y7KJX+fFOSAYU/N8Z8JJj3bJTtoAD51uO63Me
x6qStv99a8iDArhjBGAIQ2Gw1Hf9MPAtxqprooUxrYeTxwi/a0qk36JTM97z6J+BC9siu264G0cs
8wG8xRcuSgtYnjbVNi9ZlV7DwpBnZXs8oDjFNc2NPJXJxhxNAsPNQu7abu5AEySLXn/587IZLU/E
R1agq5MMSWZyj5OSpniB99Jkocbl2vdnO9XZMTDN6m5WTCIInq/TaRBh/2O9kxcBks/l3JMJ5UXW
dh6TsqpMInZus9ErMFlJJWcNWxqeIhMcznDxCu0UwkBEEg3bV05pSF85mpHxUKm11NfWTTC8Io3/
wXgeaTH13rOhzgUBXeY5OYZacbLIyAaXgmECVqYXOzgij8QekUqw9ASe12BfYsZ6JsTxrODen+R7
Xs1mdW6aIpgMliTB05jUTiW44MxHgBQDbp0yyYQE4UTeaWjKja/kgjkvBndAyafxkjAhgrBcY+Ue
SfsOHSaDHVXATPoJhNyaF0iz4Cj743731k6jtkiyATV+BLfSR23ZCjRStoQ03svR74b7H4XB6dzI
XGNFpl1OAQBE1DihocPGn3MKchJFfYJ4vZ8a0ZAWhDme2sN3d1A3zYujDKdBlNagzZF4zIgwj+kR
aEuNDB2iSmo5FRtkhlfM2+XhZX9z6Dhpt+rDp5rOXdtKoJFEqYLNbRcuwTDdDe5vyMAIBfTvf8ZQ
8tYzFJhWzgpqvlwNd4k9tmpRMLchGQGLnejfU8IeTF8IJ/HyGHt38nRDJNYoPbbh1sUvnSFBGK4j
VFI8QgcHmHUxuY8dm7uKQI4uynhLj0V6bl3et2Mje03QTmfPvrJpuHBbErg7UYekxrg5pdR7sVrD
VcjWrUOcMck2oeV8eK4wrGQEYgT/8IkPNqVqAVBMvTOhKAHuh/T72QXXcFzw2Hd0cP3e6TYqT8ld
mE5dBghDCXMSgFM4X3EpcgUKA+l4W5KwOMITO7K7kR16SGCFcNwNOXsCBQf27MeMKShkNfeiLfT3
twutPtG26MryldRVvn6pYzFD2qdyqL38m2XRpvaT6HOLVLMfPJcIqCeMAnLPEQ2mqwFUVDz53m3y
Vodlh5h3Wl3ULXk5uR0884MGi76nc+Y5a5fkgTtEX8Hk7yJt4yI3Cn5qBneF0Ckvri3w5B0MtJCG
X2LP1Y5GUli3/nvTMyuxShB4OIkYGk6Gdg5QsrSutcCnkAD5cnCw45cDmo9aBeIPiVL4hMM5DDlv
QP58GKo/XOoaH0kLu+EMWI6mRsXBmUkX+ZRKw8MG8S0LXBJa/OtbLDtFRrU6wMYHRT8/EwnVmCnr
qO8l+RgUSwZMK7V7B4ZBkVOQtcTSa3nZMWre3kqJi1A33ZHk/qCNMNMVcFdtD1Nht1YfgCISLspH
8SP6aUlhZmVK5LDMz85GLh+Av3ShX986xpF3CpoKUvkQHi/wViRE7hsqAXcSUzFZ8bWLNKWb4gMl
4qW/muWSh6o1KACVRIqmCO3E9qObHjL2c6Y2Dz4t0YxCQQeliBGvSjX9LfFjaMAL91tkpmNVT7F2
pYFDmHsaxVAh8iBegefWpc6zJz8wlYhSYzZ9B2Y75+gCQihwbphmGb1ou3wjf27uQgw0M0aGwne/
iFWAK8mb406Kwa2AYr8ZO1516O0nZDoQ4Ch7LwQx+ghpYx67isRqC+CTnBeb1IWgZyvicqVjTiOs
1EVJ/4IvxHJXytEuWqdI82rSATqCU4MR9VaCF1cppOb/ttZo2oEB08p5k/DinaPgqX7x9KT+6uwo
/QeXYAhBTm/qSHpGKqz+Aza7KwAnc28LnXbY+CLZAYXVSUzfgZFrPMqt6OPFZVlLUVUPhgM7pOc7
E6JjBLeHVxhQ9gdTqi5/iaUW/TU9+SLvbmUlVd3IzCq7ghDoBKfRabwLF7evV+ZnoGrYRJl1rAdw
AyAMiSvtRXIebGmOh2rYWeFkbyPQ7jlLTIlnoJX/qwv+ki1Mi/xHSFZZzKNsbnexcYFmJy7/6Cju
IYyGkvmV2p8UifFoja3XsD/4Fw965wjWn4yj2T8ORIDcHpOCURmmyw6bWwurgFA5KAW/PUmE4/CK
1qrQ13Pd1+vLIOxJfDmMx2WLTzXRQkJepHehJo4WZJWhOGiEbr0rQxZ5CX9lfNqrYS9KbOS+ABAo
mSyyVRM47XF+pfmZLkni6Ht9+6FgAuf6S9WFck8Yez5QsxYD/oY/k+kJGtMYoglzTzwXfEDjhrSv
BLdyKYc4I1f29D3/CoqYBGCMPRo4qwmmDzWM3aI8AAEue6Gb3SBn0won/Ygs31tic0M/Jmq+jJLe
ykTIIsTpC3tfHOYym90Ioim/JytG2I8HzjUJ3KnD5k4146cwz6xdlvlMv+rI/g3uIo2i8PnA+A9r
28HrY5GbKiKNMntF91nKz8Lzv4WxMRzoxTCLuBrI1yOBKvpTkKcDqfyvhVj7K4UGFDKu8M6FLr4C
r5Mmk+fv1n0t/fFTlrWSgBdi5CyN5ZTaaZx7oo2cDBZ4yn7+Q3RKMTF4bR5PIWXWXdoVjYQ1YEXF
cxn0dX6+M8PhKzC3CuW/V/9HJK/TK3v0+4u54OINd2yg6YJ5BJvlhFZyCkwf891b1BBQMj/bLVAz
QEHAcL4Lp8rFV26GETZq+08cgQSbZm/6VBEDaW3GmT1fpMKhljeXW8AdXHtGe8PvQ5fV6WD5AO8V
jiHT3niHAPxo/auo6tKyP77o2C1JmLUfheU24msZ1LSSYD3TOd02yHCEW7qZsmn/7L8Tn1qNh7be
Xdax3x/J/uhJakbVMNHOGy1KTZwHGP7MUPiFqQ0S3z9QeE6dEiLBCDEgknvsZSFUMOGHCvxjrDBm
X2Oe9Qj1TIhq5fDWu89eZKTXAiJ4nJy0t3EKFvMvVKGwbRvFEoxWFA2jX9sxZAc6wXZsCgrqZcm0
Hf1dJt+fo2I9UCZzlpN7+BBvrPms8xvTOPrWW7wJfhefc1zfNp9LVJHiTfZjFLutaiOenqwnfegb
qN5YMjHAkdND3DeLGA9I19fFoMYABcgsBR8tcfqdZt/delA+3d6Yk3pl/KAtQQQRaCcxqB0phqu9
JNIuSSzM8HeshJxbrR0pv/IdlT6N6Vl669n10x5RUJ94Dow/UNQBBR82KWU+KwfMt7XVKy8rwWtq
i/Vq1Tr2W9joWTzYJHqMBfWX5YVlEK8dVpPvWKK5oIal6Tdf0n4g0HLkUgukhwqEiRXZo+OT06tS
yzmGIim9JLHul2NwRQ0+2zw63lYScNuFmi96+nYEdpmXm/Cd3q+e4QtHm5xNw/mmMSDmeFaMy0QR
R9ghjm2xRTtTQJhgdrPltJGaER31Y7czjvKqLmr1TUlzFF2v/xiclytSST7qwOrixaoOJyQ9qM66
9f2Fv2ek+3tOK1JvPfj96Go4haOahHZZHTz66GexBMqSkRUa03A1YLQjuVrTO0q4yf6MfZOT8Zpx
0lN8effcSdU8rI/TW0JI0JHx6p2+iRkLpFTPiL5PRQigYmN/7nZ5Ej+kQsRNj5cikzXEy1JazwYv
YtuRNUy3SQu5JFva6nwtM85AMB0ssVxiFmE5e2MOmSrFQXX7RAYe6tiiMMlSEK/E3bveFB4rTej4
HqoJa3uh/1VCSnt2OGaTzZIpntmI5lcstLDXwIquQYPT5BJImp9unIGZODXBg0YhGt3JtQVggwdd
Oa2pHTBqswvF8etNtpvNY0ZJtX56vHSuZ18yQfSyjYgNpMBV1uaIuiVPY3hHsE+qYEP38rIRxdyg
meQ7/YDK6jLP9ImPqFQyZjAfA7QlDTsqzgko2EYfOYA2J3DwrjDxmcsUo3egRxac/j8308xr7F8C
aCd23lheabe9yuHr6wKt8nOn3w8I+Y4Pojj5Noh1atf6W7IzoLmFfg/kQBSF9Ept0t70VxvZB3k9
9czfrhOsJ0Q9QLWilir76Oonz0JS0RNOXT/i1saJISijl/N9m2ZGXke6Ci01smyv78XKTfovcZ5+
yO8TJdyPzxioMWui4p2m+mFN/1E1siOaoXyMVQDoyl248P+kekdAdSbRpKJVQbwMS2o/6Upp28yH
3uGkCgcK/GQUB9vwzu4iMzaJgNaWRmuDgL1tbQ86wCmfZTBFIK05t3uJDh4dHJDRhCIVEXStNYBI
Ti6YFTiqyeYsUHkJ09GFi55V/EkA846AjJGjDKx5GiobI6GFYjXNbZdd7ii/mPg31FRyvcoDuDIr
vhfWufQrkGr39w8EGcWs8eUsqEwOfwQNbiN2eTEaCYcIbTat3DnrdHxmITetBSWTOAZdRTQyg5I3
8e4SzOOGrf6cU57o0DfcHSOxhIts8djHiUsuLxjzhEVFobJ9U0PZSuvGD6P02+R7hbN4sKWVI3M/
jkdD1qLujml6kax0JNNwrO/r+aybz6D6GlKnlblKdSvPZaZYdfbJ9KGNkmffVhtr62pr0VljMwFe
UOee+Cy1mONYoxZkxRePS+X0KiJ0qTHO47f/aQk9W+l32kd/EcZfLpYHNn2y8KxXgD1FIHTIm2BB
DD3M/AcbENnaVsZrLgcoSSiQJGrPvH6V5NNsKPDOn/a6AITiXGSJ/AsqM4X3uE95WWdTJZV/cPa2
sA+s6XpKw3V6Qw2IOTn9cF031oGsJ5zMJEOZGROmMFyhRTAbGWYNVHDd0mKKzFsvANqRc9Is9Q+j
V2NqIT13Z9JNCu9l9KCaKY1Eg/Qk/sqw0l3OXTpQ45ILqtNiyx4lifAKLYibmyDsymIV9qctWgu7
ooundJI3g+F+c3F1EY26WotRBfqTTwGUHc2nM2TJABSZ9UUGwcqUqpKKwD/DNJLGmSSg8GGQM4yW
YZK9v2chFzrKd/LAtXYDRo+1tdj3QE8rilQ5KIDQ97tZ7zvUrmK5tmDQGix6Jmyw65InJS0kWuj6
fuPbplYEXty83l/OqM3RLq1XxgreYJMPb4uBL1JwABpiNwVnTDjbhqPZXU8eLZpwRabKnABrMpb3
jOOmZ8IwcUxLiErURt9xOlDb1/C7lVcuU6z1YiwmtGy/TGqxqs3wN/VIzbILvkgxj7DLHfJoZ9dH
00MsTBecNeW03+gwZRy3kQDeydQ68GPiolVS5fhuiY9CXfC1RrP2lrPclzUxopLXk+eM4YigEZ4V
K/bh0nELB99oxcRI/X5XzwNMUEzlAOjcTNdqBxoZCKpffcdduwJQoysS89dcDguBnUv0mey7+gSf
j6IF0O7XSjRlD0Gx95ECku4TGjDB4XQZ7YyWV4e669ZpNJQ6N4Iw+zVj7rT9xSDpozU26gQQ3dIa
aVROpUP5EkY1RrbHJQL9wm3JICvyvZrRdFW0ilmtligwf9Drj1Ym5FQHHmqcSeEN2Fisq98oliZf
iCN15w5+22vMi3TnOGTYwU471KZILS3xXz8hlNOmgBNLAHsbIg3wtbQcM/Wb7u8TDk2S19gfmVeS
Mq4MbxS+lrmjM8HvhQaUoMandzzE9wY8QdaihYg8hDM48If1a0oJvnFOREWaIZIf379hxLs0fRrn
200dQCUc/5JxOikO64U2/hOgcNyTKZGKFZbodB2JRj/KBcaq44uO1GDj7iQZ4Fq3kmVApOXgmMRQ
qaKD+k0alJz461DMFuzcQZUczfx08pkSdl+zsVLmM/jLJmYznfM7LCLXq2DXFV2sz648/vQmd8sS
wxCadg8Kog+xaJvxdLvO4BXfmpL6gJ1ELjzd9cgeUiO5PRf3SjRTYUbfvziSs6JUvwZiXrzsd/VX
+PVLIIBar29RcFRyMMEXZGMcDqEgxMM4VQSqtFtlnjM0OE1Vvl0+fWXs9x3EuM3tmZU4SS8Bj7qr
OAedLyORpGDSpGsI41hr21qW1qXC3uaeouQzXOxGzUp5QVJs/L+i8KcB2HVEqtn9ScNZ+6mzMnRH
vdX1WJfVq1sSC4R3Fh6OOf75Riyvks0sCFMtZwqO9sgFwr1xtgSk3p9jOIZ0zTpmBURApuGr3eT3
ln0FLbwo3yffxyNOYBuyzparbeW0tia24SON40q5sOZQY5XUSzPUOa8bVguiZFc4wnuBHuQrwiIg
22hB6Fp2scEiNbD43V+LPGDST6IM9iWZmKk3uhNg2J4TdGYk+EjUjaRPhiJ2vIZ+FYM9xSchbq74
tsJj0s08EcegUGPAmPleEpPgirbJIGNfS1uHMyn99DWgl2x3LTFBFCfploS4LLqqKFIL9UL3Ds2E
+VbRZbLnje36u7AwydJYg/ZNI5XkztBQsHaMn3evO84q4RoY1rt9MwQrBGGQxkXflfIJg8E6LH9g
U0dn6qjuq6wUrGWp17/VOxi0kisO0045J4yEZXos4QxXhUlyMFqLakqPZG08KiRoX72mRoKHE+3o
OcuhI6iWyd4d9AtEOqXqS9YWPOEKb5+yKhsDkUa3T8pBeekORt5gO7hHNhH6yj9WAc2wOFIeTvkN
bK98gT79asfC9vkAN2K9L+wy91GwY4ZQNBNe6cn69+FOjOXX9S24MIUiZoCWhvtqZZZP9kuQbx1/
4Pwf2DG4s+KH1Ixb8CHNOSL+yejcqKV5AOjrTy5VmyWngZ1DQQd4y4jfqddcCH/PMOOds6rCHdk5
CZm7EGR+NTYzizfPI/lURuSfEpMkfvV5rq4qbGpk3TgUY+pe9DKOhnMrGtV4BfAkhCLtB+uuWdDm
b3JU4DmH4pAFv1xXsgwsZJzzqGDHdNaz+V8rqqtsyFo+66xC8qs1meWMn47SxzK2pocG70J2Z+N0
w6tFeiIFQtlpZjZpt1O2TYxjHTlDx5WntZ7IPdm3TnE+QUOnC35GuDnknOtJ1S7ycaz6ACaTwZBp
mj9qZvKmXJv6MLkBOe5f8BQH2EtquqYCCBE8ypQYLqDdYNSeVjDDwkUxMEkvgxvHURHIPkg6UUzf
VMQD7GT3r7kmsOAmmoP0iGr2EQP4q37dyhRtNtr4ITFMG3ZHd4HkK8UhWcO+slV1jHSMSpW0sbUh
hGj4AYwYEpiQBhTI2KtQAwvCk9OfIE5xAv/C9j1/5aEKBkLJbHqDtV92OuJW89Qm5rgwFk/t/Lw/
3RfkUKTthFycIVrU8mj8f1vND1frK+KpxL9M8SuhUq7NJCFqG0UDhSUKEGqHjh/wgMGagkSwA/0M
gFPms5XN6LJmXVzHSHv0H65KAPxuhjUeLMyU9uxUkyQcJX4LYsdUfBqq07SderHBfIxXUdRG69i2
/lpJTuAN9tu3bcRQf2e6yyMgRBjq0epsd6cIv9L1WD+GowizmnKqgmuUcaoXV2CcXR11sNtfuUhS
ZMNMXb3zGMZA9+nrd1q0Ryqp0d/Mu5SUJ9j31I19xwnxLt31Vz8jxFukYFUVQzupqquWTN8RrEfd
VREu+Sj/TfwxO6TZmSL3NUVvQsYoXH3RLX6Wn7JbClNk8iT6G9PIs1CK1HM+8KgEbsuahT7ryCso
z+7FILudakU/sFAr06zLEZJrqm8d06Rqp0308aqFwWo5uwUkGXmayfAP/4NoVV6SUZ/NPT0FDeGu
99BgCiZbGvaPwoBfbrcdAfeXgz3KxfRI/GqTY/EwjMgyCFmAELTQjKnUFQNm0E5OROawp2p9DQmc
fdbv71crFKpy3Xj1wGxcWUQKG/+XPPiJcaB4/XI7uVdhJimc4EEuFDeSw/4mQCsn8v5WbzLNaqEZ
yK49BfCbpqtR2Nn0RDyCneTnsb0Sf9wIzm81C84ynM+k8BV7weFdFETcrYby3Uz5D7YiLObfIYlm
lLAEa46jmRbCvPG0ZVhwPowZDV+gcpY3KjAwu0uklLtUZU41+tKLP6WLON8t1j8+Ux4A0B9ZkrH6
JDHtgwCSoO4/q3QYP+3QPVvkvphN61hmHSwFCO4z0Zdq4BUA9PBMouN10d6sxNT7tRvzXfcjZugc
XSDjIrx0urkMtMsPHE09IeKiJNkb7wN/8JEWC+Jaj8Q9Y62hUqcEwHOACMV//IUbGLBT+sAfvJRZ
JO48sYyDOPHKowm2tMk9yW3qR8zRCEkC57YLmH2JhsCh0IbbAxPHATAjIVMp6Xn2Ya+AmuC73IsW
QYCGzrt1U4xr5EwZ936ReXxGqVOcX8EESIY/d9qj79eivX3XurqUtNja8u1f8Bo4kM8f8FFiwY7L
TJMDfli5scy/yOTVyD4dZcRLXNH4wWzSYBIUeyO7B8zmOHudwXgJvazZkA9puEFoajV/7wJWRxOT
MjzCox9BNLRhJHxdOfJjBKImae7QQYtvIs8mJXo/0yGXUizMK+NTbHgtzS1vzMagNClyQgwtYyg7
Lc1M1f8HIKcvzoK+4HMgFFLPhv7S1HDYcPmECpbZmCJzY028To3n+E2UrSrMPU0rhORSBBn22e3P
XdVBSIEDS4dZFAMdehWSR5Ccqk+KnXiMQiy6lDW9R4+wu1Qs3SXUyIDAVB4S8JrjaYEH9kz0FdlM
mRcGdpUIuJKrKMg7Wtt9GznLQLs2+MWlKpu+CwgoLtv9HTzEzsrdB1FrNItatKo5oNe5Y6lng3v3
tARtDIAzUY94qiK6VBlK6X2z4lp6qwGRelY0oH0zG5q2gFkiE1avEgAVm6R9oPle4ED09ELRlkVv
4eFsEgu1kqblS4Q0TzXmHBbxbntsOtj8B3bAm3dyxhazAu9gIoZZjV8bNA6YHU5H+Jlia4VR3t3P
YuaC2wNXE47eLDE51Abj68n2UcXL2Pineg7PHUA51MUBoTmM3kK5oUxej6mEOgVJrU1YS4bE7peQ
viuiWggEoqqGxcoqhOul7M/RYsN+v+u0WdffgLX0YNWQOkXnGBLzaXGsrhzpu7pno3wC6zckp039
4wYHEp4DgiZKgD+ZV73i2NQVqY9wFuu0shivgwpRCXmmK5U0dKnBMC3Tg1bdecgnbC+m0O0+VxE1
7Ga8OaxFodnwl9uBorkHsX4wiHaiswY+MU1F0epjmyd7r4eiTqci4KqaJVOT46rx9cxbuQj+K64L
BNpSMLA/MkQu1MZmgGUVz28nEzaIBzZ2RcQkZlkPzbjeQI2NEoI6YXeIF6PAzgBgsMwU24omub6b
DydBp5Yh/EtBWu5U07669/4HUGXtg5fyKmspdPQZFfSyFIqWDbkVOOAFwY7TlMZGmyDMHcmA07YM
4i3KnCzwretpam/CG3O2QhVOAEXBRYOD7le4CEEQ3j+w9Cv6qPAll54iDYhK8XYahcnvFF29eCw2
QnJY7c3BL3GhdWiJVYRmndBuAIpVBC5TCpeKsl6wvmX1s3ww1IxallS6oUy5mIo9Qhys4bHAUnnI
iJcRu707FNOcWBxKMdi3lQCZ29pARJCY9KAfF308XXom0jZTBevZhbUsSwTDJd+Xp4J8SBGDY8M5
gw78Mu2YgsDgR0DCNCD+b0Ht/W+QEihArXK0f2frrjImj9nGT0Dm/DxoGFy8BtSATLAtT2LlKTB8
s8uk8Z0DAHXuW+k0PzNnj2kVGSqsMp5QK0hcUpr7qQcdkOD5M/FiaBsQqUWhWOF5Nkm56PcsdSWN
hDwKf5Gm/XNgu2ZbYTlxRyVyWIB0W9Q1bI+uv+VbdJa0PinmP+kpPW9AvRennyHqQ5PsFh1aGLDt
ZgKHeNtsAQGUff9gjd4CJEp8RqNnKwUyX34Qs8MgmDwwzAij1NCqot9ygwLg9IUsih0VOjJYyVdO
ynmmS0EFdh8pngYbfMtLVE8hbH/aH0qMon+H2iMa4akX7g88SyWavSd+HrBS62XG3neInGaBrTZ3
viVUD5deciWUxeH6aFtpgFjMo435fD3XhI8+53SFLR0qedNhOb/jNYNNRF/HYtl5GOfS3hiQmDhx
8TSD64lzhfpBA1FZ6BvpaIjHrpGY5HoMXtjzKb39fou2iPckRCGR9QYb3qETSufHrH8Rr8dqnHlU
85hXtg1YIUjqbJcX1IlJqpfjfK8t4ukz3F4MY7zarNKfDcyIlLMm2SRgNjdAnqiuNcRnnkM5TMa1
nzWlvX5Y1eGutIedsyR5ullI9mubzA3pfTPEOz9iAAWj0eZVjhxUOiaxRuQBaN2UneglH1bv0ezw
aVeZtu3D1sX8lb0TLw5Lio8kPF0Knvc+a3jjPZMcrm93cW+HcblNR7RBLQ9l6WgSlbmcjc+sG4o6
fNuRQMzTQMzJJeJVCGsOfUYLymdyH0q2qiHLtYxO3QqeRfrihajxkixusCNlLbix8JocqPYVLxWU
sHkmYmFDoYUWGPM9FefTaa4qH6xV7E68RDpL5iqxXsGeNH8VgomHeXSweoM90i14w5Evya3GEEaQ
TeMflwwqPKag7jiFix3HIc6WGCfdL47sr1fx2fyHKQbvdS46yR3KWkSawgZHHLXTtWaNonzQm3GF
h5u94MtaOyBj0kNcaTUOwkMees7T51I1piNA60EeJMtGendoqi0kOuQike64njUAhKQd/4nR4rEu
hC+PsZFegK70GWJjmrgYd9i7YiCIwFCffecZ4u98uxr6WKH0xT2b1oj2nS0rorqBOOx9AlA30Wbr
5ywRVz3louASTeg/Y38MAoTid/E3f9mOUZmlF8TwidM2SZh7kUzFne++3c8tb5Mqy1OFI9rWW9CK
bkeT/K4Zl/r4dxVaGalxJBd781C2BTmPsXUR2AvU2b43317PdjsRyHjSTBsRE4pIfkmAkrUeT5bs
RtmjbUT+ByxWSb9o7ziWpkX34g767RfIYwXAFyUqbvoFE6cv49MAeBeloIypK86r9d+hqxjUSK2k
o98J9UmL6JnnB256wSzmdrLXB2jmucTMVHrVR6YNmZV2USs5A2KCN1zWyud0ymmYqkfROicJwzD5
f6V/f7PNaMVssplb0xudT83vYSiA1DSXQoJ1ZMz+rk122YQrTFJJf0wTc0zZbjFSNuZX4YD0EZaC
W0SMWoqhvMCyD9lWzvRI79sO+zf8zeZr7LKSnbM2ypDk81U4zwxrXENqF0tYanyCyVlIB0YVsjoR
ph23u7rzaevk70sCCFlvGxunyA77n+1VuCEOuiXiRj9wGLSQxsQmYXUT+j+1VSmfkhdqqa4w6hOF
sVnp/kyx8cpR/uei4RI3bz1gqAje7jrWYUP7nBSakNaZ5WTo43xkp3oWrtG3Jpq9KOak7vDJb8A/
VAtDO6CIb9lTVZzqLRApQQT01fmqzYrcjmybVustR1jsefuRevQaZfXmYZzgK0Id7sjwyCA3elsS
EIzE+lotp3S0pTAhAXDJ0wHorfSxObiu+ZtN/x93XUwEMXy3ZtsDABN7oC/V3UB590M3IxeSF2b/
64MiH913FYjiOMvZh18z3XC4ZroNhY58HXHIv+5BAdzMCVcQxsnYNU8/SFvtuquj0uRFMA1zhg4V
vbNrGb7sMNdBBBim8UiLGZA9xLWKVF0RFtlRZ9xelJ9/p8Nqi6mZhwGwFaMgCuaNW2YLJORLs8Ur
zb3xnjOU0mzqlZc5dyCorW/EkesVN2ZrYWm/rdQtiP/Fq/9Jsv7BroUTtWCjV/WY/1fL8VgkQzR+
IlI93ICEnfjl+ZZtzWdPB5iYDbV/k1+75aKUZCqQrRTG1xB6IHT9dA0HhibIvDQ7pnfYPBbqSWEs
mS84DkTobK8LmSWCMRQepM4KPWz4YZhQ9Pc/NM10CwqScBqPZClx1rRqQfbmOLOaZX/+uVRcQYLb
hANMyqKRX+szeuuffyTMbEv98I/bSOPPytCc5yA3HxHpG6kC3pNWHgh7Ty9HXNtSZSxt9TBYkl9t
PFSPG3UkKrftdi02s7gYFgcQYFAXLOuZmw2XtZk/T3+xKLsLVqH0JSejBH7QBjjFVZkRlInqf51S
rjmN9d3ftTNRSHynpjza4tzIjb4ZhppNgUA5cMpl4St8p9mLP3h+5JkoDm4jhKFwRrzsdeVErGv6
c/iIJOXDfj2T9DaXHsiHHGrZ09sO47i/Re7MbHX+h/dq7z9U7NzaM2WZpismP95pukliOiCXvZG3
tTUQFBJqtwCncJC3trUoRoFuQuuuFet/ERO+yezlT0mCo5SSu6fmijSNCo1fo+23aWnv7NYe9ZRy
9MYJSJca0gq+u4ow2ojNtXMa1jIT13Qa7AcGpCqYejxRf+7p7vjVRGjeDYeKcBr2yYpvGJEwMcJV
D0BITih07TJuybH4NeFPzR9538K94WieO7SwM1FE4TwNuK6JtDgPTQ5X7jyQvsI60jTylWT8r4tX
3tphtxZcx0npqwGW0ffAZ+rePRg+ptxt1peVqCAntdK/CXN4D4JQCcAy3FmlnTSAI0JL6NOKCPum
iWqSqWKlz5iOPaWg+xcIrjB8Y4IQSwFPQb5H+UAc26u98DlPpAJgtCke5Be1twWRKJb0AArCkc66
GlFdbRmw5OA4Yv9+zbt+GNxQ02wqjQ51jSU74eJjcRav15d/a/zAyYI2RozCxJVMv4HSV8kEKEWO
QDlSVZNxZv4zOi1JHb6k3Cmu8aXQ+7Opa9Sw7Qr/I5Z87CUapWPzlm+NWigt1dbWz9mGpwdoTun0
GxwFBhl2XR/xxGn7AWKT2ydo5yI+i+E7/zgQoGwx2WGGUNY8oXLhVvzrOJSEoNXV3FaVhPtRrjsw
lbfmM/ziqxQSvbZLN+jPgh0ZR0QkezBney21VdMxFGcZfsoPzpjW/1qGUMdLQ2gnF4D8whoPGVvO
ikM6tU26Jru4ST6ahmVCtsIK/Z2Hd2lx6KMNgMrF+upVbNiuJmbSgwfUlyC3wQQBt+JREfghvCkr
F+WxDS4ZGaESZyl+xY7jzmL8yxC/8Wo4a5xSGX6XKCVyxcP3lcx4Vuz5bREJz7X6OqR3+oeAcr2I
+yvWiShXYWHLQ+TyDHezhBxw9B7A3NDfz2pJJ6vaPKS2R+JEwtk+Rrsyy4XgxG/vYpgFf6+i1JF4
8Hp9Sxg3s04lB7NIK0VY5B7s3pGE+RCBLyLh8LTaeOTiHgOVC6Qq4fjhWWJ1cM4tXvfeHY7aRzvN
xAnVkYsx0BoY5AqSeiIZpUFVVkXe2WJD6IZoUrs0/j0WDrq6MYoQ0BYT+J6LZT6DC6VOQpaOlg+w
aBjHoEL2FMssyGXwm6zadzMg9agGbMPqvXlPh0FbGizN981lvCLMgQyswG2hy9RdMKkEk296rifQ
HllYbV+T5PPyBRay9y8X+Y8hIoSM6ROPKgl4hS1B2/N/vpI/T5MdMr8CCrKyfrPBCjCITMPrqPMX
bGohznKjXu97V+anIYQ5avaWw0Z70NGACAV+d8001uuLbrnGWkPgkC8rmANCrbmGq+Fx2qdgLgkT
rYmAF9yxLwz9IV4Yjzx/A2lGiGlcFOteqh9Ii7GVC5ynH17xQN4/pJfnbEXOnwws4u39sftsbIzk
dGIYEGM6k9Ir1GATRT9bC+BK+/1GX2MTvbQze3jQ7lsaBYYwEWZ1Tj3XfCnz9TV/sbOeBpFT/EgG
JIu9FaJ6IVCEY3NRQoCOvHNuIJw4QL2ExTpAdUPlb1c5ylpP8xVqL8Y0CrEICsit7iHlNgI8sf0a
RbL3vmD1OYv2HEnrUpkO12rzRYk8cupL8d8jJVab/DrBbw1wqjaGQwQfrgbng7Xa5h1AbYOxvGbs
djMV5+t3WN1BTCAtda7HGJGE9drc6f+DIqp2Kbe2xMNZdb9CNbu9RtfIEtMmmFsrUL5NB8r8FwE1
6uelJ1hfy9kc/rLF9XLiv9j/UlF2PAkjem7Bq1AxsFHWgdZrlkRz+aru+6kVWzR4lhwlKsreQnDR
bTrCXsFhK/4AP05zl6Lmeloni4orJJR8iWRbdV0qLeX7bIynU7CNndHYOBX09lWxbZuBzGlrajl0
H9Up8NMk3YnZvvGTdurcA1GHe3d9PYxSDjdaWhD7A+4mIVdurgpvLjIpCGi5OhjkijnbkMmy/PsZ
hla8eHNM3dX+ed8MfQBRFkeRBDa8g9pgy+OCT8WgBuU4zbBQfVpbN/IUl/VEkD89au+86m6nGS4z
pRRQOfa7V69DWHcq/hBFnz8PxCwcaAyTE/+GRSyny+xLKJD148pcb2ad/aLtSRaDkWVUN7xsP1Hk
Kruhma+YOLRm0LOxoDmWU6uZ+EX/dqLh+C5dKoMFKMP1RUb3deEIjWLrcEimTQocB7pyUXJxFdU4
mex9ok9q5xI0NCxK1KjPE9t2Li9kAZ59stkknyXsZ4GLx3jtEYGOLanQSrlu+U4k3tZkCUHs+i17
kGyM5i1EbAOwHBvm0sJjxjkYr+uKDp+gRCowTD6pNTIRBGLmtKZzRRinTK+p9pQzwc/RnwUMqa5z
bVcKN5rcJKn53Eg0UnQC4onoUAEMNAaJ8ROKmV+2leYl9/jBweNLwJqJocMr+YsKmCfaIQpS/9mH
ncnStmORFUUl2rHBR2UL/Hmq0pY5h13zKoEvuj1pzRdtMaL6IdrQhZi1D4BDxXJI5aFdzBUJ0UBp
tbeMTf+EwTQaz4WLi0MJtitRfjwof4XgXgo4JJY1csW6LD/eAJOwbywaHnMmlomRa5b1hWolnRUO
R1GBx3y+xNqPJR5+40UTulNuF7487I5jgp/GJzdMWjT5UWB0w7ONcZFSzhffBZXptXntY1kv1mVJ
/wutKXyRksSJ5+UwP3eaWmkQDxhop3YronxeNCJWJMPmYlCSKpWoTSTSekLsE9CEq/m/ROihKot5
aIkComYxnX4MJhhoWiVD5GClg/0IpQ4nnkjc/Qce5dAZTvktZO2DD5OC/NWH/XZRT6Z9TglJpMyn
0NeMLq92C+7X14s+ukNDPufTbiwHH2A7TFmxlTHT0BBa1pHlWBYxzsQnpWK659Zw1Pf/llt+4Ehc
6AnZrFq9Y6m+dPN9Fy1Czq24NFN4Gez/74sGOP12x1G6OftuO22IujHkm71o7zNA2etAi/L+isWZ
cBXv72WEqzihGnhtbTRtZiyQW0McscT8tf9RNAwYwihGtLIqbrNVvVbTXsCCUk52EmsufKfLO8Hw
rd5ife6egbn75e+ZoDVZpKlwgwig79/XrVAcf6GM3NCJMUyMZgy2ptA1vnJ/yZb3vea8LdvbSIj7
pCzWShbwxml/8fZlOlye45ek3XQmeU4rXNBfss2b2nLbrD9vzuaZLxr+nseAPCHQMofCvJ342Tvk
zo4RlUa3XaPxSV5NFDM+u9e7qjbGplCUl2T0nQuJ7uiSj9FA5i4arOtGuWGYvMX7A4YI5RoZQ6Lf
yU3OnUCTfQKz6G71TKZbw8F9CgWARTjDEvhHFqHIvnStq5LyI9SO8eoo2S21L+KKHkkyW3wRrWnj
RB6fEK1R/8R+zTLjrLezg5xh3Dac6K+LES2VHI2sSGtQge5Li7sksVeAV/e/5+tSWu9P2IB0Vmjg
ARSRixUvg3yGh5NLfr+YaQcQuwDrEl92A5gdpBa5JsqJFllXXMDZuU50Wokq/JIrexf5eXHeiYHb
ScwPGsmJ9eArpfM/LtXL2hQJ3cYYatsPVA9cLwJwSItTUFcicq0FHRMnowBPTp03DuLmCD0aJdET
FSv0WC1J9R/GSB2/NkUJE44DayGtYSYjwRsBP/chplB61H8l1jvMclMyouOZXenWZB+j/A/3a2uw
6z2enbJVu8LmAVea7c0fEikmlb2tWmEYEtf2QEgq1fZETRnTmrCZGZyjxSAjVug//X1HkgPhZ0pd
oVJiChTMbMuloKhQvivyVZcy6f3k119vTkQxl+p7ilktZ8LkZE5b1ayGZmcFncHetsQz2d5uq0j/
x7eAvNJFHVdmwWmdPZy99v5z+Nog/zAj7AcepxwNRMJUFTLmJwfvqls9ys8VNvmCYf3o6EpziqTU
HsGMf/slW2Z6wtO+zRNKI8DLHcUvOWwiX8ehRhe3sBDaK9r2QapqtM/lpsVA2Z9iaL6cRrncp4vO
rzI5+ecny629v7sBmkqlwOMw5R0vKOPjb70sLrNLkPkFGTU4yzIi1SCwtVxiHdFiI1VkqPMTYmyr
dUDGVbdi7cgXsIqEYVhcEoX9LR4gOr7DFSODpPSPoc/GUhDAxzHiEIHfAHBYO60VvBY/01Bi/dwi
SBqjkg3N3hqsAfYGa4qnObdImTHkso46Z9dKfs4bY8NSvImr4CEQYPqjBDSQHT5giWxQT5YSdB/R
PsNgl+MCOOcGlOE9K1WaqT6GeDX8NOObDDAbmUGPrpf/DXuc67QqMjYz4wiMwa5cSwYOo7pZbkz2
OGldgFKCDdqBY0iv2KN8ErF76HwN41rTcsRP7LBDx4XzGZwvB1medrH04S+SK61MLQukDRSpX68D
ktqHVwYd5dUIVtkK/Oh023XA0hhtjH47nvcgye4bOu+0YuIKhnDAIhGoMQl5HP35C0dU6ffgDgCE
gzsqJ9eesZ5Ua2TACcwB7kEPBtz5gKbYlWFtxudLwXbHdFWCSHjdfqM7zPsFz6LSYP3u1qUHeunB
PXiMuyjv0YCcKYdppgnQpdoTePMFQOFFCXnj3Cu5IutxurcmnJON8dJIYDEu4Ewe1di6HbUCN6/h
Fm1MlxJB/m9Amc9Kg+nGCEr3WlPlp19hoPO5NmC9rNdCIO9tdpZr/2QRMZN+BKBQl30UpcZlfFc+
NR/nBUhNVAj/uNmczKWAPDRC+bjmAgZo0hqhVeCPCsTetAUkA4txxwiHC2QATfLXZ1V2k1nXlC/o
aNSDlDLsmmGvGrtlecxbjQgwgK9qqVDKONv1UO3IMqnYLD+YDcoxasBEHIXNC7amLj6eDCmqXL10
aoYi/KFow1vht7D7KSb4vCAGg89swrbcs8cBknPuub8xvo+rnbonxwM+Rl5rwclt0b/rG7VgApn0
9oCAHx68iHFtypa7TiVwxRphi/wwJAClFgA+4w7b3JGUweGBEbkV7PSckwQo/Ez7bmfJFbOjIPRd
/PKEBk85mTI8Wj884zKfSASYmhnYZ6QYUNpoNFJU4BN026QAzFmNVlK+EL5I3D60qWr/3Z3Ybgtq
JJakvGOLk9fQSaHL5K9C0SZbosc0KjTjhAs3sUM1rhezmmRR9JLLQtByAZg1upcsZAo5dlCWKz25
dmaPTzYf17dNAppnR6cUih9AfepC71bH5Z5da/EXx+gr/zyQYXx0oE42MoK03DN8IVBDv/M+hsm+
NfYlw8OUdNKOWiD++FyKGse5LzmYV8XXa5p1z6ZWuKjcwbuw6dtcmho7n/1WLj/BHUJwTUVuSJdi
Vr4/Fw243NG6VfZn13ys+FJ+li2cK88bbetTavJ1CK5+YgcmooIufDYVVTawPS5OPRflHFhbtq+j
/R2xrWYQtMDqWj0tEwQZou8sz7mQ8iETYk+hcMZUG2Icv/zFLx6OSt6TOwhdvp0MaDUoTTlBZXYM
BtGnGW2swn1z64K2FKYTUap/gTgMOZXl8pdu+3TA29I4X0IxUi8S631YWU8Y4Kj8ynxQPQBiySGW
3LMFjloqk+0N+BphLpkK6Tm8gOhCpfvqIO7ODUHT5VF8CKiZMZD2sHP+y7RS295FraIOhRc7xlfJ
Ij+rbVbaKiprDMMhENJlltGHbO5hNUD1G1HlF8BPX/4/nVZV04UJIFkCQYdHJHEdQv6a+idm1QDt
NBaqqYQct+HJ5cT0o7WDg/0HH6ypmAzdnwjSuXBJuTOeppOo2r0t65NWxvn9s5RXAiUXnTLUyyCx
3SeVczLIXN8NHRvwIa71E24SkuuFmpcYKfsTIoEq5vpuI+3IzqMu5bL71ZXhoR4U7nUCxPEW9mls
B5t85fWuyh4S7A1GFRZ0WcrBDgAE+Elq3jGtUPMmL1rTzYaM6jK/ScMjUHGVr9olRy4j3WcEC5AD
GCbkC9HZ9sPeVA+xleC3G1E3NQlNAXkpZUstFt0XleFmjtKsvO4ASsK5fHpzbXu7O2pn/LP7UB7a
BTsZj/yy2AK9+GJvQPum+t2KtLXiJlJ2U9v3g+RBLDh9F6k5ngoWmuo0K6XH7SCNjIF/TPfO95hM
gDX9Ry30EOVKolUdL/x2Gf6r1ZY8xIvlRxl0Tlg28Zapa0MJhfmR7iEhJG0LG6kqVwwMgS9Vw8gt
SReO1lCa4hY6QG5eTNkWTKxJhrHZpDCrNtVjScWFHLA0RtTCpYhki38Wrg309jYRj5DY5mEQAVJW
f1+VZMppfYJ47LdI9Yn+3BBE7XR9HOwzHyqaEXIJovfyVH2ItxpJzvfUNMzPph2L+TfXGC8HoLfS
YLQrJ7OBTxcEaVxNO98EP906xTNZqduTNwb5n6trqDMNN8XN+UpSulXddW5jCcovnNxt5V7MvkRy
tuH72nWqKe3k437Ptx+Wt4Z2pOrnZ4mqMmLqZ+Chq2hssyQU9l4s2O20a5TXt10wtjlrmoay2BP6
Na1oDMvo0rvDRY4nhjHgsoUKo8YOTTBYuKmBYh7H/a6UABfzh5Q6sf6IBRCw4AlpSZCxXx+d6Pv9
9i/cuco78oMzuUey0E7PeO2wNV/3yW2OLfOneCNoO7MtBVcBSkgTQmCO51Zyw8otNHytY2VEL/4k
vTu72M2yZRIBhATiEp2EAQbJXS29elpzsTJJYpAZXleZJc/j55T2rbUuRKnemKuwkN58QZKYY77E
+5MfwRTA+e5ZG/c+dO6EfqGsOAvdJ+oiYjkDjGFDbnasibRHaW9Smf9somb6EhoOhbd4GhCAj1e1
J6pJI9cnN1g4DUjDmZ1qAF2lHZgC6oANRlGdejqK3CzmoZCgGNgAtXYwBnF1lpK+hDxcguU3sQf2
7aIZR5udWpUUTe3gxgJopoFma1EYN7FnY+kr55lrifHTu018rOpvP6IVBAfuOXPN+MNpEitxA2FF
+6+wkYRQBR/65Ruixc3l3KmInWBnKP1yP9yI7XyFsqVUwIGq3dCJCu9iM8HaJu/SEavykbYiWRf8
055jTImCDHxIDM9rnq5Zsoh+ljCfHN2ac7YbUG7VGtR3tTmGZtKGMslWZknb2roXTgCK4H2i8Nmp
4mnOi93dhFMT+UjY7y/YY/QBqeqHodkUHjDbJ1EkPK3F7iRnGNW5M2CzUcgqQ6jIaQ+HGYA8Fgt7
fAupDeWn2qa1ajN99EPVQBbOSxBud0mHNOvXeg+HvhwA008uGH2wTC81HK6QmgWpkB6NAO0mFAqN
I2ohb97RlEFbwScKn8HAnZHq6/IcjQ7N//SAWf1oQ+4Oc6cFf2n5FekMoPQTnuvHnuZ9dPTHd1Hv
LXc3z++FzqIRRNzXUUGxiWhMuehXFfpK5bFu26jp2HUTMvms8GPgfF2pvnRuMhuSu9kpSnZH9bpc
AAKRFduPtYUQvtUIf6UdmEHctUeE4OexjCIMsbyC68muAUVD8NPJibzGmN6IJd67w/Da2ZDUMVoj
hJb52kNqhqgUdPxMkXSNR4MlAmEBHUyPxTNto70GhZkDDKUiQ/2wgmeGlhi48kss0rp0hI5epge2
SwG9IBLSQ2DsANc9So/y5Yl8Rd4AN5glXLhPeWo5AtnZfnRH5D29IAst9tOxLA65rYUOEFksslYT
BlIkRpnSno7/cog7phQbTx+LCFZirPKbPDkZExO0VS98dmUOU0/Uw4fQWcuL/x6gEwEk064Cc0RJ
bGM/L+KdXDix/m7jAE1Usla1WfDASUX4bPqe3AeiEz/9llxu8h/MP/8vg5oA8jWmxjGpg1gMKkWO
b88Al/aRVqToAoxUxH7Z2Sav9Mu3V34yR2gcRFdK0kgrOXFSufbSUc1NxixceuYZmTrk7o+pO8RD
CuHcdXckGG2g9qELQoGV+5JigljtfK15HZnRXfjskMWlGZhEn3Pk5pqPO+abaaZjwPSL7xqW1RSC
L81tm1wqzVKB6na/LsQicF2sIdVU2GBDoUDwh/v9ehxXj3NaV34J4IlIC8Dt6oZLU0Aa3F8i8ila
Q5ohXelJa4ehPnB84I3S4lj/Zxoyz5t0sVGZIPxJktVS4j7Sz+y/oNAocS1JnJfWGFPRP/bknbVn
QCMwlUYX/CmQT5vaAi9izOkg6cuNs8UYdN6DKflkBR8jphlRzrmK+fYHrV5S7rmQeqAHzgtHrfZi
niuh2o9fVGmXL9vQcA9Vt2k4oUxXghIGEI6jlTsveTXGFrsd0DhPVersc5S84qB0xDWRIygiGusm
hP1w48bptMKvT6xXPpoaCQj9VNME8jSMCs1hKOyK85S/Qcb13zhJR0gzpQKOJvy180QAQ0iLeYry
rjphqiJ+Hh5rQ3NU4ZhT5MZc0qbaxEd+q3IXk0poeV6LPoKXT7X8mccvQ/zKIRnadsaqdRelaLqh
igOGbsf/bFRK8PiCF8Lun5C9syJAloz2yXmYmyUqk8sl0+CcLtZh5rJqxxfbchqFpH6jfBqCmt/x
L1fDILxreaBXhXzaIsTp9AQsbdyZSxIZTCUNMu995hepyLQHpsDv+xsBg3kp6vL5cHJUt7ce+8KF
Q6yea5AR7jQpvFHgaqqhfSKYMQx/2bS8CU8qhll8F5aTsoAXjBDNz/ujBV15//low7IyPRJ4nq3a
t8cqEa7nrEUTcW8A/wtOzzmutjM295HqCHuIgungowXN+bM8EjFThVKLjWI0psKkIVK/CLtWTzea
1M6vrbvRYEvBaYNP+cyXLwgc6zNTNowwbNdlghSwq4+cyX3yH98D7mcbB9ttSBVHVEfrt5qskI8y
ZTXQmeuQIVw3NaCv/nSJwjCN/DFxn1ogh7RCUXMiWiz7XY5YQ9Q8zo8afkuZinUaX/1wRTmnaTRW
phNhadDXkjcUVnMunUOVoZ8f6TQwt5X65VSGwXN125JS4HMErPDQ17hM+S8zt7mNpsob2eWkdRpc
TDGJ4PuVaoGPydAMtk4K2ZdkV/NB9ht1FIwss8vifuVHLuDYC2+8FUmRc/fpQV43RTsXcIX6VgHr
B/wblREK/P5qSstHui8SNfWMuFAOQYuEj6cD2Vtb1XJnSS+Kgr05DA4O78BlZrkTZaRkkp/fU/3S
1aj+BqS30xOC9Gy6ft42KFMZ/mkxEtoOha3ByRlXjAyvFX44czM4UoOBQqhGfneslf7kSX+XWTlc
IpM4g3MuAHvaykmSmdzHOuGNwCR9Wpdy2tnLwOKt3hq/UXcJRUiWVYPCyQ9KsXJD3iW5z95TXwYg
gN/QQMXou0PpPOz3GSlBLaAHv01u/bFjTC6SZkCScMoUSS+TwIBLC14s41HhirfKL2xXMUrXpC0o
90AaqcGXJaC8Co5HItPoMUTHqo7ig5b9uaTp20gggSwIgRA+3RNXXXXHf5nC79UD/hFnEkH7Pogb
q8yJ1x1arjL/mjdEoEPgs82aagYinRUEsBS4WXGSHzuf2yq0Z8C3VdcbWocroeAIuHbjDcprQ/QV
xM5aXGtpMnYtl1uhGHSaduJIfyECh6eH5T+tBG8xCS3wIX/zCEEmpk/hYFpFj1GPSlax2kyY4S/j
z8goTVtAT/ahPAJ4BM5wfMh4Jueh5kJQGu61BNsyrbpKykjf1dsCFYo/h5PhNwV9cp8Ljl8DLgfj
lt7wYNaiLYY7bFTqiaX8evUqwjV6VRep8wxzQVoAgLps1T5KVBU3BDAVLdo1dvftoHQE8kJn47yd
HEM+mlToj2i7NRScMjjTjVTEj+4gkCgMTahmk5T3RZhovoCypFKVypayOKfriKGiWKHm9SWNhd9m
yKjTimJxhPNkdgWTnCtsBV6+ujnEjH0hGX3VS/A74K3iatedUodpzR/8Wtehn3GPZcSgxY4HAkWP
72+gpZ8ZbxlaJeIvyHTZOyqzLTpnyI8de2XUsKMQXQvg84PKD0emublhIKR+/lddiDXhSG5lEweL
4+2Xd5ppdNCjpllg7bY3M4rkKbWiQ/BDN+VE2kkuIpyTaGPQY6Nj0PLhabw27NOBb4SaOUtNS03D
zf5JWFy3VnPQ0nWnNc7tr+ZFYHZdF+nHVNG4HKOp3M84mX+SDCkp6/pTzr9SAn7noHdc3bxIcSX9
0q6cvO4lznyby0kJAURFuVBbekgKKPN++1SXW59NmRrhuyeKa77fWGw2Qvl5b+3TJP82zVIUyCeH
HxfCevQLEgYH2Oo/wij1xzFGs0nXLqGz4C7u9rRWNXQJVuIEjIqY5P5diuSwpK2fcgJOztYWfwrE
fggn48ugpH53QtDFrExYOHMAQSYaViNaH4tPcPhW1koUjF3Wnmf4ocBKT4+cUEXuOBgLTkQICryf
oyk4/6TowOBzCsT4KkOz0dRlqJB0X4DTIaAGOZma3Ocoi02QzQ31beT2G6wq36xQ3BZPiDgy7imG
neYwXwhWxcBV9AA+UBiz2HEzKhz3Rtk/0ExQGX0RQQS3oprMmoxzco4FMO6hEJ0+vSc7BX0Rn3+k
teMfUVKBTkHO33FH98Um/MbsCVdwMqunmosRbMcacekhCoazahla+ryp482zN+GalhnLJeMRP17/
Ne04syxC4QfN2b75726hK1LleH3vKwQ4iifUVRnwEeOqYqk0dNd7yzF5s7E0UPwhBwRris/8hcN0
tALc3vQkxUBfjm+J0dm/aFPUft/xB/Ozl23ZZOfYNvFoxmT2xYxlIydv91u/+eEaavtsXSNDrhHw
5KUQNK7+cl90idE2TRyUMIDoYsgC5M2nnSX1G/80bvlCa725x3lFdGTsPxQZgZgy7AZxzOtSDGvI
Bp6zcSwZeHfx5HRdVNsOR2veHFP51yaAyc7wSXTzM+bfFRfOQasNobCwSPbnLoUeUpGwtxXcLYAh
EmmrCCOJkAdH8jaPz/e4fJddIoCEPhYsMzBIpWG8qFac9ZEQHUjfw8rfKyFy6yWFonjeiIWN6BNI
6vEb+pQR2iZpaULVAstdyUf7B0IEb49Sq3rJSf5QjDVNPGPBdDph1xBqHFUfE/OuQZKzooC37eQY
zWTRQ+aOYxt3fMoyCpXAwvKUIJ/G6wbZG4PIxKzLo1Z4EFXmLGMF5GoWv+b6WhhQIyoCeZlyInuS
lFPbbYJ7H6QuuYzZTqlhV/bGT6alsHELkVI9zGCkZDdGMrU37eJYjHJQlMjhIieo3Byyqq4FP6na
S7qRtr05yYRa8CTes3yXOUC6vLLbxWnVJ8ZOu/u0c/QU4LAe3CY1D6TP1rKRElit36xG53oSmaeA
WQDmquc9Weaz1BWOXH6YEDOeqUABsJV9Q/gLBCIvvsWnV8XU0PlImqJ466r1y4oT4QY4ZjXKDWtH
M/Bx5BqEJulIKfI7ENGeunT/7N8Zh6dhyHK6ef3yrlEVCWw5pGZb3XFRp4JwtdvPNO3T+OAYCO2V
B9q81qPifB7+yFQmOsyE7kUIhfl5Gx7nWu9D+KNu8hmKcWlgqMFRjNRC/OThsmN1Ceo2huH/UN+h
kP75kKL6pxEZTPDfb69F/qnVOQjEKyorb3qVKwwCYA447Uh2ZS2EZFZLC773eYYDZvh/AAvA2T5h
+1Fg3v3+Xlnj4+VCOgjgy4f8ULMgE7ZnYTrds9d84sXL56SiuO4aPpjk1dGm+ORKulnTwn8o+VZN
kMvKGXePv3YXfj8T7MxcVA74oaz6UO5H2F7sC/5NmgQVYkvLS43XSFI8R1hNT7V05qZ6Cfo+UlyS
U7V1Fkb+t29UWbqNr6qk5clcJvtDOVyfcaZ6clyEeoI7UJc4A+YNELBLNBdrx2su+vcS/3gr5zPd
uwFy9fhNuB9IarZxSLM4vF6THLrck7I5N0BHkp0Dchhbx5qX+YMPZWsXJhhSFw4fprKJ/DvJPaXv
iXRRUQnfVQUqW3cuV0i/sXHRr/0ErrtooZG2/RwPZqN/qLe6rFUh4C+UKbyw6668KZtX2UvbVjHJ
pme6+EAG9ewk6XidA8OF658S9zBZ/f/BORtuuWnkwvDAUCI1eqlaLHQiP/SjsVRA94hCotMC3Pae
kEAiTiRZBY4fLOySaDkcMHYlf8nei1/whvUN/NoJyww4CbzPdKyZ93B4FA72bHBIxvCANQ9p7uNc
Z1xlbA3HSG03vU1W9N/3PiPiVicPtECKo2pYOZdkByjrjLXgKmmIm2XNXfXQvogvYpkW88/xpMWH
VLU5f1z1PrA8En27pKi0BLzuZ2/HkQAJrflh5Eb6QBAgaP86GZzgXKeIJ4FXDX/Ek8cesAssZgS+
hREt47EOFdIyGyk3zpjB1wkCXMHS2J9SixxbvYtbyl48rAnezbtIqt6HcDc8sBi4p7Yxr/JDa+on
Fix8dtBPCc8fAyg33Nbm4KUi/ZFY7qx+7Xju888Nri95ndHeWRrCo1Bucr9haMFqK8ObLNzAjpOl
D9MGzl5WPbcykurEFV5aFFXSmdiT4hYhXZg9bDL8cXy8Bs/nOanMtgotqPlB9CNIsIt60lamjCzs
FhF0HdtzMyRoISkPOUYlqzm3Gru1sJ1lUlyzRwSMC5nYO4pT+RDQD+ZO6b7cVICB5boQpTXstzeA
OV92lHx5GqrzXAG4ccGbEWDLxAEkW1ummEwW+n6wQdy0NJRfV7Jd3qweK0jYNec0tQ+RiyJaFAem
BIv0hMQVV6RfDVaQ7SQV9s2cLGKEwzCeznEG66l/Eh5VQboYlokAKZ7XiXZpEzSqXI1xZQ6DtI6t
Spx64wvcmnPDzW0R3rl4QGXr1OkDOYQ00mu/y9Ys/Zzt9XF6Puu2EyyWsBjo5YHtH90J/8nRntqI
WSHrF2YvIoLYxLCiKshdOmFNT0DzkRvuTnvj1nWmHT705jG2xGM7G9bF4gF5WlZatJxpOEC34FVE
zI1+bnKjV+qkmbSCj9kxGvMlAvXu6nL8fqwayYRMJGqO5CABPsOOY049/59YhFX93RxzW6Ht9Sgn
R9+9JZOgNgV7G8deEBmRgg9LzvV/qD/eDL1YCZkK3V06qxfU8jiHJB456blojhij94zUn0A4YXot
nRHfHj0j0fOdDLhlac4n7NlXGjkspwA1c4lpmAlcLzPoEb3dWyvBMQsw1yxixhUEBMJIhK1Kng+W
T0Mt6AbhGj6S8+jEInD3MiGUighGvCWo8nb7k1oyKuY/2ZfJiPqfLPWTjVG2o55XgunycKPwx6IV
PWgZjSxPSaKUyEBGvFn1Znw6J3OqxKfOX2e7cYTLKPPpOVOtKtGN9IFjVW1Kv33BnEDxpCQBtsWB
z6nnEcA8dmwPbbrycEkHQ6F74ZbpUtg68LIeR9CAymYR29E9mmF6DB487ziKk8HALQrVkPFzC2f+
gsxUgxC7qU8Z+1bx9/x1R3GxxQ+U4CkHB1u6gcwXGQQwAVJSALSQ6QfQ2NnuI9r3l/jEgRD7v0pS
U8mR5YHCql4xUXTFWJrXVr3Qaxt4EKDxNGpt2gk3nEoV246zfdU9GDxzo2nVVnti+/+iGEuIohkn
7OLHTBsBoUaQJoZ2fxEEOYb0Hl9CsOiaBpKs/Hc7nmaIPtONYnA2jFPRnfPvCQBRQtV2Y1DXsG2n
B/Nj2BFfkB1zEKHW4IWOV5gOsEHl/sAVuvNAyTYNhu45S99yBTWVKbxBl/Nr7r8pcJVWfFIXslhG
BquEpORoRFsITFzjrA+YOj1vd9jkhmOxZA1jQzjoKQo0KbAi/a+E6hkDV6HfxvaX9E7L0H6UlxwY
RFsV3oHGwqfxSPIl1Zhuu1jSHDGwliJNbth9Uz4Bl5THLeL5pLffcESWyXhq2WLYf1VWkER/qyRy
qEMFXuqGlYTh2mkIcJ9XZ/C6R6PZ7zv810/ogtxSnh3dTEk/za6D7exSSSYSbskvyg69yEpvTHKL
PTZBVo9g7JdLRbRcqUhNOFhC3F4DcwoY26A1LWHWmgGbJ2KbjNobPac4gM0ncsKxay6llxr7tl6I
5BffIsKzBbt46z2lwSnU4GL92yXU6le7goSL+ric9JiXFDuaaZguBOsu7yAqzgJODrKHgqmdAUdW
BJOhCdWCrDG54wVVGIJ2yx+996t2PTsdkNFHp3uv/N6LIvtGw3wP5hG5ayNMjRal2cdCMvSy65qB
hIeFUY2U1/ziAvPWNGOWSgyaotDdNOodNiaJEwm9iReLWgogQM9Y+x7z9MUuhYDefJLGokWmOQt3
39wvH/jZgOJutQEbDyYKnD12xr/uwxQrLYDFo0WsyuLziuwyVyk98CT2++m941JjLVgSGuwWpfaU
Zl3rx2J0FFq2AQwT74xpZ3QOmwFlatS402iexzmmHpe9j3lqq9To8xIREzwTvcMW4GKyZMn/+MPW
o4uZ/qcDO8I8fZ7az+TqFBBrf1aThaPtxwjLrIgV+n/byzhSWBUB1QXgH8QdFVu+UO2QWAIvbW8l
0LuxW0MBnJQzyRS+VzQubQmfuq1RpuBlLJQlbQwqai9+uMOzc1FG7+5V7PqMjZt+YGnOhNUJ4W/U
tVnRrlZ+/G5fBp2ezwe0asBPUsbwDk21AVbiPRSfTz1KlnL//Zw9ft9Zs83vi+R0Gsak9y6AGHcZ
GXeGSFQDCdvrtFG41Do6JUXUT3MGVNFhbq7HIDFvMQtOlgqAPKEWho3791+CtC4YYShexeacdKAu
Ky1+siXDlgDSDrRcIr44qtqGZ/wpMQjaY4pj0T066QcX1VjhcSvVBsPp4JY2TBnqN+Q1jiPfclqz
ojqilbXTJcJDIoyXG9rtNbRbN4lhfBGsNpGPNICrSbbnE1L2gR1ouQE23GBGle5H0P0xTDas7bWe
qOcxZtoNUF2FzEKMjHU9OQ1RN7daHzjXO2xvRhu4dX+quD+0oIvmptrGB9i+gwpbutlEQ7P1AOnu
NE4Z9S9AGeVgfrl8LpXPnUVbHCl5QFDxFPSXEtmLxYXnj3YgEUi0kLPzb5QOP698h6QCN6oq5qcD
qkilkSTrs+BD8BzqOCAb14280vd8cHu+XULDU8o3v1XyIaRx5KfFfZCbrcW1QmRmaK5Nl2bx1I1X
d0+px5nJAOLTSz7Cj31x30tpHcSItceXsKgCbtrGjGmadVFlyHkaejVwrF4iEh5j8+TqAl2BzPxl
uh5RbnvDgWR8T/sZjH9Dm7ih7wuxtK+uh4wsaGZN1jnZybFMHa7WePEuEwnq9Ywv4Gn4OeNhvwtF
4yQ7RIn0N36qEdkQ7/D3mYku/q/TL2ibyISvNk//iuegF2lLr7bDXllra2R0/EvmeZqxe3YvHmzG
am/mThiXH13BGXyG/sdeXZFyIh/FyHm02QS0qNNZXbdqC2Fqw8aGhxx8nMIcZt1UVyiIstQrl1ct
zv6fVRSqc9/okzrZmp3wE/1g7gM1LHKMv8cEcYkeKaPtlpmJnGrxHyn8OL49kBHmbr7pDYJsRJEU
nxZj4rDXJD0GFuVLVCsEhkZVEI0/nXn7X9i9LG2XtN1BGn9QCp2wNpnl5nv/2MS1702RYX6GvlMF
J3CUE+vnMP5+oz/UxN3Tuu4xk5c2C65smx9Azm0drCvVIYECQBnxq6LPc1SuWAMVOEyKvCW//zmM
hQ0/r28NgkcbOxxlj+NOq6CuD9T2AbekVwChSGB2FAmEd1tHrWWceP5iP3EFuYKRnl3ubQbXlKRm
honchlMnZsDGYyjXPC8ktZCkxq8w+o3uZmSDBgyiZTaQngPwvi9YsZROYZgYXZb52EzQyFZpHg6T
ZxMXNe7yssvja5hY8OeWxhmVMYOqiLHLrmLb1eQNSNxzkH4apBdg5iOfsvlGpppkROqQtVm16oG9
/mm2U8cI35VZVxFQXeqOfAoyIwEgX4tggz+m0oPqOCqKDLZ3VxuofToxXOvRqoLeFunurUGQZD88
Irps16Q7lgwIXmKjjet/uxBdxTj87Ryk6GEXWSOGx5HaAvrs7grp8ELIA9rvtfO8yJZajnVz/Cjo
gc8rlexZYLRll57GUAlGJxGnAdp0Kqpxym9L8iNlx2eJJrx0Di/kkOuhETyQn4ONVuXIVsBbMWfI
wkNi044weayP6dPN376pUlO9nC+AwBItMUZ1pspBq2FlQg2S4FYCcuR/8SFseDUnnCgmON4Ed4VB
t6+jdUEaB7dJjcI/WNqdjM0YaUzATcAs4Xo9KdqGgTe6HXdczDFUCX+ziHCbxs9nA4M7pa8kzEHw
yIQV42ROn4/qA0YJNucTm4W7qFPAK0GUeIBW43eluCott8AA03SsffwhPmmd9ouCshTaeMEQGvRj
yjCOx2+vNO0fjIt4Rc8PItbP4woEZzxZ1BJsqxv3WnFWT7k4mkoOwbbqnwXaHe+xdvydwVBXcvzP
bd/W8brMtcwRrbJVByDHW6Undtt6IGDnmsCnujTiFZxmFYBKzqZ+pMFCmSZzTqXtZsyd0vP9QGqg
wdYaGFB+or4p8vY3lNqiMXNh8cFGYt2ts1/m2Z59FdDzu+iQ8Goap8chclNB0eXTtC5RwSd/5Y+o
kFLG2X4dtA/kkfaJ2M63/h9R0OWGppw/w9Mh4oKOE1e4Ry5H0NraCe/2CNZfWcBRIsT3Sz1X30nl
IggodNRJOCEs5WfyYMjH6ohLqbyXtNTxFK0j/t/KogbA8E1LojzRFtCtTB+GXpNTLWn8UANuTHHT
Q/g9xRWffjq8VC6SkCAlsIN7obtWsgFm0j2lS7VsXTK5KmCbGpG9vivJpEKC5zHdZMfuivQw/gdo
XzEM4a82oOVG1jeMXHvWDpGZQO2z62TOC3RQN2kiUMTiMv0+9ecUWBx/qIWtR6DAXPMGEvSQqHfQ
XNqynl/XHRYoxn9HcLD1BtbK+aJu4DtC5Nl6Ol+oFFY0hRhCvv5ftEFFlArkEuuuyTtINH6WVLzX
yO8jmtmYRNzjP5DLivZCc4PS8S4N8gRTUkA0sOeHwPs2GKWcS129O4Kl+G5SyhXl6KanDihjkP6g
shA5RbwHKxUC8Vz6joLVunT9RrmxjnX7WdrnrF9HcrU3wMed2TAlc086HY+Q+699EOfJBVoUgz/c
/qtpIavqbbyicJIGCOSJjK94FeDeLKmwwx8SDNreJ5NaG7dcfCqBpE1ku/qSr+FBf7phG5H0O6tP
+AwpyUPiTWEpQaHdlK2Q03Bhd2WS2FCN4Dp9iKij+bb2V8ERaTR0V1O+TugzscIQ8wkPHRy5iD7h
WNi8UvYadUdmyA2P+9zTmvqE6Nz9PAjcC22QoJGRP4Iof1HmkYuiznBH1DWvay5NPHBpHzJuBv/N
rDAzB8g+pkWsCAn8BgJ0MkfkNUefXAH8QTv3IgPZe8ZTRRQ6+5crAGOZPgXr03JDCiBu220R+1Zi
Ra3OlAE9qb3V7tNbZCR8wzLd8mSo6xEOVg/NtNMX5WzLyEJx6M1ek9Zkgm4eW2nWIBEE/NI/o4vD
CLFlz0Uwx28HsvoAbzwCHGFRq6FX5sf95+XlVwQ1ULtkWI3byWfxICNOer9+wjrFyWumEykKK1ro
1Cj32RYe03Q9VRTMkJiAlFhQg+/Pw9Lf5ytz6zLeBgQDKDwCBZUMgo+EIjmgW47ne1PuiAKBVKV6
vhaFm+0WFWdRf3jj/xjMqq2ySnS/aZVubqTKWS94mp8B3pqTWVmbkHa8DamYUFVJDZMYLYc4QsbG
BlMb7A5IgL2FN9PafUKvrMIX/KgrEqM0sbL1b0/K8R8mi10K6epJAEBMEKjoLRVTedWCxc+UIdw9
zj//gPGwaO7qb9VwT1Pdq3i8Y6h/NKahoUMWMbWaomD2fjpLqig76wUTIQE2INytyUl7GWJklKcB
uWH0H5L2GH5dpVJFTxLF6KlPDeg3LFZKuopGmR5EIZJc0VAFeSApRJ05zWU/uQn6ohpbAihMaqEX
cGHn9Uc8EImZ5ojU0NjZ+TKIaMS/U9t/1o7nnGDOB1gEzoh3zcKzmw1/wgWiXc4I/esFZXl939tk
mICdPQQnHzqFrJ0p9c16/KZEp1KV7P5nrswYMWMSmo1QHjCcqGlkYpGBxvC2WVD7wAlUydmiY6Cr
DaICOUAmeZSiiQYfxVV3qoGb3PrAGlwwFg4Dmca+W/lq9XxJT8514oNK/HdgCJK6Fyh998D1nTLy
xZOZX37DOrmcrVPd5RHr9ZCBDNLjadW4qXmDjdpZynbo/yIXhHJuji1ov9o5ACd1FmMIAbcbETwk
jVhfTtVr9921l8pqTlpBaGgrKD2wA56yWBCasPmti8mSqtQScXhpERqCyQUUqZspzHqTI5UHd1T/
a+/pUvZgQ9iLu82l6WtDMHCRRvJSIJN/SlY0uGOqXuaHaAgF9XneDQ/zsDkb5adgr2gzhmZjcmw1
trBnvWkQkBJAqHqrzqXXko9SJ0dUwaUZmrf+kFWpcf4n1QOPNrQocickJrzwguch+ZF2S7YmtrlX
YOyhjdDCFBBws//acyK84WgHh3dsGOqxCJonxUC4c7nyg+t4Lkv8GoTkQ4q+noXe/GU3RLbtYQIm
flGYcnkW6g6+e+lF7TvjqXMNimgoF6un7rS5hdHvD+oCQVzDF8tLT6JKoK4M5EVQenMrXg8/fpYJ
G8Uh20yAGUwrINF9JQeYrlxDkbOnnrcmo+g1wBgWFEkAQ9ykmpyzf6BL6CGxwCmLvOYpLfwYbIu2
KuuMNX/KZl6XLdDK1s6xAYl4d0MMsXVXLBw/2GBIj6B0/Jp4pEwqLk+8X4Di19HHxx8cf3sfdZ9i
8ZlrCK1FBTh9BaXcu1Ox2NK0cRr31pWxSVLO0/SCoOJd5+c/Zm2suH6wPoh9Ktw0SAviXgz/D/bY
188M8N6CEuNXY/Atnd9gd6bYzBhspDNnjbFb0IPnsrrZZmqaLru8Zc1vI5BZnuQ3tQzF1JZ/vVpQ
ntX98lxsRbMYR4N5vKe4/lziNlpnNTwAmDRJK4yVbpMp725zZ6vXKD8R2DE6ks9xm3JgKBMTqBP3
AEKX7fqyNiJJV6mLtrKUNjzJT4nzCksQwYDQKbanhtYFYw947L77RUYORS8t4dQ37LBqE4cOPhGK
QfmkPdNIkx1BWVv+6LXDxlLWjUrqN8sawbrr77iCkMCLUNhidSCqKE4KvPqF6IOcvJLgPhdbtZvC
JfrmpL3scV2oUT998R5kZwhEZtGfC+yMZIbKWM50Y7pri669EE6YiG0OTrxJFa+c1QTTy/eh2s1J
iy/W5wDPQds/rPUxUDOkZ6ftdGlMBQwW9w1oyeLmZNLceC/Gd7a6TKicpJhSzhQyMSH3rEZ//B8D
GjGLgB1dUgzn6QCSWUqEqHiSf6kNabQtORD5ZTGSpwSp9wu1pMs4XYrOsN79SPRgmQVNz0wDYxjX
zjvjKUGo3UA/Nn6/9KfiZ4SEWRGJdms3QSIHu2g/HyrwKiFN97l/SJKLqV+eqNEN6H9keGU9T/4p
XZq3gdGR09drWahMxPjgCsVYplcOrLfpWMVKykmCdAFp8+guloM8NlGJBrbJvnmEW3NwxVIs/1aE
02T5z4NKzoHhMrKE9gXTn1Ubvo2sNBqEl0uvpeAAwWlNVPet47sZ/K5r+T9VRa/r3MnFDlWlNxuK
zAnnTU7Hkm6FXHcCXqbxtKC1Qxz8i2ZbKk6N/DQwm6s5003gJ+q7zVsa0ibSFLuc9v0W12fFS7YQ
VJi6MgFLoZlnlhVIyt/SVh7ByBsEkd0JQnCJZHlsscdCZHDlvQ+PlSGJ/trni4Ftiu9873ekUK3Q
ki+Is2Q4UE9Iak5pXLqqDL2DXt/xOxNuMWG/K+BkAKF+yu2Gm/S4cRoARHdo9URFswNiZRjcVmQY
bFwdfBubjSTp66gMn/MPzAdmZ4LjFCEM0rRkgvGaspThhD2tT2M4Vf7bmFEtgPtGTjY/CNVBgmdn
JP9VI2o51nhJ4p9G73QScYZYmOqyTXbu91rHy3rjYDeyfwM/w/cY5eFzRJBPwMLjz/kixTJQgOuV
tDMAURguD59HxliggyAaUUNPQxurHx2CO2ypKR1CXSBJXDeXshWEMNjNl5IhziAIkefANdkwByqP
24w4n5B3vx1Hv90h14IRqm4Q3M04Plf/a6jpdyhlrRrv4al/i69Q6hxMVI2oR8PHsEVzsKQF8S27
EAZuxBlp991gW8+eCZEqVVXLSYkCz0w3+D3jgL/VcfKE5BAqzahzNubMayjDv9hXfVuHhQ2OaRBU
rT/K65SBqAolUKO7AAvi1t5qcyZW+FRefXNyyVubBfGQfUXNkk1zbKJkpm3ckqDh8817Y2DnZSzu
J+9YdDKX1FCz4MkzoVXVuEMEtmFQxhFkHn8oykLtqcVfmJpoIrh2lxjQ9IN9x2q0POqPnNoz4+4t
KMN1qLHDauTsu3X+YBPuJVKMConXlZ90q3W8+T4jhDldkeWljoabH9u5q9H9SyJzYD+rOV0Acniw
V+HU0ul9ckeKM/O7kpBaIbfp2fowJmvghqnXtPG4ZH3JzK0CTRpTv8SjwzsIZt1xKGyReY5Nlmsp
2bciqFGcftA0DZvOzYdyc5uzJwyDrvaCSvUBX1fAjR2uxpWY6J+DxQ98Njk9KD2N2SJvrCiXmbzb
cN1ng/VK/neHVLilWD1GPdw51gL6f0RHvLtm3L9KjNMUKQxmTajW+pVUWIRX60UN21ZcECxkJiZ/
y1ioEOgbTFonWZQeD8CB/Zeajp3SBsJwL0BcxfyD4kmzVx6JQKLr+DEMbOsYiq1MyD7OKUMJPf7F
Lmxv4o8HBK8r2wAgKvVoT19plIme4ssgUDYQsz1kuDrVa0+7aiy2WMN8seaww0LNpUcdEwydtRvF
FAKUA3RWXLXCZpaPDAgkG7boaX3OcJVXfZa+7k9pxfUQ/37SDkqEmRE8/ZlDJG0Bbc9i7BLDgB6O
7jvrPEQQd5IWf8mHeNvZNZ+oGOOrR8XdBxddkkfVfJuRuvjXHCXH+80HDvzg61V9+9Cu6K3xd46m
K0oeegMGDFdoGZRHZpsFBppXydsAtI20bQ7ZlIxKlvp25q3JW8LZOrszYgBsqhgpPShCjX/BtWsI
MT09vJtBP65hMnjCKsUMbkwF2yYWeSSY5jdDjmPhJDLtryVJo4t6oqKvbkmaJ5ZggTrlyn/tF3rz
AnO0qAQPwOvZnhxGLbwYZf9b1mdR3Yh1PzF6e7SFkIaBpJENYQb+xo3QrAR+G7PI7LpQ20c2ncok
16J3dHN35z2mxk084KqN4vfRTJiIy+PjgLu4wvGWpoupTZgrFpNIkYU/dKHjz/Slv6m1VMv8Trr+
is9HfQo5TmVUHx8OKDTg7p/Or1S2ML7nMRyIQZ6tXIeLhkQKEG3gNBGRWfyqejVe83BRDE8B5XIA
HjDeL2GegaZHQKowXRo++CjVZ/F0ZYKkFxCUE+HoL7JqtKQA+2tVhJ+rPpItrwGsrobFDFLgy7kl
p/zVw8bJVKfVNDo6i27OmnmaJ6UTEN6bb7ovrXIwgxba6YwawwKaGcV5qvcrlqD3poyfWMHn1xXx
0xFjtiX2ilq6VztGRsvLRO7E37G3Hl8cBm1XWPpEjHOLJXUO0oaEE3Yhzlg9LBtQFL0RQu20FMkE
6Qqf5aUvwqLkMhCP3LPQdMwp7z4yVpN9I5cM0dwsgMamfXjLF6MVCecMElfnCSIhm+md00cRC6Zg
CqJTqCCmzmiqCyUbOQx47YeRUM9KWY1omRL241uyWvWozjGDtoflZY+gycvD1mKHM4rXRk0RyAtP
Popq4xOzoGMZiMgfJkyr4HqwdCReeY+krb9QW+uEbz+qjGI9FwvlHuHU1THjaolGsL96dQa7AZy2
CobkUolaoyEkw3aYjDkAGFr60qiktQ6WtXwLXEJ+Lq1x0MrRQzbp4UxXuOUR0j97ehcWsSRA1Gv4
vtCVQdUuGr+O4IlLtMlrug53PuAKwSCt/oIwWttBGLbmE+awaDQqA8t1ZvezLirQ/IQMWJxuZXdz
ypBBMaMOxHQ6Vlt2yaLPnf8SO0MjOVX9dyUANAyspms5xQYiUMa5bETmTGK/Jbnb2HU3eYSM61YM
ewk7QSLavxzYF/NgsaYyTnGmw9jHK+4p/8jvZTYlJMQJqi1pLomtkuYIIMfleMMvoBKjFzEqEp+E
k777LZB4boDTIICtaU+x1DXu2p38gvH8vKVRRxqOqbfkMzQi02SSmroynn9hOlL9tgPboAXuV1Qy
Xd3+CyWtVqYazKfXZGpnUFSbro+dN202YPa/nMdau8WDVdMIP3lDsN5xBO0ClwibiTv6J/fs6tuH
BatsbdmswuHB5VQydp7gxGdZJtCLV+goo2F1ZDdspvk83hFFtnAd5i1QHUXq4WSh1vbxfZNSyPYo
dvu7ktNlq0lvNJK/FdfRujM4Ccm1+pr0FnM/MbT7TTxIKjHKzxDJX+H/IACxlCUGe4s5okm3amlj
YXZEzyhooma2bmx+iEswQNpLn96nhVMBr6NTtPle1xjRxVtT9uNPdCMuMZghv5TH28AeSsEHmkTK
tICqkcwMqehuDB8XBFEFD+OfMHcfSpmNHlwidspAaJE64mlXzthtmY0wJJv/a+PEwix1A5dTFRuT
+Hz7mLe/R+wvCzieJHM27q0WghR+nmgHt/O3Bs+HO0sSAIiSsE469kXhyV+zK5sCbKZE5O+KnXVF
vI//kgE/gaYZtD+vIigi7OvhV43HO6KlT5CWaY2YOh8mWlS1MQdwR8CJGWWAadblGq4PX09F4jQs
D7xLIupCurgffrbbpByb4C4ViLSUiIvCmsB8nxTpzOq8iZ1NGL5DfjFnPUgmuWujt6jr4ptxPBhN
9UpvbshHdFdzO+xtACU+Tvq2mPHYTl6dDL0myEs/5PS59xyHCw6SmGWZwMQ+Gr0/G+rZSOAEN3qk
gUeGGtN2mg1BjWdP3PTKhsrN6ItUsup9+RmcBwcm+2LTwNqHAHgeYmzJ/J4Bk2s5uAQx8cmdHeSq
/X/1D/NfV0U92h0BdYv2bk4gR7kopc5zovKgM/5XPlCWmD4S8/uy314N3zvv0+SeAgTwHAqOT45z
WwrppHvjxGQSCsShEe6YUxBgpYJmejdiHI9kn52EMhZ3k4hm6c8qanNwtdxGLjbaZtX0F/N9t0e9
KFZ+EwOm+9dO1sI3KMuoqqFPShtiLAiRRhwilnkqnZ5Iivrr4WpSw5J5cLI0jLtKlksvXxE/irGZ
2UsBrYo9y2HQcUrJXnOHaEJnd9dWKe+bXYL2P07gUKLUzDjBh2zAHTW3vsRy7r3dePBZ5zb80D3M
V4/p2q3pfusy1SOD+JscKPUAw0aTf3Nno04+XptnPA1DCy6p+fLe3kiyVBhA6SS8apPDbxSbYnXR
ta7SEjVYY1NJsiNr4hKjAlaGJIxjkT4R8Wj1d7I3DxY21NpYhX8rGyNRl6sp8NEQLJGt+P6E0eFr
/t8nRAM5UTfHkFckzSSmwt5nFvgaRlGVIB5ZTEXzcn+yA7NGFj/ayxXgTjOeYRU5cczZNXtVU3j8
rvqwGG7P0Jjc+Mgw1QJxrBpVh0y+k09YUZr0kEeS4w/Air0PNUh9yDIuQ/wU338hDb/x42KtjK09
51p6piuKirECdz3M9WHXnNnn2sC/2GPdYIw6HqeTVDG+qmXBjtOZ48fVei2TmcRh4m2hdaTrdNUs
ksO5lxrdzVEoa1orrLGSC3xcwHkuvzpa2KhW8t/OrMFNR4bSzqsOeW+/p8LQl5A1A+CguDQpCJR+
oXIlWs5EnCbdqHC1hSDzLb6xRAR6ocpNLK9SUkc7ry/3sT0MEd/MQEreUXYtD9+GZFF/nBdDP2Is
ixVUqRQzVDFq6pL+pjLu4SJpol7y4h32s6xBRC332Vrv7X1NFOi9Ae+ii9x26k11fqC57f75ztC/
UeVcKFSvWnAODXIb8n9n9TUWvBAB8yhL7YzA4iZPE/kckyMKhuZELAqPMSsAP1hfU7YhY56lRf6k
867qdy1cUDi6X2+9Vk+zuLFQPhfopOIb+0cDfxyXncbvea4zSqraXVziWLgFCk3SNGOcCPONmBDf
I35kJy4oEPq8IKUvmz4Db2lrraAD83kWGsks04RLvAvrKeZXHNQzYpMpugBBodbsQVnyl64D28b3
k1izNURNQru6oJpj4h/m9aru4CbSHfynfzcUS53TljmJZoSFB1wenU7rS3Ci32PxZssq89jfZuFd
sD/XnVFTlFlpyNZZ2GU3yEfsPkGJOVdqrHmlaJ4JHnsxS0EvZWKNZNpbOZgaSvf8sLsWMXrX26NY
qurmi/J9oa++lhpxkgxGb5AnSArLxuI4ToEEjElCSVY1cj87n3npj2hzCP1/yLQTKdreXzISVeIh
nqHbA9OQfEB+UIjVkHyAR/8S3FFEj7C33KjHBtCzBUQPTAmNo1qkU+SDnLDUu6StqPVXin22C6T/
VbCU1ilrRqtZZ5WRFehhKGktjlVGpC939F+AwbE5V26+T6nes2fmHIJCliqLrOZ5NBGB9v0pj/ZZ
nIyJxOE98tl2f6Ait4KofosPRub235QgtjEjkxLwNkA/ykosR5ma0Y26x2WM3213CNc2g6nSZdQ7
oTxf3ok+5kv3dTPsA8jjfoK+BOzjFiUcbDxjx5/GADe3f8hFsf0j4GMRxIbJXU8mWqGw8WWihDaQ
QqjJEzoI2bmi65Jfp0Tam14ZK6A/Th1O9r4tv61RhGs8+MjnP/vwqYyP03qbFEty0y9gDxjp1jp/
4qXWsdnSSmpWs18byXWzYwRoiRwQdsSqERiNPIJofJomvNKI5pUhkFkNaum0SUiu5i0OJpDPNLqy
6K07a1+F5ZYEayxsckMZ4oOctiKHbpRua3bOjDjz5BG5jPzL3wwTb7tfUBk+uuxfVweGrz3GtT4V
nYIF4i1gHL1AObb8fBBg7d23hMkUJw2pDRhrn32q/R15jbTjSDcp62W7a+TRbyRTjiiokbzMYbkq
NuGexDxiejK2oB+yYDZZVhaGwjFmY4KW22gZ0ThLzrQId+BXiyJauL7dusS487/bSPK3fzORLxJJ
itQjw4hI7inxlvgJpyotbcZKbHptKGCF8sJpggYSsbvr44yTluFGBFQlIHnwplFsK+1y8eazkwHH
O+ZnDAYMA6GANOGdr2uhtjEG1KYbCIJbdmyCHWxlNbu+QbvBVFKHuinJ0qwarDZvWsW252VwemBg
Da5Zb6gDwZdWxqduVIeZPGaz4BMHDx3ESBFqqJUUv631IOSZGQPtFP6C47l4IFNdl958GACD19hb
UE8lUbv7vIM64Y961E3xUm2uWlI0+Ze1R9712yCAWq1k6i5+Txnr58pUivNG2odzXdQV2Um95Z4t
oYQ7mZElrN0xbFo+JlsjkGgMaY2KT/tq4WIarrNaRu2zlcI3KUvAv+YN5UepWZg/g4FYTyluIEOl
3vsRi3QaX8HtkLEupRmsqOzXiqVzEwvxZgE9BOZHfqLxmdIPVEFRMLY5ICjuYzG7nvS+yB/CxJ95
naxm3HUGMrY8x4HUjO09E6TniEQBpls0tlq9G5169TV9pECQEucohvhmbnV6OrcUVB1qVe2LRgjf
vlAGc2QrI7tKo1YdEhmy0Sj4fc3wz9rTMtvGSKi4IGpCRki4UDcEgPFOiSyrMDS9Zmii3jRuKGLi
76tcUCXrp0KfhG2gg7A2jz+WQ5TjZCsUz1y1irfeji/kgrfOxxHr0obgMwsrCgrcI2bUF9uFTkSU
1U/vJbnLMBjuX2qa2Fq/oHppcLGLABkykL1E+iXsS3vVh03MHgtVtLb3Lt7fG+Eb8/cgzEmE5qoc
oLvJzX08l9SlX/daLc4z5C8B0ZjAUlQiniEmEtlIa+i5EuRvk6wACHqV/pVfn56pmQOLfc43NNfq
RfONi5GKNiyFvPhRQwTV3U+Jlu8WCHdQA6jDyVvDI3b+aSlZw0UPLaiyia2MRkc1K2UM20gpWwQT
p5PzHf7jZi3Ps2FPJRWH4YElZFnEy+smQAsnIadCyecEKiLUq0z5ylF+kCdAy+j/VfQS8dIQBDqQ
ZT6OoJaUhCK3X/1sz6Yk3ODQyVsANd2yaeH48ik2jXsb2Fqh89IZmRJS7N+raUYKTOjyYzFfy/nA
Yao9/YTaQG3KktQZlVg/38H0Bo7v9/rCWlD8JL4LAaFNZvT53Rs3fvlePlLqFXJ1QLuBkPulRX+i
bO/niVijhnGzpfToEUwZ7Nw7YVmKUWyAjOY/KascUZM7VYulgljNsVZ/O869XlASOdkLXcZOUqZB
h73ZURKjajc1X7mJcqBgi/LZxc4RDZHVyOkQwdaaNRus21GyeHqvBHvyiUbDelvmYh8F6wNI0Z7y
qiEKfbDhvu8FwHBPKxJKg5G12KRL34HR61UMbyhRdV7MiFx/mWaQWobzF+zqro6MU3iFks6LzGzL
UlZtzf/272Qmgnvae++U6qkw4P326GKznKoT6a+bDMcl95gHWAtmh3fKqK0baCEjOi1GIlDBH4YI
R5HyzZYsfM/tdzWn7pvQIwAoPbXLpCq7IHN6+QZNdLUUDSAP1jU9sH7GpuXXjzd2L0XGcWfnBndJ
3marf9/94xdqZAxndhsR6y7yFddSarP2HB2pOhAMD9zgJg1HkXXhW2YfMdtVds28h9v5ABURHf4Y
sGO99QcMiyeOp33xinznqI84EY1PTgMNo6wVJU4j7uA3ecOK31B81diqd/j6KAyStomCNVSlYdL2
1QFEjxHNPI1pNlTbo0e12G5d3N9B44nIgBsrKDFlPC6Tv2HB0wQAWHkTChKzUIcolAq10vD5LqJz
12Fp7t221kB5aGV0KTSQBu8ysvQ9vfq11o4dT3DpmpDVmIiQ/yJFY1QX6bpkP6k2gbWAHFILr9Gf
i9lBbhKoBqdQvZSs/AYybkNwchcOCC+kIP23vvGRRbAasUfAnhJMyOllZpjGConv7De6TYo6/gTO
3j8ROHRjRA8lHe4NvIU27dKxZEuBBv/IjB2rXyCk2IdxACw7ImKp2VbHCQuWtSA5bUpDo3raPcJ/
B6KuJBaQKhpeFDIZ1JkzM32dIMfEiIPDT9NGVaYAim1tYC+Sc5O4NxXisqI96KSkfReMwxHuNIn3
3WyEYZn+pgGJXCANXyHIMQli0lt1bbr1ycCncl2q55S8ND8EnHNrKohwJeWgPuUqEIPQ9xCocfUS
z1nIpI6oexm9OWROfNjANwIz0V7y+AmT2ODAV+RjQ2wqj1SSA8J2SgGuzF8sYj53iWHGfU6SPn3c
K5NksKPUUYrXEd7LneRsEZ5LsxJqKlPW5Oy0VXM6IlxwAz6ygy00yHhAYkvXBUcLNUqy4TuMjkvF
InmByWy2tp8OPjoe1AzTA0jSFSfzjhl8OKfJ2xMnx4dT4RWgGaMggKyVfrqQ4xKNLQMBzSIr5V7a
YvVCuUU5YqX9BEMU6WCp1kB6hdm3Wh0wfcnIZfxQ9z0RKC1OT2ciOk786Y1vlKzjDS8zhCxNPOgA
+ysVtW8tqtkRQyCuRMoVSMlL5GS+K3/jB4eT93Oy0fzPCSSiHYeDbgjMnPQrt5XKdgoXtENNeWlr
Mj/5ZbL7FCbv3Usn2sNo6jNmgC6Xa6Bf5zMhLSwlu3XDWvj4vU2CENgMmWBZoK2jsTAKOWyU/lrF
ofGS8LrYhjDpnTvZTx/I8wLvHwrYMERVrl1/bcyUSYdczQ9kW3MqHSLuJVa5uVBrmP/Of8K2I4YN
ZEIg7+OQZWUtWOHpUSnAvARJ9eu+f5yP1T7o6pCJfljM9eDMMexLzyq/O5JNn6fW3YnbTdD9Q24R
DhDcW3bBkcRipR1113a2AepWe87+O2tvi3xxKTlbzNstfkb2D71fIFGEvU08b2mqZu7BUdZA8KTB
Vt7+ZBeYqP1+HABdAPrrP/aV/QTWiUaZ7Ot7KLZSAgPkonneaQb845+LhgWKCQ/g17wRakYbAXjV
HKqWSH+RHzFn0T0rHA1H6M3m8PChguSEjTY/If94Hs0tDm6y5nCZasHF8nUsaO4SqJzM4HtFzFcy
hVplpXFCUtnvpM43VCm7PmIvZP2Z2sGLuCJGCUKmtIjdAbmburl+qZdrI0F851NFAHQYe2jcnaRl
BVhIS+HhnCth1rbExaWEPAFsSEQC76Ev6HjEFTOqx/SKuTTrqfB4QE5HszuN08FP/iPRJVMC0b3Y
DdgybTsZFYV+UwaqD91/KTmyC6sRv2XKWQkUGgkGQ0oGPvD9wY6gMDSCQy+9/0Ujdqrad1SLqGZp
v92UidgWSHsafOoVHB6uDkCNSScWByCxRIRu2ZsFIm+2Z1nzQk3EBKvv9wBaWkYUTFSHicPRrCzr
UDUzTAjK71pjfkFQwWLNhW9sMA2vlyTO+JJXps2mQUAUrYCBrgp8gkTzfAYyG8YCCJIFChmCJ1pU
iNkNaQmRnd+O47rO3WuL+qsXD5TOPQ83oEtXdI6PoCIDEvhsHqjxSn+gaQ2wreKfMDYkYeAGFBPs
vt6uK8lbdMricQE/pT3kiO9mKIX7T5K+bJnc/JpC99eGBOcpBGGewEzh9otzfchGp8pC32SQyK3f
GVbE7jFMrnCPXtdWharXMMN5fgx60ASf9uwrXLAhK6dyh7jgoTa86oQOA82liqglpbWg32xyQ8TG
+FFIpcp6HC3Gkd1cLpiLLJh61HbL70UWKlNKhD2cRGNkdb0T0Jusw1KdzlFmhWwrjr3EDpP1Sr6R
1SRTGskHMhPYfFhQzultk9KoMnOFakzDiL2dfNkMZtQT0HFxMh5wEYorRy38zfewN2W4yzyZCZ+o
4CGxUZaeaTQ6iIDwl1Gu7lFFrQjmHkwANj61/H3AEE+viyB24joszyMdQLl0e/YBuakvk8EnuJmE
TLsHcaL45kKf4Gqw+clJuf1oY8uLGu0tm4rBg2z0JBpymZjuETR5P/P8oIjWQwhQXMYrDXnGkm8x
96CFQxS4DbUQzigIIdMyXGgUUQ3qDhyuF9XWllcwrYiO4yu20maWgpYqqcR5hoC73gKdsTDIFNxR
D1YYtCPBCc85QbClOj4S3AHIxl78sOZqpwwt2GZoC5D1hMs6kwgIFAWv4Gw6Iu3bdMLK1oTJMYNs
mCIxaIeRk/6+9IfTrFvhIb6XdBpHMqvXbG3ip4yXL1Xay+Hnufoe5SMZX/wCFGuS+LefrHypKOdL
1vQxOxCercDGyFxio0Dwf1hRc5XblSgnFOp5Adm7Jhy6TVkOfpej/Kn/nmDvm0kBEUH1z5d8fzfm
nh6ZMgLjTnxekUb/sIXNtZaLES7ercjELKi/M8cOjLGF4ZBqmJMqPdPSi1ZJ4qMyQOUb3f9KaSED
xl+G4+h9BJLwvWMtMJLJEicZ8UjgH1T1N3eIyboLDa32ZOy/hKgPPlq07GqbFmyItgn/iDKSPbY8
E5hlLm8v4s0+JGV4cfEgl5ICDHb8yi28SuQGBrhb2drdItveuXeGOTtk2kbKN2yGkxP3hlhB/Zg8
WSC+QHnbNynohzoNpWWHTGlk+kIA6AnLXfeul15rEIKlp3tV2109aZW02bp/5rjDNCGP1ECejiev
jtOHgOPOKzYvtR5LxKIZzVs86LPnJk7VNlMeCwx7C5GBIk6KnQlvrcHMRd6f0niOITN04z1qVzm9
vejmIX8TSqcv+vmxOuAs+godydB+fERlSxMo/oicKvgD4lzeeCUiU1NDPASYgmSjkACfd6xbGJXN
rvQf9lT4xeie+V0EITfdedX8fjT6ebBVqm7WvtxY/FO95R520nkp1mxTBv0D/8x4guayUYWYlgek
2f7x/RrpZBPpstsRW82g9vrcK9sMUCnTwqmx6+8cinB6KyrpY+6G7vdRTyxlqgkIsnK7PCPH9i5m
l36t5LtIY9nJ38CKINprN+qbBZQvHYE8XplPa1fMjSb/wxBRFjpncLCmdWd1Kxt3jNOfd2K1SAzE
Ui4vOWVzTQgZc6Z3dkTwuKeYzejZY5wGlP06lFS3IBOvDfv2Htv6IYgMHbkibUCqqdPYFFVTiaVV
k4ihVdHk4fGjie29Ihb/zK8SUDblmZRSgC77Cc/Tx1pJzkZsNHRSFqGyXB+hr9go29QfzvhIH0Bn
nzvHCyPtoTVrQ/dSe6ZJgf3PZQkHvqKBL8MidXHJYUQpe+OnHhvnbIav/TIPk1ppf6tGENtWkiQ/
gZY7oErshUx9BBLHLRTMGFLO3Fu85ktbyySHwnN0MOCq+oIe0rV2MKzWHOD+jk/5RnLPq19yf9ow
hFqeA8uKW5p/+d8BgOpw42RiWqrDVmNyJXH+OMdvvlk6XJl9qMqIxmUokyO03Ve7Tdgx1OD6BSLb
Q/Nfymy6PzbUyOlhHb91xB382jSz/gfS8JoJSm6bOGF8rZG2QRfCDHtCbNo27SesttxOupgWcAqd
4taOPhvNQ9QiIhhvVRcL+VFlAGelRQRrB/1v5LRvY/xVdeO32F7tPkem7jV3KR4wCseb+w3PqHr7
fLWIPLkIvE5119tYXD8zEHBPI+54RgSCNO8CH/1xmMRvoEDYY5s0180gHw8oqDpxa2vQF7AVVLn3
761tMvBxLAr2jxgldVp9TACm0zvZU0eiS8IQnnm/lZTQWVNCpFtJz9cVXbtuBUigNMYrPmdmegEB
zhicLUmeqbc+cvoNntOWS3eNiDYjIcLW/e9H1oZjg0uPeyyxWGJ65Kof+/fQOLx84XVLGWB91+24
+2n0UoKKtsK9cNthjkequ7oYzT4OA3t7txneUNhxgZBFJa/Qv0+fh33P6/JOkwSaKDQZepVPGeC3
BwcJGq+Bq7ULyUK3jVMcDDP3TFHJmS5+2WjR8CqcYOYc5DP/Q0AC2imig0Jz+NYYhLTi4nBOme1q
2a5kXoIk49jgeR6YqHeTW2y6qdPZuKZMk1vYRx8Xd0EA3US7CQ5ewL9l6M+CerJsM6eZE1XxujYw
hNqeDw/ww+Fz6A7tanh9CYx3C8GkkL7S0tW7Lx4g1NTP2iMGebHJqcO5WaHvR+wE2p+0D4VrGrGY
MjHADC+6brlEMEyI+Jd3RSruKDr2rw9FGB2MmGOOnHG8O/x57sd/1WDsLRSec04Ly84jt7OoFRl0
54gnejtimj0jh4QkvUerBBMBYDyTJIbivyqa7fttD+ayK0/K+JUlufi+BXrlLSap2jl2nrqvmm3D
Kvi7ftriDxMPJodwodLfrmW8eQ4anv3iTx9rWjIw4jIOJvdFX8mq4m4WmajAFE8u4oxQPaFe3aAI
UpoEXEYUoW06k/FmX/Bbn6Up9JKXGGTJJ0OiLuStvrNDd7L9J8gPYz/CTFK4h7PeKW+OfTx/RtCZ
2fpgRj43pVYK2YyTbIXut4Jvj2XzS2BUL/Wn6pHscsL8fzKMNkMU5elSIxemjD2tjwv9UmGmbzsF
8c/p9EM7oz0RwVIImtZk8E7b3slje6Zyd1mGIiqJt9cS+8MP+GPV0AB//rq5o2xaTvCwim4UTR+n
cHCQ0/eT+BDP7sF8tjqFccdACHqbG8H76ASqIS8hbrHx5VISgWsIz+QCNfs31EJEsMZCndMB7+PT
JzhAp3GITvGfx5cVlZw/m2qBLz9a1kKW539zT/TpFHHxlLOkxIf/kfH2fM1DjO4JmNoZ9+uuLNCo
2sAtWZL899xPSpxCxVbjPZPYolPrxEs8AM4VXlLU+z/uxcTxqyEqtxOOGz1aVe9bymTHDWwecBNx
008bsDNyG8jkQAOfFjeXSrP8M/3IMmkZGCFfhgahYdRd+Pj9JhmOLv+zPFYLsZqmSFHOTZYRSGa5
a6H9WwhksxNU3bVzSl4pBMX/JkXlblF0pK5X59Bkug/HydLW657/0LQt7U7uXbFysPCHEmhlaxYd
QqU/HxivUBZUfo7K++f8er/eMNLsn3I7hijrocv19rHXwYdi2HBBRihOxhnnnKu84tWqpL3cElDX
Hr4SW5pdcjMsjMGamGSXHsRPRMcq/R59I5xmn/nr+W5vbf2mKSWrzTr3evP9PvbqNZCEeHmUhriB
yGfFCz+oAse0d23BuxrpKY9peoFC6UsLIdT0oscB3Wq5O7Gn+lP4jS4t00R1zNYqw/hD3QhFO6GL
TIUD+msTn0ErRoBkd7j296WOQaFy+CXG2KDB+0kkcGMp64CmE/2dQ2giLu1pE8mXosVrYIAKTjWh
rtvyFZkJryBMlhIm99Gr/QdFwF7+GykvI9GHXFCQ8spF7jonP1Ugd7NoejwVG4sbpPZi/SmeAsZ+
TNeSpdpwsE8OCvI/jqxXtKh+UAyvGXkd3jCB1bUFkXjLBy0bXzWbwDmBucUrsB+FiPSRyscQTaGL
dCkIsaM6iIUMG/9+bCQzA/fjSpgDT/Yn1H2mZ++FRSYomDq11c8tr08qH30rGG1JFe9Gz0kc087K
ykycnhyIrYTv3CMpMvmFDQTrzC+2leKcbnIhwAH5VBctY9Zy1WDepFbETaEDYLwwOa77OS2Y9a0U
4GZvxKXAhzRXe0gtlVMZkb+R7CAeQ/i3Yiav2hCBCQzXnQS+e9rpBAFf4yN0Tq1CeQ+CmYgLxPjt
bM1KZi+QxnoRampb4SZwHrkJueTJ/UczLCcalKia9XAhQ9ocr4rYeDAyKiYj8LLKzqFrNxXaL7vC
hXf/Vu1ciQ5efgxJkaGIGdx2ZcGBo36lX3+Okg5MVJtwZjCx38YaEJbQJj5iwJthhTzECCs+2b9u
9wjaPM8ck4jaWelS20wmz3NKJrPdmJ/V81yRLJrfd2Hrv+xjVSKgk8eZ4Od+pSs8w+Hq1vtstxiR
6CKv9qzLgRAkvSvx7X7q08yvQfbGA2/Fgp3B5hiIgjCHm4jpcwfqXlPLqr4mCjAQEJIuylDtsil3
1N/A7WtsQ/7QA5Zf+B0yzCClELgcofQMItTsT9rWmiFH8haC3BmvxSoMU2UBd3ILJIPDFh5yBYe+
zC+Ou189orLzQnLK0rLTKaE4Tz1QYsWyAE11XtKpm3XVx6Kt/ii71kIge3HK+VWZk4g+bGeOa0/p
nJbZanOOZNYeiueCiHiXflKXD8Hv3MDpvFeDUHm3Pov8BDQ3rCCYKSfmS2nBjaY3gijnYf1yglqD
G1/q/OPNwkctGkmG2V3Ld4y20616CUlGX/sJzVpboD+LYnWvQY+8SSfvknRcq4Ax/psGw/k6c8IB
eVGuai2QGfAFpoRgjijijMDuph5Iv+FB6BW1BaXNzUv/6JdsE2H/4trRGBbtC13RYv6lBwuY5Lzt
oDEDxPyY7wXcejLWRBkR3gNAJAVcVG9DjKl+5rK75ZUoSicpHqPHE/KKgsNHxtUQ3BDNNUQLZ8sB
8Azr1Jc/RrELCHYnFu2blBJG18JhQd/tbzXI3j1xy6BJtT96TLaghWI5Nqj6KByp4kI5deMIZjk5
6QGpKBlDgfpflwHqOw/fQc9EpfsaTTK3Og6OE9+2BuE4hYrUnIVd1/JQctX+bhMBmGcBHMMBSsqm
tYe8K5z9Xv6cVaZ2J94j+KANoB+GYu7kpxELtLxSrmyMt4WqJhN764n7XS/ADZB1t7pMG5TPAfh8
3BtXs1X9fzTPHUvH9a83S4piXPmXKA9nsZv0aYNMnalXCeK8gcqdypgLhgT5mLQHJZR9YGI+zosF
S+9nHs+AS12IVKCo+ueuXufs0wmfKitVqZBcqIzKCHb8iAzQcCaGcpI+grrhGTbzJc1lh6/6PzJu
OowgJC1GEwMjUQ11PADzhKp2baQs+FNec0PuYXRkbME/+pg0nkZmCix4kcYe7zqpJnVsdi/D/TYq
FiP1cXvA009w9dqFguNCnU8V0L3LxPuipxT2rU7cR4Hre3vBPVXBqIAjfCLHaATF+fXAjhmBchkP
i5QETvHjxKq/kM7VQDJsd9LPDT11yk3UHX+sZp9NS7AxDYQmzvz3EnwfCyA0TMey7VcjNp2AiioI
WBQ0b5brlniEkqJ1Hu/rTNUoXa5vvHBbIuuKAOQPdDWdYsfOBoR9Akg3xBikNtN3X2Mfhama45A3
pjDYXsylldpCX5iVl5FvJhERh5k25Q2H2bDoKtL5+97ibe5+n3ix91as2UuTv4+npnc9cBlhCEh7
wPCT4Lj9He9E0gCpMWEHH1XBSSRaFPOhgv8TkcXF7isBwmraJO86wHOaOjFK2+K1atfSTs+su2wS
zEzfT1XwhmDO1GiBMtkknS7pb2R3MEdg1NbQDe5/7wLQ19jOvcy+IaSArkaJ2YU+fJ3BcOfH+odk
7rmOLirk8uqvpaXzJnq97ZO3hRhMtrzrrU0QZen1VzOUpQ5mbkwc2qsKx1Gy5mrBGLyXdMTIqe9V
wG5zygvLMK9/3+WslyCOaS7KD0XBz+LTEAvAzLkaZd+8ejh6XDL3mIU+qOlppwvWIRCRqm97QYhE
AfWNH7g5SYMLi8dquwSaDy5ETozRxshBKF3HxUJ5GF+hwLGPcg/H8nFLvYwsbH/x+DDp3TYNHmtN
OQVu0SSsEEwMZ93xTQc/aM4O8vYyhY7BE2u4jpMDWih2R2rIckm8CzquWZAFl/3HYPbYSfpvp35v
5AF6gcJSRyPqq76eiveOtGCs1zKJhFNs9JQkUozvO6IiVNWqu47aDIxIitr1tYhOxe+a7XeMKhvJ
gTNyg/bLiejeXzVUUFL5NtupZb+s6XAdd7CRs2edXfFiYDM9h9OdY0tioTaRuVc9mSQA2GkRxbTr
Ygz5uSJUY/Tde5ZvN0Eg07K+4SCRAcruhRiJGZdwOPavyPgksnrC9sPDKSMj67M8knQasmFe+RH7
WBW6Aq8uO1Tulw3jq5tiYLJ0UgVqxd98orPbf26bZjqAEZpGda4XArLpUs3Jn0a8bfBdtRe2tOkn
mGRHeV2aWYpZ6GO87dxdGkjxzOD0hLn7iENAakv4nAigqgN/kWMpOHB6exIm/2BbOgoiqL8WiEDT
KSH9jI60x8n8lsV1i4UEUJGGZyDkd9mt3bf7r9p8b6HKS971Wx2zwDN8b4f7Z9o7IYNUOCqzbby9
LfsecequSFMIf2KZpp0gjcGTIn1fgYL+50FsA/bMFgId+cppIZaAGlumDJZm5PF2mgkD8kK+rt4D
lUG/qSCQhnuByYgz93Y8e58GZ4vXO0AgxBp14rzhul3AFzKX0Bv8fWjl115Brq9Opxf/qdZZ0oOJ
nmfQuC1NKH/v02mTNaAI73/lSbevv4k8WYc6PGauMoHT9XlKHGojLen0MIZlLGjbsM1slZK0oJve
l+QU6hA8Yhkeqv9Vcisr850HSVrkIUQNBi1pR11qECxY74ziDw60v61GM/MBxKteR2d1qBDwXuJP
3fDUgZ/qPXR0NpvA9RU7dylZdW2ELB2hWlHjhh1nNfT41lP7RDBxmiBVfxKSiFC7LORUgdN1dGor
aD7tBhtnQCu5/1FBB4vyFnY97hyZEfDDTRr0111+gQ8e80ayOhxwc/5YU/w9vdMm8Zho0wiG5zVf
mYd+cs8E91a6WjZ0Je08i7ZuV7qyePhwMNPtHeOwWyOe6HxjnIffqZFVNA1T1OWPafk3YwCGZLkl
Iub3KWUZvllgEspgWxhkODjx2DvGTs2wNlcUHcjb2KEvE5dV2476xwFosylGIh9YzDnCzPDfd2YT
Cw2oMQLemVhsBfgLhzclamqEJMkfk5B9fMinfk+jV7AWmFi5ND0xJW6JGplziHqO4XgtgcR+h9y3
pInwnnQkEk1nSlVckU5L5iKVf8hLYw9os4EVxmSNZHNiKVSsaJ+Z2+2JR21L31bZbpwsLwRXCjSS
atrHzHSB2UpAPodfQz57J73JAazuMmE4hyEIpWbkQ047X0O3yfAOEGzlQOLLukJLYvpUg7LJzPwK
WqJmZ3wih1ZXH0baUQfZfdRZR8lpCsvvEW8hXMz75I1+TgsPPkbdoMeMTOBFU4+XhukligLtYHyr
9LjzajDSEcL52bW6GefLtKZjdyvLg6rC7dROzm3rYCAKqBG9Sj7QvuhfBfQTF6SJGwtDLmSHdZtr
kQ1Fgz14/s3AJk91IJZdRKRl59N5I+X/B7GA6y2/tn3+zEg/Pk2AsGGi3hx01eW2+eu5jJQqrzjF
VI5w6rrSXyCr7S6hcpxqQLjgZV0wvu/1gzKBiX6dhhDeonXGpWtLSz0r5knvsN0d4lVZOydKs9z4
6w+vvqbdrGxzEo0lbYRIAZP3IqD6AH+UR3TXVngGfC+MOMUkCxE6bQ3k49WBV0SX+m1i6KKUfgcd
6Mkzb47rDJ4TqNMmn0PZnabsdIThaO8xQMB27yRLxEmNVDxnQVobWAH6SQsxzDLcpECdr33U5IAt
rK9yZQedrAsRjYhklkeKJ+6h/Tbl59ssnZSJoHWiPv7eajobHmSYdeiBuinFgMprIg0A2Kent0Jb
w1EpOgpz5a/yTW2wJqEbfOoNxlBl6GWvj8Gjbmo5zx0Qnt0BjyVytMOAUPuVsMElCdNOl+GPfCK4
zMAwnwcRUZpfV3Rv9AOU8IgGX2uND7BoXzBqz3ep6hagTNvdxkVhvXq+rTMIf+Fn8l8sei5zQHZp
YeVqGb6gDq8dZwrbxG4VCqj6EPnN+2v9YM1oam5eVwRsNhc+/+2LnCpRJ7S/RIIEEkxLdhZv722l
kLhu+PHbyK8c+uNrwhPVUpjdHo94W42tYv+rcmy33wpU+cnBkafyxyKC1mxnMhvbp+Hw/Pi0Nsaj
tLoKVpoj2OE2YN43ZSwOYUQxhnaraRN3SxnrwTDA3F1ATBJylkUMGBuli6Tcn+ZK3WK5eSDmsqZc
b/oc71TOIO3eogRKDM47p97TU02FYP6zFLMKIJkj4z57Ym5qRCQIl2ztNhC5vDy7VApP8rthKkye
EZ24L7HV1I0LHWwT/uxdgH0NITWyglx/xcjNXIzCFSDc8oO3zrRchzzVLvaE96wsw7udQMb5wUU0
aCRL0+x/+YSTvchzL+rV1Bq7VS+L3MhqivJ3NJpvbBt5w2OIWVl8jJmCQLsTpHvPdZmnphuaRsHl
MuYYdsj71D89cNguvrWqA2bDD5q+tzKIor/4FqqU4Zum+4N1Tgn1MECmKD4Rj4kAeRMpO8pLnfVS
57iN1hQvBQlhSWtVlwSmvkm+ngOmHTHnmaYuzrojBivkWDJ0vwckfXPmfivvphv3BWv2k5wFm93g
yiOSEYICZNHZ3vWFMwq6n2YhYZ2Mu4XIygKOdiklzEidGH4oLtjQw5pcpbGQCzTohtO8fXF9AUP5
HMUF+9PjHMO7rihykoEAUAZp6hpTHAfQaHnmvCzUatOc0obT3P6d/lHzcunjMfkBOL5MKhqTXIqV
WJDfY/b3hv/JP9eewaGLbY/bSEfTdPsU32t8K3ly9sdwdfj9GYxgH/NWiGw3/VREDawboAIdUZMo
CVbVx1bVH4CaqT20y5wm1zfNTpeX+2jzPI4LsnD93IJqgcm0Km+WwL8M4GHayx0FDA174Tg/x8C7
CQtq406PSLxwqHaQofjtl542hrQkEEL5wCl7fSK7kX0LfMF37u+1AHC+AHO7w0mt5zZBbu/z5DXf
3QCay5Jp+7m6zNYGHNTcWErEH7TUJr9bsM56weYFixssMPRZsfKcFmGNt1LTxbtopxWFdshyrJ1t
LnKPCa21TjvB9bFEJFOKbn8Qb4c3vuoM6mdUFyE0lRKNYvOst37KhmrMTt2OFv0qjdMI/gRQ2zsK
MxVMGnZooEajNdgBx/9K76VwKxhMOalGEy8i8+6ETRVF1jtqG3Lqs7g5oiUmzD32ghzi+xP08/Uq
hLIzeu4YJ+4zyIDvdsoFDT7DGqBDcpUPeQ26Sji5PXFuRbEE8vjzMs/MjWGxCjKuR7d0CWAeSWDU
FvzgmXvmfq+/zcmIa/qxlXBYVwzn4LVmSp7gafTAh5EODUCQf2Y1Q4z24lYKchBtKSOZGTReYX6F
xOOROhzLUvevZammdGq77BZFtwFgyGphmcKQMxYmLGRMQmNd1igNhvUsbY22y5xj60wYeCe/GKKC
cVxok9eDDkYQ3c6nG1AkihobV1LzKROuhL1EUPbuasTgA5lV70H45QybpDCCsWSS1KsiUgSCbpS9
WgLLH0YxykxEikjo8w3zl7gJxUCUxyp/7CKyFyj7wFBCeuGTINp2hlgdrZj4lybrhUCU/lsyD8n9
9fqCk9trL+cG3DW9YfCadyX9aJ0VhDb7J3JhDu2PZJr3/tzd9wPa/fOSFsGsAk2n0OJAjCQQ9K+r
k9UsMvMdBQnYvUFEKYfUt64UIMdC60+ipwp96aByN4TRpCuGSz6j5SPJ0UxLWQSbURlHID9SW2hT
pdkvzed0hOx+D+7WOiPXGS2Z/gHYVqoC78P1K8LoqX35gBQCCSdX3AbY6Q1PJEJcn67mVY/gzSAg
IOJN4V1KPzwpNayNPI7rhMu0wuZNVA9Qo9EpyuRoA4Y6QefqNItnCvrHKpNiKA6R5Hb9T3CKZxyT
HR8koJPn7v3hDqloI+HHnu0W1/d91FnBdPBNIW2JCbVjFhi8DUCIlhzU1DBMEo1ftSfDxDcHWRyF
zzJYNdRh7qNpmAvkGgQpI6es4OdK2HT+xGI1qykcQAkA48oIg2iNO7frQSz5g60bXV/VhsVMSyd3
SXSPJdZnDlF+JAyWxZSaxFEoz5Xf1aDKVHGpVJZ5sdaf7DHd0243kUgWWdjH5lbB12VnhkqLXUuC
Lv4xc0+O0BBQTX7gHNyDPbcr5rcWXgMxAunC+DBsvpr3LUJ+iO/nhjONwLE7TLyuQIfNiIlbj1HU
WhVz/NqlQhKeBeGOwt9hUm9Zi0q2HaWMy6UbzUJNswzt5reXI/N2crMWvHuub4trfA9A1mGvzy+b
sKJVI1bG2ywRdMkXQf9xioc54iSPl1aZQ2fafSfBqW8B71EzHF9F/HYBGrYZXWj6SxEeBaHbySFt
gPg64J/pD4qWax0Vph0uYadH0Ep+P+uBZLRy1MoiufUFSETS7JOdqJ/BxUpLKAMB85Q1ft/+EAcO
2NlYQM5UvWn3gh4uUuvGLEoB/SrOOa1WoGdBpSVG+g+NpO3Ld29LBeQ5QHW3g3CY5tdjQ9KwTzwC
OzfpJBM5Uriqg6FRnBAWlY4zR8bMyqU2QEbjODZaP220d7gnaCLLls2zdvLNePGXhMSyaVCsQ4f4
ATxGEz34OqrqU7sf682N6KEYReOMoHqJbvFaYU5N8390TmZ6fbg6scPBZUVFBtQ2qNOTsMD4C8yT
Ewvx/3ISXzYrMYsYbF0L6ekvEpnhC6N6mDe2hryVJa8/Lg6BKch9fXL+txuHl+nbW+PTS4CiulNj
bCt8bLYBw0bJjPvEGFh8oUompVp8uPmm6zstNHXzbS6Loj5iUeHVakxBSn4onBAGomjTa4ZIBz1B
wU6AxrH0nBNEyBSBVRowdM6y3V7zYDGeFXBtfnGf9olQC9BdoTWUcTiTnoZ70cmlU2Jdp7aNxv1n
Jg0d9tO9+2KSfa4E9rrOHww2TJr1LzAPX494akeoQ0G6zDvXaUtXfIZb6Rb0WWU5NEIdpGD0UbdC
MHAx8WUw1RWPcKWH2LtpVwzeOGK+W5Zcxr2fIKucYHj5OMXt+cve5Ug3CW3HbifnviIoKqxEZD1/
t/swKmo/x5w5QNfJLUdmVRvVIBhf8g6G7aBS1oz28zHQaLkUVwU7uaHM/XOAsUlTII7Qr0Evo4ba
xVha8JVQ9wGoqIY9HImwT0YwDXdAjvZpkkGEYihWTs0vSCnt8BKsuBYf8Q487WKCB6LsZvpv+J/s
D0fz3AK7LKEa1UoYVBHGxKKTp3bRR49f1k/qKUeAlxcTKOio8jru/9YVVe0DSSZ/0+KgXOYP6j9T
JylOTJHcHyPOfxU0i/DR4lZLJSxgovjLItJXdjCxtyl/oBYrskNzIoA0pZlMIrXGjcAQS90clGV1
gO3LEN9kYUvPvrNV8PYGPjYeuN+zYg1McX3Ev8EnpvK1odQjApOVamq6TFoC6lofBKt5GCuaU0sO
E6nDr9SRNrVTD3Df7kFLo4+tPyFI/2oLGGcEymVAW85kQa9WfZZ+KIvuhBXRCVcJZjO5AMHWMK0s
KlG7wDbP0kLsWKUSttqjiLnRIc60AIbRzK1vyYXObAsQY0Ja+5NWgfnoWhzf/RjXPiYbJWG6rlTi
H4zySE19P7rZ5Cq1zK6f39CkkNbmUtWw/qWsSSg5RBNmKXe8o5wC96P3vnsLL/by/5hxcLI1Grnp
67OfLPXJwa/Rq8jN5o0ZYZ6JRFPlktm/sBJ6Ar8uOYRYLPfe6MCTWTCjuyC1Bfwhjt1ucQAkQxzX
ocQcJiRtqkwZF4zPrhh0GLTG44WNKYJ9/Btw7Z902esRrMvRkXuE8JPLSihJOdEB3TSFV71SHJFK
8oDg63kVJwsD0stDC4nAt7U0T6V0N4ZPjTcU1k3NWd22bZ8S0ZC6xhIntQBnh29+plQf++SEcKuf
TFbtEpHc/hV4VKPumwJ/ecopIjN5736AWoZveMocX1WS3J/eM2Vo6kYFag366+dkRKeRuf6ogU39
buQBrJwZ3fDcuwlCXOTb2G5jK/26FD5qYgAc7Y93kqBiXSXYlsfwk33MZCUCwKP51SszD8aWGm3v
lBsxvJLxel0EgEo11S1lmj1IEkRejA80pIEyiNUlC8wBGYmzx7OdzboF4xAVLSY2LZslndlP523H
1vW/WOhCRN2MYwjbmWI+s4YghKlXvSF/vIpNyWrwsLXl8IFbX5LGBmI7QdmUuZC1i5RXk12le2Kg
VIkcboU9/h3CX/Vx75qNpgsjxQyZK6I8pukXXiSHmiOSu6YL/hI5FR0kRwgIvt0+yDvBo3vGrzr5
ewA+WSG9G/1yyx4QIPDQy49wi2GVKifv4Z7IpueMw837Mn2JLGz+unUNC6Y5yFeDVTYfFZkVZkh4
EnFeBsPf3q8XTkOh6CUI2ZojbNbTmEcTlY5A7iZzafnbJRQ0JYDu+Z1Vdmnmk1f3JR1mRJgBoqxi
KSS9l1TGxEDE5GEsesRQYJtmG2zF0qiK9jD3piAgVUbc9XLQ9x1ltUF0u51J4qYTgzM89NyWGj5M
pzkm984KkomhMSvS0wL6CjMJo49M+1QcQqRFlhcD6ZPs6fsLuMRH+3asoTGR42pZZ9+tAt9ZL75N
iJXlq766rh5qELIQ9srF+q3gWzXast9DoA74/417iDkRBm6NMe9u5NT0DMhWG0n2EQUNGZFf2snN
SFsR/M0P5JlamloT3w6g2n7DBhbo4AsfDjmTB8NmEuOihWgJEW7bTbtJU9L/LVZ4NcaUxYPYqKpP
REfaPzJJsFH6XS+KiggSYWJ5Y3kwDXHMWvtb/Az6uIBK/8BBiS+hTl+CrsBXLVs/rI3cNpB2LDq0
WaocEQxIjd/rZcelRasC9TLGnXlOv9h8fgIJbCGWLijbo/KP6J3lUuAcF+tKigr/XXOP72IrfFfJ
qlt5IVdOd/tih37ud0YGodn2rHd6hO5U72ICLam7v2wO09COvYm0d9+5u5GTOJFnVqhilvMiAaXc
W2iri862iZsLtq/bmk6r7PQ6o8Zz/8DSR1Uu6FyyPJd9nw88ZJkMhs6f3w8zvI5zlw//Qmqr4+nq
HzeZ3kjVufgBsAZ/8CqcXZsExSey5OVS5mgqxD0AIQak62vcsNYub/t5fYt1Zo62+U5I4ibtHVEN
SzcaLjuNtWg+Ni6V8/A0b9VzYgZ2G4u51j7ju7qyE7yEWuT+a33LYgBf7NB/hKCmrt3unIO/2vhn
ieuYxTOn4/EeAw7KJZ3+a8Ofv0UBGTP2LjCF8SQgg62tp1BMzCCT522dcjiS6zwWbbr6gtepF6T8
iiTVfIZ85NZq4REI8ZPFQ6DdMQDTWwpJqvuRfdI61cRmlgGSfwIL8ac0MkwW+jCCErpukoMnileG
4FNxm1LJEMhi/6kIvXOCuQ1tbxgPMLcpyupWPTBkZUw0jEY1NQ6DaEjkVTuaPNTzx+jciZR+MJ3H
zoDIgPSZ1gtpKW7Nph4laZam/favXxWcs8k+LvC3rtDlJPwu8u01cl3DP9P3peBpmG/6OTxguUHc
dB01s1wAVGWiyIcZUJIzC03t4C83ClomfDU2j2hiAJih/Caos/F28z96/ccN9KXGuvMDky4cFjAZ
NqrMDTDnHW/S5jkizaBYusb2CNUUSgGgVS3Ilr3R2jquj91D1p37WFZMYfk5jfDmFQbBlFERKLMH
VQjW91aOrmEQjXcjctPHvt9Z/MaNk5rK5fXq4eFyHUgBdPFrPeZfm05hsS3YnTCCLHHzhG+UqV7k
oMG0yzYfDwguwBguM89xi3xoio2gHYDyPzhnXf15VBLmbqJ+fQupd/cIVKJ1TE6kB4i/G1iK30H3
1BUjNuEgnMQNATEKsCNHD5RDRT/zuMIXz2xdhe0vTa3eaHyTQbA19HdBXIXRcS0fY+Zzrf2hfr3I
dYgA8PLGbs2ynONJApAMfxM3KDlqjgRkPMgn7Zd4DY/aYcHelfgkRYQV60T6gkVXbZJHAyq0Jf6X
V8uSVMh33uq+5xF5EEbHXUlxg79S7qsi3ZVU0qwW8ubje+NFwNAYsBRyFe67jy0ZBj0O9CA4hZpc
ECXaxv2AxzPrRXw9CCFdmAKKjsOCe8lqxVLAotrmVMpT3hfWCNL0KNuddbLs66kSblJ8sdl4O7DQ
+q8u6ZzhDMRFwVd5sv/htzRofZ7rQh5t1g4Rv2MnXl/N4+vpAS7ip+avN4OiJQX4zv9iDBXMQdBe
qk8Ip4Aike+HMeGs3MJBnwfl0ncmNWZEL/IFYlWfsLLa1ml0Qskc7kHVgUNnrXgd3gD9v4TXAKdL
7xEGafDlJTXxEmH+hhg77tMRq7/gqk+fiFFy1w+7KkODWVJ4uowWANneChgEOiycG9RCJdE4+hEn
Jtv5PYDo3i2/jSUJkzDRTzaZWdUtM6jvz6d97ecvLVggz3bSjzed7LWZj5NMa/az9EHUSstFQhjV
0xhCqv7ezfvt14l7s/f+EUIOyEP/Cv1zjAlzn5oIsWrk/PBViOKQjgbmHxlUYQjRB0/doEW1T5Jw
f9mvF1J6EQD8+briZlm9NSlcTw7oDLu2r9ZRbnnnem6jCoUFmdM8I5BwcYcFB0BNIm+TQCKyQNlR
Qgai1TJppONhjgIq1MAICeSO44YdpLJZ6SoRSxq/paF4/Cpuyz6fLCOUWT+wnP8otXyhtpevRN7i
ha5S+Iuxa18/6tq8nrC8qtbSTHPaj4EwwiVs43I+QXFu7ZA7BNxNFKsVISeTR/Dc56dZAbBlhTgm
S6p+l1ISt5lmjXauxykeex4/oCwa0oYG0o5IucYi3GS7sFPAivn4D36F4ZPcq52TmZpJJ89tYWyc
xSa5kX/xkZvLWXp6ypPtQ9B+TU9stNZVvm7ZmEshoubgpgkTrp8hJcin6lg4Ltw2srVnWhlGsed+
CVgpxzCr3bQvMHpA5+bblxp6bw6Fl/pZhkDma9aX8/WOaBMX4YnuceSwP24b0OANMGqJjEW4Z/QQ
mbdAkE30VNIeRFZhLb00NATeFPOlPQTefb4qlIrQPhqq7qpqwjBCuVIFZ4o6F7GG+VjZJFAIr35m
bu+MVsRxvY1twLMaWXA4HAYYnLHP1H3iZSIZbTmvTnRrulygHKyidXSBkfGQ8M+ctpGbzEABi73Q
cvoC6fE1SITQLdEZ9HwtmD0jAcdoJM80X/zuimhQIKxAglSH8rc6bqYPeMbYj/VsgxIZdAjBd//h
bnG2A3tXdk0xPZs0oWm8FdV6+evlZzmGRr1xU5yClcmFMBbDDLRrKoU7ovN8dQhJ2XnVIqiNTFpC
fS5Lgnrz60xqgqiHpgZ7yFX0X6nvCkEFbr5P2eKiZ5AWMvsIuYezPU+PmXo64UQm0Ifk/XAYH67K
LoHNNPdxG/0YLssQUQZh1ZHf/g80yMZVrDqLSA/ynyVqmv2R3RrC8AHO4QPDam5mr+WhP7BSR9Qn
ExZBEQ4xIiPtDjLGrW5d0++nCUwJP4lLlTVvZ50xzhVJPqVC5/cr5E+KW/eLJnQ8zLtzLZi/Ogys
tHmtxVrXcxpOjWyaK/+0iOhk+cE/eoPKF76sEyUPUQtIIimrcMcehVZ8z2e13P78DiqSolYBGosr
ScZ+ky+cqvX5E9popdC1b1zzBmsU35DeaJk9SPx1+Aeka2n+1VOVwkCl7OF8fyBLq+p5oAYu9ypr
0IXPJ9Iwv2GRughQwGyHGNdyYPOR4AjRt+tlhrW6RuBAgaf+okoHxjDrJCkE1JpibxRJCzXoJEn+
/W0Dg/hvjYNYUhUbdgH1aaUxHSrfWS6lbSftEM7VMVDA2jzhMExOKJTD1REajt1VSOQW95OqdVsk
jdpddQP5xiC/jR/WhYFb+gu5FwZ+fWSGaMpDFcZA8iRpBQEG9Xk4JQDwHJZtPkOnmsEQ7cvY7cSF
cwmy8SwQp/uiEkd5blXq9W0mrlx97MD1aFGx/nTNeLufCOJ0rtVGmvt8Cp6P9crxjOT1NUjHCzYJ
RtDW4pkh9KXMxzvEU7otWCcKgmd9Aj5h4JM1QH0rw8XT9VS/5bGWKcJWOMjcH5qhCB4iMWx0WVvQ
UCklIXBnGUyook48FzQv3oXzPbvKETq1RXT7tlqFUFQc0u8TrWY5wh5jaYl+mJwsrGVw+xrFevm7
vq5s9HdvIgrgBZd5q+bs/BXPPvC6QMm4GKVmAcZAGumQXB/+LY5h41jYkDooigErLgtDrBDVuzg9
Nx6av4b8vdiQODpFRsXCDsDXKqocxzOHvr33CM5y0LecjZ49qpjeYZQi/OrppeI4sMXrWMV3DMak
+6zUQ1RCWQEHCSAsjHsKBlQITDuUMuoEEqGu3Dl5cFJTJ+Q+iIfwGSGZRP7wkRv5yGW+pydnienF
2UTkzgQ7zyGONgoP3lsCOlGYmeDliZdM3x6/GnBlTArly+BIUrFca/yTvOyBS/5K7jBscEVUOf6L
22JQY7xpG/I/kntw57ufd7jhbN4yon5iGbYCvpUfNxHaqW6aegUsp/j9RH/NTRIADi5lwcsxvD3l
IrwnP3HXjEIKi2yDIvZsK/+awfprGW05j2wd30XfsRp+5yIVYBYDIygM2McC9n21mk6sqlHnmWzT
WYVSlb8jL8ycMGe0gk/etINP9wnSQ9kgLHXBb3hmjxLoPou9lfNEVomtu7zAqjdFynz39stZJu29
QvrzN1fExCETdL9W023rTfb8icpPiaCcwL8cLChQ6Pt5+OfpTIvgbwyeFJFbR1xTbHaEp2BFjyMl
0BZN6wduMG38N9lXfzszCyoqwSMTR6l4CQ3mVrcGMx7CEBhAKbs3kfCCTjv8BO1qjyAQnj5D+BI6
NZpqLHKLJNX9A1eo2DAZdOiq4M6wBX+i8w6xb9FyRMUwveZy43McMHJCHzjZBZII3UjnUEYZnwAx
/eog1ZI8vTzhaC8YJayMJh50RoKZzoO2920ylWCbWzU769qMDRL8GwbTT145oMHV4fDYv8hlhVv8
Cz2M+T8rqL/RxEp3UmtXOXfsdAk1bMdEzMq3Y8sCGWsqez3bZZDVv7Ti5vsK7B5wi0CH/YRktD/c
GMH0mfJQkO2joVC+8lnGT/jT5jJuKTImfa7FrZHJSnvmLfuymdo+c8B6hBdOyLJKtPs+6tVUafKq
bYxUyY6b5I0+eZjjXgMXRTTsIG4C7JpRJggPrqyIFuDeh7ul7bzc1bAG3J/b5z55zSwl0d+Tngkn
9DscFfTrGyouiOmWy8+5IwfBkQ59Z5G7Cv85Ne5X5HWte6Mez5g0AobbVbuJKi/071zCzMnBBNHp
2LIuWlcornaSaS/bVMYH/NtR97Zbvfknc6982CQwknJpC9LrLXO10sqPtt4nsmrVjyB+m09OwGLE
swP2cSvoPca7eCQCW5In2XxGixzTP859KiMAx+6+aC9a3GHCMyIu6fd1Di4P0rqkIcmevPIKNaVu
DhbFyj1HDcD6AtZwXsPCA3rccUaW7evOfhTL6wYZa1nrP0H1prViB6Nqoc61WR9SzfY/GowQlbAd
5ZQ489E5ojSUETsaHstCE+bWq8QvUCIxoccCGtgq0b1W3Qhu/Fl++tyCYEQQ4UzzqkrT7CIE7ggM
sPU1fdx6h/LvD8WVDHzGapuLhB7EF5BSNhPDTsEEPRY8cNjHASMQpEXI4vdbzxnIgQw53qH1H/zw
HqhE8U7XvTkJmQvBrGehrNatOvr//kdMUbJnWUEd0zii3F7YLKniSdd9PihGgHTaOYvYdPIuGUDA
tyDuWerwtVJloHje0FXS0Neuoo5Qq0glI4UQW6qwDenYKv6vB3DwdErUQztd6C/BHq2yR9hT/+6t
fUFgFCc75tN2u8XnjM2InYkXxLCbbAEfl8V2YGsFzVeJhqk0E3SLjR65+X17sGUJj3ZFV5jxgBnF
PUh+YNaBMSPaG5ifRgfJUdkcPWKYNKGBQnWh9ZwodkOE6cn2RgwWncsU0hL5JoQsxg36GnR+m+Q8
1qBxpfYgIlvPITX+bwPMR9QLHlQAiGq+eeQVjbRAQSQetylV2llWtcdmEpLJ3xLubm+Hu5NvXS9b
6pnvWmq1O6kirKMyn/J+NkS/S3ziVgfvWkb8SyAvP639TWbCInV/Zg3tgEGuYcDdtN/3fGCsHldt
kG6pGSlVLuGD5KJPeOPYlPJy3UEieDwqihgNqhyaAor5R1xi7R0ZGYEYxrOtgMrt/GfqCE+ghw2X
zQ8YARNbd4SfU4bipv8rDqjz3sk4BFT5SHDvlulZFCld7ArRksAfIUTa56Dh7KqKx0k5zz5GQUN6
iaDXbK18e4LHO+APK8zXh/T/bfk1BG2a7fDmRVbs9WJTiHfq1dIv8xOVte9EZgo6EAWGlFcWLxuI
0lBYB0boUQHnKsKIPInKCfbVhG6e0R4OJEC/5fCQ9rMURx8vv/PNvhuxvBD+CJeTvuCIzAs6/wN4
IzJq6DX/75ZUmtpmiAjuoLxWw6KHy/UXOkNGtYCyC34Yw/o8h11wmaMMbFeNHQWy4B6XH4mpeWq5
40wHp+chAT1xYp0Z+47+HCBahBVwCIjTsz7wkQzvR0gfBMPCtfCEpxQLc2YW1ZaQLib2xOvgcOtu
wk+7LGXmTY2ml1gVenDoffJTgas9t1aOvv520YkLfatuRbZ06Aj/HqqDXczY2tBBV6BpjSzZBtx5
a9NH8vgr4rC37KRLmHURCU+t9a1ggY9VLjQ82LKXcJzLc5Oo5H3b+H7mvX2xQsr+a0PBXfUyEb98
GT+8k8VzRykYC3W00kOenWOrP8URiwhXhNzEhCgOC3gdG+ljFBjT6LIAFiop+chRJIGQBxraJBiE
ELES+QZFDX/zL9jsyK92rR+lx9ZnvAOBncWxtv9XXz8Zscth5IifqGQAejdKY8TFxeUs9FRpLx2e
GzcYp5BT9GSsvnamkLoursqV5fvK14rOqglBonF/8r8qthpc83e3MKCIl/7/WTQHG/kWX0bz3EXE
vGSiwkH2R5MEk5Pd4HL4yyu3bUuF8zgkFisz6JW8tzKtIX0sqACzprBijmgmgcq9BKU1ItQD0oev
f38RTZEFMGDE1xiVMZwEDetmEiVpBI6scAl//9GBgX94WdBBfBVJHcnrdeSh2ibNPV5otM2tWgdH
CQB03Edon26JhW78HhES+BUmk/Ff78kUU0zMsbkziIa47idHLFj0DyiTARwYZaTkzZ1Q+iiYNhDp
EWo7PukWz5rG3GZ6Wwp1xc/3NnSkg1CLLvEI4Ctp4a91QOxqv0jvMQb8VodBaFqLs9/5NuGTkF7x
WPxC132gnmvYoxgyd9i5i4jSyOPhXJaggfhPfBIqVb6xfB78S6rH/XyICDeg1TSpatQ2EvtVoqDO
MdEqU8DONV9La/yn3TSfx/QDkWxN/Tuzw2R5KCxbrpavUF3MruT01ct7DxjH9yey+DzSUlm1kVSn
OZVRJ4ftbZHtxPDhU62dtxBsDRjUUw8uBKjhrG82XK9tr3Kc8nTz6Tp03mlq0QNNjQ/jFeAnWIkE
EviF/ky+PcewaR02wQ+XCfHzVcYEP8VibZUybVcCNviL5PZ5NyFvfNjlyrMGJ/VMW1EXe8A4dVOz
9dA2qcyku3vulF9xEk36pXKLV9P32e7vu82BSsR+F3p6vc/EmB304AtU+9ak6QTOSjahBksEj8eJ
Bip1Muo0SXwgr6Qph+mgA4OtbI2Wsh7G1/KbsOk8WEeJS7k1pXwc89A/1PdgbjfqaTM/UFC61/cm
cRC+AL0EgIz/+h04KFQJ4TZHddzO0tzSUWdOqhIohid4bRj3rtpFM1Pf3scg1JK0PaH2J0UJ3qiX
oz7JqO47omVb1zZU36kCaD4HRXZ/H9P01PES8PaCpFkRuhDL94QwlQYeYevSuvJSpdULn8brCfbh
frLPCiANFF0DlE7igvOYlQHHoGVJnZG2sXDFr8olUJNjcO0zgJfw8L//8Tcf5JCiM1UPFprjSmVL
SUizRX16JhWLyVoJSo1HfpLdERD+X/0o9qUXsSqLuC4/TDU7Tx5wj5ANfieAW2DvS9r6zKYfu/XR
iQiBBQmuycLI1gAfbn0X/oFaSldStmAcaAtaziAzKmJEc6Cvp7l5RSTLkeXgtxIlbwuMPkeqB9ZR
Ab/rXJcYrbqGN+b4TbrrkGOsh1t7K/o9LbeJHNzSzNnh2t2hXeGoRTG0LqmxoseEMVv82RiaSjyk
O/Vj+xnGpdrwt1koml6RUpT6ZJP5JlnE/u54S6aHFUu1uXSsSKpx0B5n4LyuK8abPStb38Oatoxj
7JVmBRnJRyFMHq5TnSpLCy/CgWH/1E+oKTXuYX+fMvABMcPEu5VNMTl3WEMS9BDoMU2Xfc3bQqKZ
5SgSAotI2Wm1Nuol3gx2aWndvCtbWz0Moeva/BPWAnTTNzGxTcnUHJAa+2czUbyLJEdBN1aguZCo
i9NdSwU1hL0nDIoC2ABQkQQViBCmYecSD7tIIRpQui+HHhOKyIKbC1g5rF5RvmX1aQ01cCHtV6jM
7XvrgBQ8nddf87ax9y1eXAjaOpymSN9bZtwXDIYFjfEwGotftISjRngcbG1ZieOkKhQ0ZVqDrcOM
rewN6RXYs0JC7OiAwQO7x893bM9MyVCrqaoM95hs684xqID42f7S+Vd8aJciAeQxJ1ZAzSmraRcI
u0l09RMCf8sJtxgB/VyKXlNce5+aSomNQtQLnJ/LWajNc5DjDSCgSmSn4xT18Gl/jDfNsEENtHEV
+GDQdDcVhB0QvutrgEld+uIGu8xK44lYUID+ZGbsRQ2lZTrlp+NRSjZLbd8WRagR8RbyCq5//hv+
IPZmr2RPanT4q5PzsT+gTBfQUO+NW3hcPz19wG+2/q823y3llHcEhPS0B5fCS6TtaaV+YNmliN+K
CfjrSy9ly0ynNaPAA1Pt/zMUeCpbF7x3yLmdHgkrXJZL56q2BlP0q6SChFZKLW+9IQRv0QcDgjBy
jBJf6u3syHOwzjfZIUvSk8XGc4+oMO0yR065+Ak3S2KV8REOVinggY0WOM/TuAC1hRFHkzVC1LnO
1+yZ8me6bBQk3/OvKjx0EVOF4KK42a10gIPcjeGwMEKsmAgTiZnDSwwwnYDbFIkRzBua3IHosojl
qCLrAETbg9kfpZd2GR677IMnUNkecUm0Hhe/EMo/eS253BRRucMkQbFOwmeI5D5rgrGqf/wPP3rK
q/mc8j3pVc08HKQKtqdBacfbtzA/eLdIwmCFj5DwgvdbH/y24boMRymVF34ap6RAbULLMdFmRc2h
QgdDDAgFFDJhehNwzg+bxcDYYyYX33U4TTXlW2eWMoKw2h0X19jJdpxJEJfaPBPM6hz3Yz4Z7/Ui
s6QSIOBlUsKdwnNVPERW9MFkc2jpWGHkfZyNIGY+iTU6gj8E9768FNScg3jcLoWrODqM8au87Vd/
p3mVoTgrqEY9cy4YPtVX9QDtLtkaGQzEql/97/hZ7auKyFTzeHnqx/y+3B+3NRkiQ/uNjEZDRG3d
kRS674vWyCwKHYmiJgNAeuvAc1FDt+uxfznrj+Jr5QcKfUEZh9vFdDIJuF04kflOEIHoGbqZlnin
851wQNx7CaUE+MJkvTUCuGvy2p84MUl/9lSmMMC9PIqxM4TvB2HkKj+P8SFf9b3PKaXh2QekhQTQ
FqZ4MxzbZVKYC4o3ZLmj2q4xWEY1dcbPlQykRHasQfHBV3anICmjFdMy9sTZauMbtd901E76Ntg6
YTNKlXngTCKKq8dlZpFA8DAVX/848LIjAzE/+Nin/i5lqpbnQ4SEv18FqL1siYHOwjb2qT3mB9VC
UEspv8MEnNMkuxXkKXC6ezFJnvaET9sJ3kFgdySCfQnuY1IMGMVZs2LYd6AKoGeE2x0sI8z5KgSt
4pwvuV1hS4k+dCElYxw3dU95f169tfez1Wf0y0uCQMjeYnRYNP61Z2zvDSqSeaiD8bmi2R7HQDM2
MPAgZ2QXF9868wUqBtKqoS5lwmqKcC/lPo04U2f4ShDii3OLAs4gJm1+Fn1zMnQnfiobtOhnP69s
FRVNGcS3Rixm0vi8rlKyCyomt5LiPHLjnWe2bt6ID+RU7lgdKP+4falkYSarrqy2sDuv3V46vmXT
98BsjVRosIeaJHzmOflkN/igG/vLT/XhB0ht/aatfXGYL3ulJZdjdbvEw/1HW1dOMP86DwyPHmxM
1d0GH7Sn3m1Bufe0OP89gTPGnypP6ce+G1ONALycZHAD78NqoQN8ai36s2Ivv2utKucoFaGXUwqV
oWKD3gArZeQu0d4Vxp5gKlIahc2zKZlSznUtsOdH6LfKpsyW1xt4lPsncYGmpeRRaB2UzAW6oKVw
g8v3P6VaXT2bq5VgoQHUSFC8rxJX1XrnaxDbf0k0DZrsbYfwW5Htbrtfi5WZCuNiMTOAJuaLadx2
yEh3RyjVB81IN27NyKMD/TZMjjzkton0STgShC7zV1hKdThX2YT1Pm/rE+sPLLYO3a/r8mch6l7R
ZR2W7CDl5rHsgGW8u19B365qZ4soGDjr/ReevI5y2Z2sXTY/ig/jHV7CrdBVZ0BGdg+804Ec1mYp
h6uTh20TlDY1iJDpGohB5+xh51hCUF9SiwfvZZ31i/+1Cf+W0ri3ofyGaoCaWly3WBljaG68/wW8
6ITBiHCtdCRoshsXZ43TWSDBT2TFVCLNoPe1zc8X70c0hiL6LUMkNAHELcN08ySUw5Bn88SCbbBH
dAixxZ01EEDg0OBb+6XmJvaASA+UktSaT3QdqXZVVDbJ7+aUotGbY48SAYL1QtwT7w56APJVPWBq
9kP0tf3DdTnS/rJ0yAqHL5tPIGCX+lsCdI5GEvOc+UjO3j16m89eQKe6ek/BYdofSJ0Z3xnrXuHe
mS94DnSTTImoNlk8GLssYiGjvsR1c3VSpqN+0YBuZTa2GOV2mLLwjwYL2qSP8bKO3FsU4PFiVV6p
YWdyDXcTuSnlSkf7SiAdm0Di5+Sx6WJiRXgbvtyo2OvDvFA5C+u5u8jm9pjq/bj5p4yof4FFxK7l
kt9slkhyK+V1aW7/W2c/lhpCz0ZMeLZRt7KOdhdKqgKrOsDqZiMho8sflH+7lnpKvBA8NGdeHT2J
pdDFfscethiciWjo1PRjhabPpHtv5GI/h31qFT3X8ZUOQpJC2ESIF9fXxIf2APcZixmPsk2YZL6Y
6e6bPkm2aePa1Al55GTrTEZXlbwNWoSkzFcIn9b12mAh5UDsRsaPqyV3n1mGeJiey8XBGb0Huiy8
F1OpggcD8SQbj5Z+4KYc0ElmvVvNCX5F96SazVagVAO1bF7iDm6/kZctCGHMEO2KiFuYl2jg4LV5
STNytIYew2xVg3D6tYcRkBic9V49EGFWTpnNcL0muT9jYi/yZTHu5X0l73YXffS2aU3QEscGalPn
+SB0sr6Bhal6lsho8iLznte2xO1SCFcV0omQzF76wcKRsMcstxddIbexVOfEBJxuwsusbPR+3CGm
OzeWF98xdgtupWVmQgFW+O5zAB35+uEsEsYlpYNTImA8BQZKDp66Fe13HTEIRrLQ8KNqBvOd07r1
MrGPbFHDxyhLBU5ZWB8AF05yeZklaaI/kIi2ndBJhnFZK0cnIyIKqu76939yPnLYlOg4FQmqnj55
ZBvcWCZCWPGFl03p+bY+WS4/ehpg4WKo84dR89FVpEiTE6fA8bUqw61UlYhzxxUZiwbrRwqWe3GR
pWZxGq2tQTAQceTpLbXYM3hLFbxdDiBaU50evaugwSrQydQyrim1JJTzOz2DiKCFRHo1y3m/tlbD
HCuZPThxnaB0IoFs5wyGeFYsN2pnB7tYtw38YJ63TUm5JKJ6q5rgiqgb/PWu2Z1nzSxpMck7UPzX
A9z06tXTSuJM/ns2/R1mt7TyJ1g/eYXqVB+n9IdXAXN7VHO5xOy/HVB15Eeke0XN9wexPNBxy9Cj
yDoxN90XOeWUD7yKpNueSXiSPoKZ1LVlaeVmzQMHmT13K1FovXGcPRVJn0Kt6jc+fjCcdGxUfauc
7YoIeL7CKKYyLM5ppo8PWwfkREhT22+JpSVPN54vZiI+/P6z8UddA8+dAMXmuN+wC+5KAnTbCjVP
yEeSe7EKGFq6s2HpgQPemurjqDHUNpqN0J43tFRNKZfCpK6IlY/42QTPC76OxLmz+Lb0SPpq32b+
Bxh8dt8JlhKGvs8++eP2345B3Iy1PFb3IEVAgdExUX0+syTr99nprhI+khtm0O+CciebyXzN8SLl
kaIt5mHLSz6K8zWI7T2tqwpk7aPAWOlWIbPKcZr9e4lSxF1oRnVA/AyG7Yv+YGGG51dmCrrlVhU9
BA2KA6ob8lEMBMVZwjNsoX/qUQVE0vRdDAqPlqSGuSFqB8N50d61W1u/jEZz/h/do9rouEWLgrf/
TmaSwPKoKzpoqQqGfrt1RCWhgrkBRQJiP26isG4K6DV2gzSfHFWteA29FzFdYYGvBDBPOhpfMjS8
m8aKI8qIQiVEKvxf5M0IkpjZNUF/flO8VrtU2alZOohDdMC8+tx+voiSWEh50rYxGAbJwmXsdLcL
c4SF+nfQb74k4xrmrcc077wW9KKCb/6k+mXiwbMyEnTgwbN2ayVjKDNoQIYG/eeqHGGOYXr97M7l
MQ2/bJGuJTpqj5w/9lnwhfff404aKpLc5Ofeo2opV9bJ0WdlmK5srb4YUqcH8IFSuChI8hhIhVWq
IaaW0cN4e9Bn5u9gvNQanJNTrdJSlM4oiKbvXW8wVMll8ZHdd9FwuYAERy9B90WBUWilCvJhpuof
YiOz87jnFSBKQOfAzeXba1YfBoRvuNTC0dpjR2uflmCzlqGM5mb2zr9Ip39QUgenm2l/gEWGH/86
m0RMo2sTKhQCeuunPui2f+YYz9FarV9FPQPAfmVQvJ6uYrKwToM28TFRWmB/cJgJx8w3Z7zJL3WM
hauziNMoL1Vts8iK3FtV0ojzDTr+BEK3MP73OSH+Rj/OA000MkE8NL2oUIF+eOv+7FnphCAJx6Lo
UC4WGAHrtm03DjpHA6iOYdoV3pgYIiyHiTTssnx2hEPMhsBblj+fRhmUyQKaq3bin79WslDYcK8T
yXzdaGrVh1qEDrncDh7yf+3s+HVlEciTEzNSqD/I42ofhjUQc72drq77BcWwTfLczbpdCttiYBQC
aSAwsLMstHzsDC1oB0e0S7BcJQL/x5CLN0/Mkst1bVDLIkzKQmVQDtGDsfhUe02dLn533RU9g304
WZ+E07OHwTntdJDO62uovqMknFA6AJRB7USQXOBvXmGQPlTIIPn22LHMQWFAGDJhIhCchkxP0ZYs
9AgCNJHD8StqPb5TFcowPrH5h1QZ0GVCM0m2tJlr0E3p2pnbW4qYUH5eMd41MlzBOQ8hoUyZNthJ
WkO9kiGXyxYUl3owC4F7TspHXknuOyQKnp/iQeO9IF74QCDlqNbmwHvS2U3j7Xx96FB37dn6UY8y
JrQ4OCKJlX1Fx355J3K+7Ar/0Hn+Fvg01Dlhhecl+LS8GKgiDqj4D7SXEoyL3IhNhhbPdAjkiHBn
gZS0JEmi0WuroHxO+lEOGnq181YS1t97EX0jvQXkT+Q9vrD4xAu1uLLY68DflX+iNuwsEbwA6WCz
H4yYKw0+0Q1gb50H8LHhaGY8xSzEhMLiVzJ7BPpQX+vNHrfKplkg/+DGU0Vop9yRsl5bMqbYI2X7
SHZhbagLEAxi0lgkeC4N2AjSeaIcfAHBbYj+B0byqDzDvDMVlDxwwDWwSou/BGU8iVXWlY0ywhFM
96sgyxK4+zmL9Dh/9M12YA5wqd1EHNQwGztq7GMol6ad/AupCyNqfgx0eGg7pUHXQUQA2fXDZiwg
JWsMpHHLknlOtPASz/mR9Pr1LjszwrBWahXF+EgsKYoFiiuILcmJXASbyBehpsnj9XgwOsGhIxb7
gOy1o39trPqidEkx6wDW9PHKNpPTJNyt5q2X7atnShaMoHGs48BlcwVIALsnzYhTNfchpSMPGYrf
mXXtnpDKnGDUwEgZooHmsVAOgeVVZ/rk9vB+HWk8qFIOtfFJzKNP3Fd/zAVWJW/ClvI39+HGGw9p
9WHia8r9e+N19TNEYtHRM981Drr5ZUvpuCM+WCMn0X81CHRqJpVF3HAKZPwF+ieoS15KVzED80UA
rZvjjcx2fe+6Nokbk00zwtBh+1Z03h0Zi9zQFBFrdi1R+D3NNswp8GsPXnkDWO2mIvR/JM2K2xUg
DxB38ghmB3rkWnmyp/1jzF03lCOtylvn7AWu6dvTYvSON03D4L6W1cBbFuv+/0hskPLcJwWqndvn
x1eDAM1gtLyoEf8bM0bR5X1EgVyK2OLOemzIMv6tHi1h0jV8Gtyw8CylnOQBtGhTShj1d6pniHa/
6YGHlUMGYll1pLwF4cWJDm1qx4lo37yu3b+cyAilQKL9MmehO4a47bKxTWpz/CvDB2O5OR5Asnb3
9Btl8PMkdNcSxe9ppNWnWP8LiPVYir8hWHXeIl5XnG1zWfpTx7R7K2APcEtQ/ZKwPJYZSM81vcNG
lO8yGW+zN9cy62hTYvdzjRhuE3dvY6GNDR3JmjCpmvSbLsbpAi8V2uXkkSkukl4EHkp417MsS+bI
1EGlIiiWvh6a43vJWLQNnSkyYSIfOArBH8ZGi0XHoICbSXi2aXJ8Rx5j35wWiNUDfQEqdozlyPRF
Bu7LBtLmgKTWPHFl3hQT7GoHdfD140IP5xuh5pZb6klT/S5BbzU5kkkxp8sNbNwjpA3EOovBO1bY
LVRf+QO/7MCU8RGLvX/8oVrJ0TXGhQIxghkUEImVVPT/u7OwKY9wVExzDxBOY/m4r5+qPIVgBXh0
9gQZ1IN51OKf2kSr6siTvnKoGGrMHpJxR9QN0QAH4itS7IHPJ4mWpiNktAH2HBpQ3CXrwvSzs0+0
imWYW4CEl049FwPhjR23CPnmTlOwC9jIccK6/BNXP4HLws4n77BgsCIae3/UDsAnvB4YpA9ue9v1
NGf/BjRgCHC2bin5aVNSJ0V2U+TdcxiogjjBikYlRn+SbIaBKi4rCrBpKXMekLtQvuAwMVjUkzXs
qC+yanePYLUhKA95rUm3l1CqFL/RuYYkUYvOiGZJogHenYMlt5RTTfiEECHpIdrvt9GX+FO+KgXe
zGja7jOWEdLaO3szrnEi0Yc/wTvoKeav/rI6ra1buF6b/2Wh1QFl2qi6L/55F0P6CcS1iQTfv0nO
CkgL/hdjvsv/1eocjYDNTUzhF1KUilhOguWLxmLuH0g1Wl+vCEv6DpECeaIjrKvVa1Cg2jxr+Xat
+k3eT628Vql0m/5DandEhvgwpzsyupQufsD4w7EQ5i7YyaN7IBEVDbhD+ztudvEzklgOp0Uh1keg
9LJTFuOcvlKUgYAWzuqP2HcOl/4gzr9l5VzdOVK0SSX7NYT5vvbVvPzxHwSq28UtZUZU5Kqq17Tx
VETc2EAAjAUKoUfAtWf7N6bis95wGmc1WmufOKQAQsbgESMhS3ciXNq3/D9YjvqG5hzWHthFgccl
brBmlw3VLFO1D/8/xq88T/YxH0PPPp8r0lEAfqIqzQ+LtJenZht4O+F112Kv5tySax8awsJOw+qf
K01Tx6Vwnn9UBJVZQkdyjLn4qqg29UlfdqPga5PPK3ryhaw+0Ei6Lu8OL8NMmodyeHw1PFBnU9mP
31BRCMizvgM98OhUrWtA8lTwFNGpNeRJn5a0Ns+YebTm9nh0byu5r8vT3IqgdQ/Ay5/s6DjdywR5
f5qujp0VxG+UXDCzo0MYfRxahBwD7CZxSPLfXpjOjvIJLdMdGTloJYC5/MOghHtWYE54dTFrplP3
LvI29NR9AyJf7DkTwnBw3eKVDKTmEWKz7NRQ4RG7St9hnQpCT4MAS9q/WMFVp46rW0oLy03Q5FQa
oOIFRMKQdG+vBJ5LTcR0/N7YKWw71QIuJtGZUpso43vGTIxcpRbuqA/vZHqt0y+HPZpJNrvET8HG
kw5NIYyJLUi3ewub5mZSSiadK4jX49obb47KzO4KGQloyoEVHd+hCEMj4rqQVs4rjVUa2ePvHwLb
USfpweRP69tfEc0rpZ0fuoCXkZ5kUB9VAJfh5dRNoyAvPTmX+wnU5/aKgVLx0spUZJzYDEbKh4WA
YYMbJ7l94Eghx7KVqWzjvdt/bud5fyavHXTqvnePrBuwZMJ71ebfCnRgBvYSf9vINA18nC43eTjZ
+p/8B5hx9f6UdVvkrbE2oC2hQn8Hn56TRuuARTzCtNzNbK/rydYz1oXvUnl0BTgWcMl4Y6gbdbMC
CYE8KEyLGuZghgXtKedLldoAXVtkQ/M3jF8+9pN2I8Gf5OYd9B2XbStUVhKaza5sVQqO3ASlBzzZ
XaHhHjmjO/Hm8RULBOgtgy83TzBcMkxCshd9NdePJ/bxEmOORRZvkCI/9l/lKW6TdsqKd6S9lxf2
8xoZGu+C9tNEsuAqH4Z4EMR3MzHpfOEyxTeBEvyLDXeFTyuGQ0F//HUhyIoLRPgX5Yli942G5Onw
CqOot52a/FEajeMy8vEyoTxjVtyD1xWrwno2xckkNMPlwIDSbZQR/wbl+1IjWkZdrKHJI4J+uAXP
Gn5UMjHJgmSETseWY/LxZSr3+6IeZo82uyT1dYahu/NGrvrJ/StcC69IMPQz6EHaniP7b/EM8hnK
z7F+g1wXV7yVOxxB1r0M82roTCngaptsV4KLgzTJj75Snv+I4sLmDYXjdWxyy6HcSW3NVm8k6JYb
QcBuTh60jvlOBIhbG0yrDIzj8lWlXTt0hCID82tY2tGFFOeAvM6inJjmuHLE9xT8I3uh+5kQ01SP
ZZGG7RMZ7GHBtURCBAgT+VXK7QkDGQJhwu5KkUGW9xywmqibt3Lzw6XwLZC7lelSSfHF0Wt5rJXj
ToVPeK9YHwFWb6kCL+SegfdjHyzWu04zVeATnEfSZDyizVVdpOuHi20M8gsTmAgAA5+UEmEkj/AU
IlGZMY8Fwg8NywsesfP94hBzhnesuEq3QDEV7GVGhlMFYleyR9CXoC0NtVVYDUXyX6zRfqbfEQ0L
F0uxFnyAn7rpYlOa7Qr1+jQikMAqvTavWMh16l2RTstrX1uhSMdSOv9m1w8SeQxvKt8jUBGA8luu
ZvFCVwG0ZYddRFoNeI9ikqYXJxHuhHNsAv0NiZvKl2QJsI5V2DXuvOqr+PTX0s0h3KgfPSWLinL4
y9zu5Mm3rKC47nmm0OFAt2rcpLJfCz+391dij4xXzArLrMTSqhBan/b2oj3AgZ5OKJBGM5dbRKBu
weN1CYJsXKiATSCVXdgav9lH3Yj0WkcPUnYSlp9AF3+BMcNicL9EiB5d/4Goi5NqVmB/gUzZRG5x
IN2Q+wAsjBhqK2D+i5JviNJzeUHb/EhyRJ0ZZYjRRf3/lnEoSDELROmi3umz/03UlSImNpggrOqj
tlr1RaM7ZlWurJEmgCyRmqviX0/AnzFudNrb3p+Qzv2s+1Tg0xrS4/A9nawI4tUjsTad1djKTaOG
tw1I46sT02EpBDJNaATpa3iaP0PiQLs+/3sL9dnFs0odVA8+6Au7x1ooQYP4vc08iGsbW8lvNE81
QQ09YogMNp/Gq8MprRLAxCpTpyiMg2wutiviP3obzrRN7pPm8orul8flcheLd8HJ/kqp+rAdqiBC
RC8Ye4TMMFQxjNn3QhgPgaZ8QOqSJBkvTqv8aAx4elaodwMoZGX1QKiz7S3LCecgT6SRdiGCrkrE
M40zL/2ghjLC0LIJbH/u06Z/Y8EM9Eb6ny64soAPniNp8X5YPbbltq95oHS1hIYjnzyiLOQouNrr
TjKgwsmU4Z2UgdLYcvc0rHAg/jYKAIpA8em6L91qxDhHhvQEE4eapEs3FUpLYLMUHw9dsgRsvPSW
TLRAInaWtjhMka70P4BvApGGmdrDU985o+ZhFq1vIOIuJ1JsaMUW5lqW7auXtLzVGYaX8iq+Ld68
9MomKt6hcVaw3kBLK4yD8MEV6eQOwNE2Gjd4iGf8EHgwR4rEFVqUqBXCGt8ulgc+0qavObtLjU/T
Ysj/Ky/8F2x3Qg9+kMpvNntoDsqRzD7f4WZsvxiSOS/YvhrAQ2YrZ1fS2XW7k8z+syOaHdgtlcUq
S5QMNNKVBux9nkCg2goDaUOxE4s3ct3CpSvyPbz0+inyUgeyhyGW2MSWP0pbsOMgXUuXGhMuqWl6
+0lSvVKVmPa0vcS1sW8vzoO5ziOz9gxU9cEAw+m+8Kqd9efSrMuCP4dUm2/Ek1zSNNeFex3wsPfX
5dq2pX3g7nzXV0sCDmIzxxCgLbJ17ih8DrwPEefcBpv5DzWYutePjR+YGyzluamXFCzGSLWUh8jf
cOyujFccN5OCQckri3gg64nzjXzcl5fmhhZFdz3D/M419/OkatuqUTfcNe7qoTzDGukgoslmAhb5
X1Ygrg0UG1NFHWqrDxCc+hIlMGuqfGnzuox3C+LJ+vXA8x3JZZUdzvA41knpT+STHXgUCjdcerKP
G0FTPaaxuST1ETCmXC3MAyErKdr8Rx93Bp+xp69wJjyqS8TVZtQMhQM2AApc0hbfUvGS2Ia3Cy0S
MthKoGMP6+D1WpnUlf3tQ1TRGnE1FSL/OA2M3zfChBof7eYVnZGE0BIeVrK3RpH4X6CySlsdP1OJ
IwxFz/NopQrixbiRwvb05Tm3pYbS2DzfoYSqxZGkpNV2Z/EyRSTdq1uouLKewv7rL+MvhebfC7Fs
oYwOIokq15b3FVwkPbLJUEok0dweYnI0ACRqxyH6uf+W1VkscIzbj3YJhpis3ag0gcd3a4hzpqjp
cpsO7NxmwqUVIRPZpQTBwDtWzW8m+dl4kgoTchF2hKnQ4qeB86ek/DuK1mE27HZRV1OiLdc27fPT
ez6vWlxxij2bpJHshcFVmXUMlBsQvyplFramVqfahyJdcpeJ6zSYuaZVVHkRUSop350z2vfL+9Tr
QnrT8JQj2gQU8vacK5KxVCgi4ruFXauyXfNIC0AqACv0NRDVc6dwWvhMLiteqOXK0AnXS3I1aRyt
991/UFp/K3zBon5AV2xNzNemrSDdeA2pXC7/s7oQnCJfYMxZO07cd2W51qgdTjqgChmlgEJbJVuR
eYavN/jHEH8cXh+WBEqDtmDAxRhdJmf4esmGtENMQrf2YRFIMlDUmieD8LbGnil0RiMqYj02w2f1
HUp4HZczPtS0BAcYhqYcKGg4XvRzfEgBrZs9i8h55zB8YGbLaBCn8CSxpR8KXZp4865geI5Nk2Cg
GwIKomxjusMY6c2Vr2U8RdxkNkb57w7c8Qk7rPlgX1nerZpQBBJd4Q6ct+B9szgRTiHyfQ4/HQTr
11Dme5d7bU7abKet9K9oX6pruHTzDBV80oNdJd8IEC3GqzaLzprkPAtFBLXUjYjk/5ZE/tdEXacq
QfrIixmafbnn7Tjg9O763nXldterCEXA2ZR5Yc3XWU+vDSKJmb1LzQLoHGbznEoKYokgWH8tBmhM
9aIDoZjS1D2Q3Dk4AfSn37t8qL6OQHIrLEr4hnfxYzhZr6qQAVCJ0fA6dkf+2VlALUZrH48feMIu
F0hS1zmJth78jaLDN91Hl/WUQBs0tbJud3CiCNVCKG3ycb1IuJ+e09AsDDPY5PSnRHlHGDHpEuJu
N3h/bOdSh7S3sF7eRWdrqMJFFgierpQOZ7074JcDiON4taPAaIr6Fv+QrPMKlLRaYFQzHm9389gu
Bx03kAUKldjc3BX9m6eL6B2qi94s5VolwsZ4pWvYTSMku2+1+jN8Q+RjjPdxVz5mnECkGIkXcQND
DflKxXX+gtZhpS+Ffg7ZmlKcjpYCzJP0GnFGxNUsAAPr+M31UGiKFnjD1kNDk99VXq9IjReQF0yK
3QooSKblOK0iRQaMZsNh7xfOJbldFMrdGBIKfJpaDM4f0XPc4b0PEvR7JtD1Wkicr7wfb4RnCQkp
DVkPGIsNqtHeHqj4pTZ4u7zZHkJ5HKQ70dkUJUijRCNlg6BJwg5vjEPkkzD5QtsZbcYS9jYqG7uw
9B27gteqVkteIoF6z7ERSaKBqBtLoy4kPMtw9e1BEp470d9dpE3fNT1cjRpstOqflVISulP2A6qZ
U6jfLhiNcdf+I8ButIQpNV1z86WDJGZ/BIZ0Mjn6rGePpIKCYhqPyxWVWoTbu0A07c/45MQKy62S
K6tVZ3e/RhlKmk5caQkyzddXHGUvFtejv4rn7uGPSK63vIClzmMbHdMpSoH/Bni49S3hE6Km4ksv
eFdMWngGTNxx+9PsT71x/ssfV4oDy6gME6qU4qONMZywidCJhes3GSHXQt7lOPi2vrQXveiTnfnJ
Ukr/XFjiBolGn322+cTO14Efss95Fkj4Nl4ngVcf6an5LFYKxy68bL8P1SAfg5NFpE4RvpHttXCt
c1itUyzyZoBfdFJXKGglLJqjsKqcszLLFseZvc6/IA5KRULODpKCY6NEAkMDRbmPY9wny48cw+ZN
mqtXdZlOkAdzPPaSkKrDwj2YaSoVTFL68IFIK4s0D1ibTuQHFxydSM7FTqV1fAuzqL/Wb03ZTEE9
XzFYBd3NTeX1KoFitQgsTLfNE+Yq6vLRSB/BvkkqQ9WGqNg4uv53zrsGpnqUrYJPckre9BQ9X9gL
CZoNZQ1J2p1NXeT05JymXkA1Etj1BH3pwQwoYT40Zk5AVD57H+MLa0mBb3ICl02xJjH6AHxVuk9t
N9C+AEBLGeY8MVaSDyEbsqa2biVq6OIvi6A82IXX2TVYnDciwevA5uZSETlQt8bflAK6YxAJpuCa
/eY3r8JQ9lfGOwnGnKjc+idskY2GIz5PtBWc1W14ZoNlOa3+8ZPLan2xUMojGyTkCrIx8PgMkqms
Q1pfx+OsX7pqyVlE1X1mRq17qtFbGRMO61/opSmj/qmmM0DvrkLiE5onYR5cQuSFs0g7DTpuGBsI
fAj3a+BWt+8CiuL+pIowTAHkakPwhg+BkXIlC8VK2S1V9GMkyY60gVQJW+0PABvA58vBxV/YpUZR
69MOcrqwUrtnizD8yeOQ45+Xp22P7oAxkHAmU0L2d8ip3Z99DO+t5lEt3kdqsyyVOM5mOvvDDjqL
/GIZYT7Z5jIJlxQ0ZRBYL+9CIgQsFE26fibx0fg3FmP3hN/batzQkQOqMQakz5QEiK+yBqxAY41h
AUsbcf6T+m+FG27z273keoMgFh4vHGYxCVxTmr/6oGkhsr7UYdWUXaqSHLA2ztq4CmASeKuNV1C1
LsM3k9ZHFBe1yoiSYcduBizaqR6p39hCJdyT6ZcaFFpFJmKx7OynLI7J/GjL8svnPXNIAUb+NZkT
b2ieGUoEjoVuh9umWWxFinujYD4rOMxCmhHcnEbRJMEMQgP5DIViJaIPsKol2bY4gj8SUUZ1yYX7
49M3qXLnz9I2RzGhLTd8RZxNP1X1L+s74feA3duGoWLcqXKtiCFdw3cb2BIIz2WQM4RUw0lMDG6J
N8OahqUxrWVRTZXQsGmgjMVidWFj622G9jYaM8X3W8s7XAwpqGZQQWSS7wGQSKIgmOsbH9MPFvty
fpyXrATf4QCb9nLgOH55Z1hYeAYO1kRQTKgk0FVl4OeF+NFkDU13SvASaSb5+5ggMNTKT/wl8S9v
BNc7023ZJHfDXy4ZQK+IPlVECPjZ8k65XNa5iYf81SKla8W6NbKkv4H7kFRyxrnyEK8PZ3RPEW4N
wC8NCrCljvmQVRCNnG95GFh+ncsjcMnrAdYrHUtHNBuEkWWp1IcJVN7VCdbbLN0Kl9EJQEchLL64
CLM5EY7VIed6w6JfmJXOe4q2bYrRsf52GcxlQHDplWVjF8EtRVsc5t2quTVnJLbiRPEJUFtR1Mrf
f0lEP63Yeoeq04orZ03m/IcjhXwhRJkNded1a38AujiU/VaQ0gUFmbOpQ8GUX/oZ35sny2fvDUK5
N1Ksh/ElKCQ2onAhZ9k/RX8vWwBgddCF4Uubr2oXHahg84xRcrVZV777gLvVbL7JT1OqMDe9U6iB
WiwLS/tozFjFC0oQwxqunpB+2jmqvSW8qZBjA15aoPROXeJccOE895DM4G9fjUp/Ewf6udruI9Nd
Ii95TBragG0x1nr4ShYnei0gwCEphTxfoZjB9NbyKVEGYouhxmamNXce5tf2vR9lF+mW8yZY36ll
1G4uJOxY94UnwvVSQXe2J2jfGGIx9+V9gItqORtcJQstY8QdWZH/Sm81VLUUIt1uqcHNHTjTfGyK
p/MYVlN91bHm/Ccxth3uXKGMuTGkz91TZZBWjhyVYgM8p8MY0YpnrzBM5XXpYYl6ompk1io9IwvE
hWmvS2q3upoKrzui9TQAsgvclKW2aRA/uzO3RBsdLFYRSNszNlI/Axk/8+rMUislJEq/gzRmv3m2
bbbpPVtGFF0zcDOY54YwWbWrDG9eMjYEp8zNhPm8oQ5UHeO50DxfsnGmJ4PpcEVgevd4/0OyL0zn
r6rDE5LGUM1Bw0a6FrIawlqdiMn8RUdxfE6FbWgxx6JkSaLAuulbWhfBmRTX6UVAbrMivz/R14ZH
2B4TDt+gVyPqtZRMdL2ZkBqzzLf+lkeOj1BXFa8QvI0QDeDHZaicIzzy9YaHlvXXi6LhHDJ43Cg+
V+O+6gSwx1LLO7Da4WtF68TGnis/PsaGykf8Jza9B7iOZ0XKlGcqPj9pQJadxO/rDjHqB9VnE9K3
vuRT9C8bg/l2PE9OvgjQDEKnAdgemliNcMUtQD/J7oA/FhJZDlD140M6b/so2lSEbuXPJNT9LpEt
FhW/94eBCI+HNWFaDuGhbPVvU5AiooStk+FLef2HtDDxCopmLCQ6Gotm6awVxiXZjq5Ys2+chjML
KjD6S1wjp4GURg6iwRgqVoeWYzJ6d4dMGct0f46fkgFEuXwMfQBTEE23lgG3f9pS7XVXeLpYDgIG
llAAKeNcDxQs0uRxw9umXl6Vpmo+09iGI9+HZfL3ef4wx0nafKMU6Yf48+B88+Bqk5fghZT3oxM7
t69CRacdVk8my7FihkHulOiB3a/SsCQ4BSvtOEQa+vdbEZUxz78u/CF/RCEGgOymlk9cu8WWK+5C
B3XX9IXp5aedzEmjwSYWtHiPp+8rReCUXL+XDDCsw/t42qnmU2Tf3nS9m9K3Deq1rcFtm4jSLCKe
dQ03Icu6L6RtvsNrRA+qYPtENfzNwYEYNNmvzU86X+H0w0tHvJ+QZ5XBEqfhJ/f8E4PdUF/wTmk9
AP5OSn510aT9IlHznFRwSNwFsX2AhETaGJj7DcOboQY0oandzUBj5WDaVuM55n+jaN17stB2/erW
05Z2nQJcljD/fmoyc+PkW6cAxDdaIgTDv9T7TUTsWQvCg5AMpwBOcB7L27Wb2AK2VY8txg20XxDe
mfuSUgIe89UrYSko2/OPnmiPyQQjE09NKshphxHrpvyfipH7k272X24mrBiwyEmNpL63+YfEi0f6
67K0TCkpQttBGwWTm2XNHFpbj6G+pwGT4memif6w9sAuS6Q9d6ddpMDSPhMYTrZohykw1LLceHU+
fqjPOX1E+EX3/oQc38cKydqwM2LEernUyf7BM6qnCyK1VKnHaxXimWhhZBpHRYUI692AsNROdNCu
G9t0rRf2hwuxYv1bCFoOU7qWZGfKyOdpl82xV8hjwJt3SnktCiPJ7bq7sxxTpk/dke8O+tvHAMkV
dug9J481u76oK7bsVzik6LHgF3xOMCngTC9ailyD/uPzoSytRxIP/mKmJD8qGddB9oj0fNp9ppMX
3PG4zpTnEmVeKnyF+owUpKVHckO8kfDeJcnBK+DSawEEnAbxWR0uTJYexXyu8zHloorZcPaqaSMR
Dgmw+a+QWuhV0SNCA7oEqDn60Vyjfvdh9Qhm0ptI6gJ8MNCdxyZUf0sDYAEY0sV+BamhK9a7Jw6n
N03vAAG8Fd2dMx5k1r/CYzviHshmcuGrnrCb1zZ1Bq7Dhi7c7WckKFOPGtf8GZhGZtbDCCCnYFUC
WXAct2jUAHGPKdoV5QZUBrCgp3Nun0AIjXGQvURLv15V9LIUF71RIRoFKtb6EUGq9zxwt8bT93Mz
aKOTPyBH0jHpw/dm9ppZk3HzbZybZtrOR5kpv1AtUMVy7MmREUMGWahVeC0Csk2b2AARm8sHebaP
FyG3ql2M53u2TxihKFVOjiipV3ydSJcUJTMLLi4u1OpJmW5dmLDWn7MEaJbAcCdvqiKrLz5S1dVc
dK4NTBDI695V8b3bSa2eZXHI3NGKUMeqYb7joFcF0+zOa3d+WlI+f2RthPJxXiMVUznzrF8JbnP5
/Aq6hHw0mwL8tpR8lMDTalwOAf3UJvWkYkhTKOAFtHdKFvrn//l+WC9Ujb36ET3OwwLUQ4UvR8XW
p+/nOvmwH4fj/qpu7Ut46WnsJCkCCuSlZSkzLJCtqDiZFCCh5JsSm7eyWUY2IFEiA1Stwh4euAaP
FQypeHw6w4+6FNsiX+6xYIWamzRdNNN8nl7X+mx/Jt6H8AHrmcm5xSVMA23kOIOnldgkhJJBYYzA
dNsTgIXKSheDYesDWwb0VaWva4ZK7xHoqBiml2JwWSRq1UvzMalsqF1DVop/FvQ/m8JEEoIHOFsf
LQQIWuucD0LeNIaHsbr5ytpUNt6j67/+B4NX/cXkRMdRF3H1nXq2CAHOvCIFIujiDu1DJEne43kv
qQpk6s2OdJvjvmOUaDzT5JHQfu4UUOvw8gHTp4REZU3BPpSmKCOWc6ONsPYT4YIVBEAttqNwA1Y3
T+AcB/+kYbCZLsW0MfKP3Fwz+0xD1XmfvyXEyPUFofab/5Gyr3r2LEVzUBNBdjGtYTZeeD9vuPXk
hT2jOxsI6QQwvX5SMN/IUSprMf1wnJxLDTKu+6/OwQvl1eGNHygSPhRe27TQkT3P1/UnVQSNeKVi
iQLOiq4ujpTF6hJFEhk+1yrsdMhNjCN4YlhiLikIqxXl1QqX+cmreVHR1AfzBZYtlkyTkZk1lkmk
zLz+brDrOzHJA939QVZhlZI3QC0fcrSI589xYI1ywGKaadeCvim2j4Ld0Aw4GwFVfpakMlEStuGo
AbU6XbzKyx4mDB8OgfMIcG6TdvXZ0Oj7hniQUmT7l+2PEhxQW5ilLqM8hL0f0qCOAFiu2WLyj7Ip
Oolyt4dNu5UvknnLaCMvx9ozjII0MjjyFJF6+oOPEZUEDtMn17Ob0dql/VxsMQ/9RZsPE1pE6KJi
WGCBA9KKqtzEQ8s5wfjqnzBCM6h/rkTU6qbt1z3+cIZUecBE9LGlYghSUMiq7RC+rN2ZVkPcB310
MpTJvEdTaNnoGVjNgfq8FsMzcKxwVEJVSqZel1FHWtl2BWdAwj/61Q5JmDPjGoimRtR1GH4Jrsj1
9hfol9mwl2oycUA/30/nC+zWXi/2M3M85ZY6AOe6DqWI6KStLzRHb54nHuCfOjeGo5WB23tL7XK/
tW5l09QF0orXiFG2uO6MkZQkzvkK8f1N+16x0GFOCfZHNQNpXderUi9urEK7SCxamAc8OrrRDguY
StBKKG1OoKYaU5leZ69f0e/dspSiv2ltU+9TG/sw0F8Zd9KZEAQFM3sdmvGqetqPRNzChp7yzpQf
OJj0BvySP2Z3dyBho9klwRkKr4NsLwTYQVtXc4+wuUiBd+AL0QQqmpSdKhyauadHKbKckzEW12B2
UkElAuhqtCeJ9kDy58Yq0875qGb+QqJIfbrHyGIT3wcrRrXJOUepehu0vVc6xRhfH+xlRtWgmWXe
ujiI7oH2Y7423Oa44acpnamglWkcew50bDjuizR/gr3dslXfMbsrMyS/K5vZ+AAToddOFVtCxvwX
DQZsFyH1IvIK1L8fpa2RkbRG0zKH7vaXzrlHZnE5STMgcgDW0qPbSjugKOESMt0ryjvtQPUMhGhQ
NZCNlL22SaGgoILltjVroMEkCoX9ZY9H0XifwqNkoz1R2wQW+4emaAeyuuA7nav0cCmVqMH43u/R
3vEgPSmCwZe2pkoUVyW5O/59R4NP8ZWtprnj+/kse1fNvdttNrHWqUhyxfArZNCzLoWvjVU5Hanp
1rkAcmteMmcHH67gfHBhmPU6vJMf409R29sAkwH9YRG6q9BQoWZPYRRxFQy3U9xx4hDekpUEYFh+
6FasNVeBlQIvCLkOguPjdYgHlJsH2D7jrDjQUjlublBOBCPa6CPOKsRSkqoL6WFCi//3rIk51zz0
DdnQ0YLhJwg4OyKatwJ9TdzbC8tMB6NYohj9EJQGh+zZhRC58p9TekC9oEiXWJKr+PouVNaktPlo
EuT99OLZT+JV+lheQ3p4M+ge0DrwPh/BtmVWjHvTXGnnUoGcrM2OmquruEtzxK2oMCY/uRtODoA+
tQUqJfxYJ4Zxw2pBEu/G4lI2tRIa+FtYNYl8pou8iC+kquaCr0z1FlZR90WRDbV7LdNWr0XKaBBJ
cOCbLP9zRkzdQwRTlHhB5zw4MkSG53F82tkBj04XCc8qB5+IHTrSeMOA7glim48hnT+QhOyPIvOQ
GqDOniEs+z+L/fZOekQ7ol0S2QacqnQ6RFVjIu0hesngVI5tWafgiZnKuOw1Dk3oMMWawxjz0nJe
NBJIgZEojBcid/T+5x+X4xLx71FSeBP41VKEvVwT4Htp5qmjijlaYjlbXVOhQCoetyZuJGgnZus4
fed1QgdjQe+ndqXLxeDGEt0TqbNplz1LL5gOvqQps8VscyNZYZRLL6BENwmmd9nH0aBaAyE/ULjd
MN2FlVqXZvwxACR+gmUR4lMNDwnV+weT1NMWE72s7luZEwrxdi9wMwd/v18Jzh1CIUspGRyTOn3S
/QECt35OlDjUkeEuLmQpiMWwddl2SYaRnP/ymfTXzRQx7KVeOyWqSdYFE3KS3SLUptOuVBgthy2i
Pwhev/0FImc+W1z9Uco/A6h4dfwWSG3w23b6K7fPSQJeMLEI34OglHjYzXtAaUnU/0/8fxttKB8H
fnB4u+kURnEaaJHZ4OLbEKl2hjkJPzj5cSMlddhmalq8/ahjaHgpRjA4VFGmDNFEodVmjB3QXUyP
vou0HugwYsz1IVagltVf7AuSH0rqbNzGEBvj3yASgSozA2QYTyTUB1q8w/6k0KX/a3HD2PzEcWRK
UR66Pddvm4B+YkaflJ1ucttoDhOLokH3YrdU1hWuqh8Flk/7caXUzPYKQXwvrdseoCqz96jo/qQ+
iFpto6e+RGKEDJXqsIzS27No1RUfNo2Dko8gmt3V9OrY9lcnv+2BWfaX15HEqFocVZlIGUlEwVRf
wloD6JuQTb+5NJ8vh6y9m93AhXxqF2g/4pgY70yiq5EHhHel3S1xd8UAuxlmS9tcijPkQMvi8iZe
U4aoDRe2RkZFIucGXmbiTCrm5K2Xtlew5MrA5ptHvn4aRw0y/W2F0tCqxRw8P7YX/CHT9aZ+aYQH
SQK+hoqsDPDHBVU4O5hXrC6g4DXHXyYPK7WMssOLx+NgwuDVN7lvtXm0VFu7EbFB1R9fC0tpp2q5
rReBOjh1+42J6jcTJIHOXWtePpSwybBy9ZIkZMzk14TDRNbtzSh66VEPpzsXnui6haDYW7TGWkS0
FQdCahWM9Kaw77ClOazHS4QtEF+v00wDRzeSRMwxga55YN9lUJCv65iN7Z55Jt+yaeqM41InUchl
S9MLF2gx+ZCgy3WWCzLLDX6X2cdh/K3DmpnbnSDZoTO4ytpQm2m1kKz+U/wumSCBOtMmS15XacR9
CtgJYoyg4hn4dGIGMhGTicWy8k6TyHBFFLmFCrd2gHyYyj4n4R26t1oCzsgjRYD2leZgTLeiSmSj
pg3qN+V+TmLLHHJUDKwHfTI4pjQGuKcmOK+IhENGmMkDfv786HC4nWafHurlaErESaKD5jMrkYDk
wTUZl5Tg1sdW0uzUhGFDnMkDaqGTsB99JocVxNZLmQptVp5lsOqfmauNZQU2Z3q+pLc/PWtymUl9
NBAmMxMIqbZq+zZ1uiW3rpiYfIghe7/j1BFW6sz1ZrczdJ/duo15DF1lnEFwYGS9NdOX6t2Eafc5
FPm/6ExeWnnaeewxzrCCGWmYPSgsZy25lGGDU0LVo+BpT1Zm9nzB7Kb01RtUAsp0KDRHbZQBiea4
DOI123a8BDWLoEAQ4wyvZG28pzE/23A9uC+9jjM258uMdSO4X7a84a4vd+ESDycbdtlbOuPmkbF+
tPofRsfXKUmmWbcMX/QIrBuiwkXAehFlPKU/ERbHQnJAIfuD2QE1R65Lvn6qKU5HIF3OWifChOzt
/2O28Zj6JC4awe7z0PftemWeca/WXvIG4QxQTOSUtWjOdG6tVq2qlpq42ht5y4yzcD6ZlwxrgjrI
haqStLRTHgDQx9TsLaDxeFgUEinEwclnrKnYSTJBanyjl0r/gZr6HKTOziSTxsX4VLl9yr8T8B2G
GxL5iALBMUYRzLcW+9anP9HRjlXoGj0wtlHX8QQ35a8qFiWZd35NtK97JwlNvHryfmz7b5uiAo/q
FDbEcgOzfFz0tOxKKhkYmUiZgph/TxmjD3TZT2tTiwKPPLa8sQuKwoDIl1gWYBdIKTll7X2ei6tW
2uMHZx6TNCminTnLNTkJVZXO3lKZCG+jfMYnOybToNQpOvjMvnNTvWil3s7X1m3S26JBuTVA2O+L
4kjQ8eufIQiWHIupdk7BmDHo7tkFqQFhj9evBNRqtb3BsYy1szpvdu7elCvNkYVi+U2Jlb4wju08
mvZkRmsUG/gRe8r4KndxCgzEohJy4hz4ghv6Q1co2p+bhWSZchtROh87KreNJGrsu8yydXCtoPiS
R3+yXYHVvdRg4BikwU1zcrabMV5xqW9pL6k89hvzPqOf3v0GoxNRWb+0EGY4r7dgInPJ3+RRciEm
86G54lzkZ+pMaO0SGecWXOaAEhY3PdK7httSIvgvm8ZMdPTK8Ktvp47oEC7rGAy2ikmUL4rOIy8j
M6Yd/MuRP78xI+/2Cl5XUykuiuPAl2IH1mqWf21T/VlNKx3fcRSo87cxEmYGI+suF0TyBzYYIgsa
Dgm4+3XJDEUsN9Mf3F1CPdQKnoDqxMpQoeLqp6khIvkfGmiAXlwHfxhwChM6Qj63VVfRDdEdwnZj
Cm8EinOPuf/4cfLeIaTm5+R9g/tzk433E4eHRWeNSj/T1VNWdvGmv8aNFghyNPwg1egkCyqiCU5U
W+e9feuG2ku6P5ufB5JpIJiX+CI9Z/2WtWzw7JmsXsrx1W2rQTz4Pl1n4UE+j8QVeQJ+b+rAQA7A
TDYIhIi/jpIPiLhdEqb5OoUBlmg/jyVIknfJgjVOf9FMbGqgTTPcdgrUQeRgEfMkFwg9Q0u25+bZ
RSmzQAoRIxySsQu4oKfuDIjTFwAKgteVWodmzaE7jYLdp2iEirIc1prfNiiUs5TSSGii5XsYNbk8
+aP+8XK2iS6MZ0xYwmw1ayhWROY6tvJ+sXZFlMj6y70sYAN89TsnvzrvdMpZGVP0k6jZUTTVDHZF
x2+UevIZiVQT4AQpPjJv7/dEkCrFqV/lsPm3oaBbb7U8agGesVb9rRk6N3OzOzoh8eXjwSHVlIBJ
KFtiK6Qf+6go0ZElFa2MebTSvl6wgok0BHSvsyd99Id4tSAlF1aXjVrcGaE/V9OmDSA2ZNAnjWr1
XlM7fEpO3iLXpdMAAoN8v6/dSLDrwM150UEZr7jOE26En1QwDG63r98fSG9WV7i65+VRy+p/TcPz
qJi9GdggdYH7E9Sextm6gcSw3onS7uUDYs8KqPkKZEN+UtnXQZHiXIVGblaMnXFCqbGk49inrvFy
E+tDQ0A7ndBHfcl3r3hmmGOaXvcoNbS9WV1EOg0NPppNiOSGYWKmTtavCJmPtjFe46jhmAZWxdK3
qCVStI7TmzIYKsaD8FGjYIQNbS1mX8lOWqY0bxI0qrbLaqNEgjYaefTNqxXTGrDwj7weihNW92CP
teS47SdKN04zkzaFt9oJwr3PWpuhgmx518BnLVjKrHnm6zv6wpsCRGidr9c0rXQYeFVDbTkOit5V
tdT9bu+ejiRsUj7gbbafVOI8o/rXtIY/BN2XLj21YhzemLLQH1CG6OW28XgpqbuOsJzLrulO7vfs
3/+KJeUTUfv65BRqgB84gTi4g1/QP1OTE5O7K3tEDwhDcSI3y01zNIfDo0ZgYO7OatR7D4k+tXQ3
0KqrDAMampxkFp66i1TN1Ituoa8qw1kX3UiA+KkzIkRs0lYhKlRT+IDvV2xzo7C07w6o9uvFQUCj
WF+JjCYi2igPQIByUipG/5+tTXWlaJOWWSGm+RAAKxJQQc8LejgQvpEfvu25KgPu2H/piK0lWGC1
Fu0GxgmP4QripS6HKmI/r/rsL/RvG9/5eEjatXTUWA/l6fNNP8+5+6Cv3zWVKAsoBpmdDZ4Zok3p
63Uuy0UUmU1zL7KY9neeSAtyl1Xu9yjkq9flm70qbOpI6zK07fe3wOdeorkYFq7ECiEiiiIizPIU
JWNLvtpfodZgO2LVQjTveBSg5r02prorOHK36HzVlMFGHHhESKBRpeIkYMbGBokkCtuIf1KMqY9Z
BLN3NCCXvA1x5sGxJfNOc6W53ej6fUwjFeZabyGJoaOh/NF+Eew5XDJBZgeti/JK//i8pOTMzzPC
nOwEUH1z3Xmtj8qmuRphHm0A5vgaqJnYZm32uXZYNd04lY0RiTOikHdEv/aESSHQOlzqcSREj0fv
h2HuSGOAHHKlaKEiujhA73MbJirpOY/Scn8W6pBhRLlrDyzIGYHrECFpWrAk7uYLrv67Wpdke5Hs
FaU5DgNCUx9libzmZGeq6WfKJgxvb4B/1LdWbmXtFd8gZXNV9XQw+5sXpcQnRhx5pLpUaUV1+O/D
12STQrR1ReT3p+xMSItJfxW0v39bjQ//eGtqTJd4BJPvBCgNQRzXm5YF6dvPFmaGczvcRZFTgDmJ
0H7RNJQDx7Gj82FZexEJRoXZ3EslsRGodqpLfwt0yu2OAlmex5pL3qns4mPcITxslnV6kwdG8KJC
EYJCGtxu2oCvEN/VkDI0taHr8f0KOEzaogg4Yrw06bESAFiPomP4ii9ZWajkcSL3v7lpY+qU1kjb
OFQ/QoNz97XYG/Dluxmejt42hx6o6n30NndCWVA+GtV3Mum8C0kwez+NeTUTtOx/Mw/MMUkFVwKE
6VwZ///uXOriJv1VqX1jKOm2Q4ghqIKtnVajriPtD+p4D+QfvdAnmgKtaIVPMuOj67pFH4nKoz7Z
82VAKkVsHtSj6XoX05odwDBDMg39tKCOq4NsAKoiFR5WZSpy4RTK/2c9paXTHaKez6iybkMu1FTk
agRYY79ZOZBttUoCd2Vne95akiIpW5G9JxjK07MMXpDp5Kt9/NAhk1yGZ941zqNkXG266sWnBKMb
+h/C/FPnVFY/8re2TUKEJ1GmN5b3XSBwXj8Nw9CIVfigZqNoIfzmxqdqnA+6iBVhY53/JmDkm6Ye
JG4nBiaiTQ/r7/6/UbAdu7/JSv2+eNXKpFQaz5Oy4pN8pvoWVWDocAIjl6lP4qg2mi7rfQd1nfxJ
aeoFKLbqQ8a4DOZ8VYMMFE0RZhojpwzZzhDSnDtFcGffXwxj5OorgXrhOn77v7oSnKxZ5eaqG7un
8gOoRYKjOGBj8Jj0WX+wkiEyOxGO4jG131aBGGJxVRzd3VSd9G2nQMfrapb2kRsY0mpLHv1onTU6
tlmNy9w+La4jnMxx4ep5dI9tI53e0urV6zUICfcRKnTEjRQqRZG757HcEhMLXV4aPYpktMYjQBSD
adIMentgG3eMdpN89dYbprrC34+o9bVHVcx49E9NVikc9Q3JSkqzf4QUvufDwCgcMYnAmr27TqlD
SqCC5DnUHXg1skZFEVThQKlOaGXOS3fZB9IqdLFjPZYotrM1elTl5+v/q8A32OGc5cwA+Y3TYGBL
HPJB0ceMKqBrZ6dWDPISe94kUtYw1U/OtTopbXvMLEIJ1AB4MgdjraeJxPfsbJEdCSJHLy1uLFfM
atxSP3xVQhtqALWur6YatSTSbDZjYyWFiri+GWY++tjkgBXd+vsujqEB84OoQbl6tjcRexqHAvSG
jFWjG10mP5Df9PHKwcTM3RxXEpKFbIgViScNvh+7uolTfdcVZ2t8W3ev07HSjGPJV2ium7f3+Taf
l1WxSAcwmUVLSGjwpHAKUW/EWBpBDKsRlvfCPKU3nbzJFl2qeFFLjhYsISkcn43TNiDj+Qx++U3b
8DzlpkihSoh2/EFs5NP4WhVtTxfFqxhusw9zJVo51VIFmrmBSk+U8Grcs9CEfgypXoq1K9uaMSLT
PTHgAOZvUJfq5sttza+mL0qCgpL2kfcmnD23Nz8yYuMccqlYT++BkDy33QdWM7bZl0g6HLeHCS1K
KrCAInymNQFYJXikQ8rmzbr71dkwD66uSDJzQWpDrkmSBpmlhWD57ZWGSAHNIstbvsOaRS3Q8p+f
PRpZLhs485dgzJ8sZUl51TEMJG5zjna8f2uLMe7wXZk1+R2aVkSGA3dL4WgRAM3Mr/DsrXvejWsU
Trv7F7zsYD0xxDcqI+lxcg9D0GPsxppiLNuX/g0CDwk/KhM7QrI3QNBxjpJLFGDtX4fj/PNf3abd
sVwcwKHICL296tFmtL+I/MZJ+ZxmpHJUhYu1V7TAY8zXzYEvkpuYClv7ElZYYN8wJXoApCftY+LT
zoFu49Q4WZ6CC/9G7XnvQ1tR8w4GJgU3yx6lvo3Ed0s2H9A45iks/Ixm0ZBueOrXnKhzBjvuqS/e
F0mhpKKIxRwCpqzmYgLL5oR8m316yOD0Nnef9NZ9nclQP4fKg1w1SXIPtvJjLKKHVU5oaJAb2pX9
kNtwXJl6VqWekQaIRFFIWd1o56b0JUiL6FrpIhxz9R3P7MfkptsDKWO/zsAJJS3VVKfYP80TvoTo
3WOwnVz2/im39erNOnCkH48ra7C30xkMatnwurV6JZEgF1ByBuPXiFqGighAi48cIgC+ZtUXj6JS
t4TZzdKZ5nsbfMyq9U8IBsaXEl7W5XbYE/Ny4J8oaxVygS8+wb5UgSxqDLn0QQt/HrhsIxEUNDlB
kEXAxBKwuLqOrni6XE9g7ZpjaH2Pn6S5m9LZdVHERbxLa1ANdwNz0OCRbULzNO5lS0BAq64HMvKw
sIsZK11QjX1ZzL/1g4ct1DVvQi5k0aSrESZdP3qkTCjusSGAZHk54U75AoSaa5G9fXfrwd35AHxN
SO/PtCh5A/CDgbB2MmJo0RHSS/zs4J7Cay3XhFFdIe6bNwRQNcy1uTBEMnXysFVFAtK+ps4FN+eo
m6GApxyFEKu+kvBzs9gq2iqb38KpsDNgBQy554STBwRmLLFpJhoMp+yatKZG7fpi1/qYzdMQXE3o
tyShFFlm0GX1+eb8GbYd/Jru4KInGrEMDyZ/InFWnfqUbezUugH/1TZz5hO+Q7K3d5R5sK5l4UYK
zOG2y/ZlFlJJQgWabOg6XTWeIsVlvvm8YyMRo8yQuaFCYTuWYwM+un/W0tgWJIBG9OF/vWczSKoC
fmsenknl6uKydamgGtN9yDwULlA1pMftGoaJJyZ6xSo0bjbCTz7EQKBjql+tdSB/w8ERL3O7YJ7n
FIUQ6eiVmquvm/SX77MGdN9neIIUsqHKWc8M/jXhZK+ARJyne5ZRii/vvJtQfBRIXUpqDYYQQKDZ
uEtE3WtgTURFpmQlCxIcmdKAq90NVfvZ2o9aYUYVZPCAj0A+Wp9YBdeU6S1oRnrJPFSelhIRUrI0
pKQTQ+WGpXDMf0UJURH0+VfTzgFixkAsEDyR7LzTIniM6Wr31Xh16FcjfRGZ/l4QIgK84EfT0O/J
oPl6aYweE7B/sn3lR8ZEYmhzOtRmMuyqiuu0aHJ5xc25UP21UChPy9mvX8+HusYOWz2ZbI3Q8dLB
IcwdDhyCWVJyGuw9Joc9ZFODjAc7og8j/ChAaDuMonfRjsfT4AoS2lBMPKWL0X8z4mYfN3ECRhPv
ntInl3F9Tn89PM6hcWxHYv3uh6pnpibx+nL/T/+Rba5xMRVE3uJCoisndtIpW4hNL92hpU+bnmk5
7wJi5yRhMqiXvVc/xz67l5SE58jHVCp6V7ZzgvNImtzjoWPetEGkdNyOmq4Qkjdn8yCxHyoRK8Yx
63ToHYxouD2X4kb78kNcnfhqq98rgdmSj4NUigG7rH0LPjVf26dIkbQkM5BNbVctK1Az7D2f0p6T
HcaL6VqL914GkSA+wfBiZYHZNNZ0NIsshYZlSST8UhPWlz+F4JfgrjfsQ41cgy9j6i9Qs5wg5vsz
FTr3u2eJ/TWW0gFZbDd2jHuWL4ldk99PIafkgHo0877osZkNAMSkEvZNGPV6AKMTdJYRkxRpwM1b
4chWZIcmJdubUP8HXehAIOldNd5PBhBqP5lihFbiQOvOcrbd+GSRu5xaHmYF7za+KBRegLMIa86w
R1FI7y3R630+2PtSmwdutKr/m8fD7Se/GR4yX9z7hpOX3G3wYyR/3cvqVYBI4JfHBLKwE5HCrJ9G
gxP4s0+HmeA2gul3iK4e5eK8scv4auIQIwKhgmm5tvRQRmhKAjwnPDM8D+AV5NHi+sT57rex06i6
KwJlqi7UXbNyGrGAmDspWborItCNAoH5+RKOLcbCJWVBx6EZpib5sAdf85aW37Iv3ytKkQ7PjF4I
u6isNbF6svcDmKg3mMc1a8oFN2sFt20i8rDiWnm1bxVzZJq54GvtnE2WCZ/UpDaDpNJ+HloNSR1z
FFZu2ZqX6sHPLqk+tUgjK02jg8VBwYNX9eNgzY1hRbQ4p4v4YuSx42BOjoNXYB7TTDztu++mK85q
mWZdQCwRQg+AiMErCraIE1hLsOavV83PA++mPPZSUN4gAq2tmp/SctjlgwK77TjPIPmgxiVkQDhM
zklk8x8vImMUk2lzfDvMFjehC4/C0mp+r+lPwYSCp+xznUpeYXkGh76iAYIb7Zt8BAzJvlDgWPm1
GoeanzIqEJE3wopaFdf0zmzcXxeznqpoe9WcU/IoMcGrIcZ4Qgbs3oo+3xnY++23arAOmNjg6fMR
6/b4j1auKsOK5EMad0mAYJTE67/EVh1rIMTACEPJP3m5jHO3Aa/MBzdUXyu1tQ638YE8G2VTfgXp
cqte81jG2pfyJN3yD7uQRuxsYX9wf/UrIrQBMTKojlmDOk8EIQCRZ1O9P4r19RwLPOn1WTp39Nqr
8P+FhKK7ZccX3qekKRIvdTmhpWFT4Mz6oAMuVVS9qGN5SrFZa/k99WQ7hakWqP3rPdR0+xKuNtbM
ed9NZp+wrA+/bKqPfjDJHI243lOJ3SNo6kzT0MEixANxB9qRiBVpE+O1Vt7OBvkmj76Ld117F/Ag
csEqZVHT9ePWfWDbu2oGDXbOef3jkx1QaT+eH/rFotqlLMCZltpFUQ8WR3MSVM6QTFRU8ZDdIErB
PPgTqeEEYY6rNzT33cd8x70KM5BgPgtdoL9gbd+pCBoamxx4DtST4S0dBASuEJ/3Cu5x0iNb7DPM
apewHKutLQ/djdoiE8IwZm8xAmfn0BU2j6BSCMuPfRQY5Bnbv/irp6kL/z5MxPgBlSKoqi2VOnfV
Dy4qs13ywy8HGRQalfhWAp4Y0iAv3EtSWJq08ET+d8fEQOHDi2VPXtieNHVIkHxsd7IwKMo2tQR2
aRZos/ltqrE/cL/r6jACMRFD1A/o9JbG9POS6qL/lVX3E3yO9ni/zeNt1w486m0CZjjAmYVA8XmV
6rkOdHt+ylvz6yGGbbWspSwekWRhnIjbaovKOSFQQUqSQJ/3ERD2y8liw7hUc40VC9zID2UxCf8l
Zqf6u7S9+7yc4kR+i9h6yhb10D7yuzOyojlhE6GWJKf7DE2743MvIwXrAIa7Q9gwO5/t0lxYSiP4
v/KS/YK0nghDW8HRjbIHWsDXBebg5sEQlXXrrfwwwgCxYVdx/CxNUNtaTDfqNo319jYGswEyGC60
XySKiq8xf95QKphVXbFfalTw9bJutAOt8r52mctDnOlm557Inirit5JhUwR9zIjjr/nsdUak+CVv
+T9oMCR0hwzeYNmDrosRZaFsq3ty/px1P4Mdypfme7QpKcy1FqPOPZoKU/7V1X2fNooeZBWo+HnJ
PQk1deSFa4ELi+mMs3jRt8J/QxLtXruZZGz8K9228UlZzIDEvgJdkZQjXWZ//RRskcQfBJJGdj+v
bLTd/cOtc1QQEkLHnD0e5LomdLckES5dVW4GA9HArDxsnGbkUS+ZPa54VliLl1B/GwXey0rPhxPT
hz8+plXKoaN4VBJl873KmpGSpP8AK8lQOwaTrSxVKtFanlQzXDK2JsmdkrLjIWVJvlfPLb2xW5Ll
nQSCqb1WjPwnulBdQkVBPldjaMq8PgBB+nr5+2u3kRb9XXADGQ799rPmbj1Av9Cl9EwsiCKWr1kz
7IrYs3mCO4FQEzaFyj3CRNhyBrc8KM5f71C6qrhJt1WADx2FzW6Pbam2skMixW0RCW+ZgEjikddM
UNFXam1Hp5jZhQxCXmIsf7kNhyF24rNbta5aXLPNGx2ayIlCj4I43R/CyT3lzsrLx3GYjPRAVCmq
aEwc3HsMMplEm/+zQKm5fenhpJcFNuaBDGfnXOVX+Mjfn6YP8qztYUHI7E53po6M0airXYvAZcA4
6ZieC5CTER7NIFnjhZU4CmwBzD6bat02isLgHGGwuFwG2qg37JnBLdoPdIuVrZ9kgdTgpOYxL4rp
6Lup5YnUv9NVSWH603bNdXo11TMVTrDE7hVXuU1gLU3vr0bNjq2WGdJSAfmOLs28VznmHGlzbTtN
9iKyhAJ5M/v3/mxkxtW1RDWTJ3oJ3kpiTae6o+Bh/n+DYnS8b03XUVP66j4/zPhYQn3bHETLRgsE
QBEvq1lTy6fwdGVDCNbZFrd7nWeLlRxZxPKt9pdV6kcYqxeSDx91Xj7UxQW+Vk2EpunOnzhTS/Y1
TxunPG3i5KEG1Kj0nBRy5+gPA5ifF03UnitBmNfC8D0oK8GPah8iBgm/kDOU7URjTDoA7AfM99bq
OK6crSnUrE247OLWTU76qAHu9onp0MlulXTQ7YaI4v3YTe5vNLJkmHgA8I3gIYAabc2Sbdzk1K6Z
6Ow4THeL8w1USwWPSXwelKW7fSYj02AuoHDpkF0L4hXBAPs28s9J1g5zUBrIKKeU0BRwRUAs9pcf
FVu1ooqvJIpnD0P6krWupSKI9NH51ZdUERIGUMhaGnt2rkhiburYc5UMVJ1+Okd6ZiKQDAPmTM4n
OCrfUkqGWUNosxJs6z36NHPgFwXAyYm968Hb7GkIrIeVjiw9m56ffhYz59Dmb6LcyrOIUKsKNI2J
lY/CoitrSmrsRyKrQXPS/P1xc0zGqqbNEUyQSeFIBTOgrSTKOV4m0fsfnO5L1Ax5T95IbHVK3fKH
n5CZpBK0n9ykkt30yjzDxlN3S8i1j3p6Bs4B33SCuHEDok6wwd96HPWEQMcYSk1oxuSQo5OENc66
vzKpY9G+EfKBxOK30paJJH7NS+HAYhO2JRBBgnnzzCaKttI4nFVlKRyitnG8stklFzwl1qRBs3iF
NNjhF78yH8tqeCF5jSYAW4nOSKIf5f9Bl1GY3xS44wpjuOgnlfYioDgUkpDWsf3xElgq1KNEey7l
SnQHUeXib90E87d5zbkc3wBdpCIv2pMNE8qkqfrBW7RrKN4pWdx3T1PIk7Gy+q7KjdGTd8K+YYr8
mAGzHS+APHe5dAEWwYEt/OxzbHk/sEoNpoaqHB2LawQd3qTzlWiJBpyscks8z06nU+N27A0iFVfP
DV6MgsTurPrxuzXMaZCdUoxPcvgZu2ovnBgR5i2CmQrMFMfPpRhxiocSvZR/CH4gMRn5fIZHzkjG
EwmU6TNJ7PVSg0JS1ezZkTONgIQB5YcsyFYc45SzJwHxNgcK0C1DiJzAi6J30wXNnyby7C73fhuk
vfPB/esaGBgYoeUUDi36wKrAsbWSOt3efLhAJdh3lMNVQsqh0jk9FJim/qlM6JHfhSwBSdEpY3PV
F7YMGa/IUT40Zlpy/lHnIHTOMXyqSUdolLV7nSrT7KOhABL7AtGubAAfl3X2O89zfKOZQYetJA1r
wPoHrka4G9+omrusXtkauKV9wwSdgR500WFMZ5tBRdlr2IBxEzU+qwEweJfFZwjRK4z/nbGLUosi
Fvxw2NM89W3iB1ev99dRO8PrNfspsnv3FxZVINiBat4Zu7dQZ9pR7hMp9AdEei09dwuQWUusHCUS
EEgDbGA77i5cFpVMfm0AS+IDEY/dp1J7JJ8I/7qBtB0/JZDjmxH2PY68U7nxCyqrevFSWeNfw9w6
Zxi96C4mL+JwD5OGi/lmZXZGPnWJD1293Bz0IZt2kjzYBJTJB/fHu6ZY1HI6nLLnNVmyq1gOvsXl
sYtwKMgKQ8xvnW4G7hCM1brgVUlSpMev4yzlPvHKT2R8qN7jowIy3xHY1sqWl1F5QqFGCq+iQuwL
uyrLzrZDIh9mjbMrK80ZLygIySUI36it783tfaObhDj/YTJ/1Q02ob9P0SzREGxQvFDECTjBocZs
qwVGpsLtGBkYvZqwPx4DnVmTiXoQ9B6mODnjyB8QO4qQfJaOBD4mmgB27f9vIhhujMSybmW8UAP2
tsbdU34ccoDj5B03mA63wLs/OMZxYT3a4q7GM+z50nqsOPsNWg/S0vdfhHhJSR2b0NLx8iDXhnVZ
DuulZvLjcftl6u5Yhurq1XM1Wen6JxqxrnHqPS0E05sZOu5JcmoT/7oRb78Wa7bEL0NRy0lYv2W+
SduNZ2GwnmR4t5ues54Rzvc4stK7qeWYZJ389eRQC9Px+yDG0x2NpCtdvvKp/L7N73s5WQmik3Ba
vfdB4apiLX0XrubA1Uq0PvF1gbpKNOF/ITHC++gu3NV/qJI1yVTOvn6i1HK/07oYIDeDOY8au4pe
+piVKbfDwCdrJY7FQi/n1pviOMFCDO1AGoC4gJGDFwxuxIpI6Qcqz7NH8s8Wuqx5rCYnA4Wf4Rvq
4SYiiuPI68J8ab1JjJG28NXmQB9hl+VqFoJZvCn/i2wt1v+sAmGqk0KS4ezat2SfdM8uJXPTcpmu
6L+dmSI3vN6SQHd7FPViRlC/hCVGsXFfYobfcgV/QQ7gItbH2zTC3vpA0qirERQc0ae30vkEp9lb
EnJ/DG2Yl3aRTIUVqfwAc9lQbVDkr6+1tErK0giMk3CCw6VuGsp1558FoVGTigSiB/OwWMhUqpAt
VDJo+hp2QcbWwzDY4frzjrt6PsuhexHsXjOUqNJ4uvkaBJB1jFwEjPLU3JTeOsTuL3QbLSa92RAJ
H250XNiFcQcSf+lQHqztoABoTeqFY+WqXq29wPEhHRTSBvONDfv2hQsJE+RiSGdeAZpvdHl1dS1C
F86w14j+3vQiwQGNf43AZz3UigV51civ854QJwN0IDXDw0XD/yEiHOYPzXC8GC+Y+fMuGx4JGWkc
ueBYBYh9J7oPZEYnxgBO+qsoUeHMPTSBELwfZfucYeszMjm85VuKcWSG5EEWeL7UoiPN6Q79e0OD
q8jG1DtquEycg5TfdMWO6Es4Yfb6UWGTn/WE8WEpkAGGGPDI56txoaoGDjsbnS/zhLzBHCg9skDR
kBejHEMv3U+6auxC8xqevePQGlLYl63iGRUNgFIMpzrP1nmQu4D04CIuiWo/wUWFTsBP7d6IYqI3
FM4ZPIKRrBGjzkIL4jn2LAnlQbYKpXoiKip8YeWX2LXo9bo5Nuk+EPrn4vL1frcsRAn3ANttC+fz
50hBEtUpJitwHKhiMji/3U1sDeRv7+sS7mGNQDCriwiXEWkGayI78N9IfX3R9/IOHq+FmNOwpqrN
zd+iJ97/B+6nVoC1giZBRSPtp+F9vDeZOHrSv7TXPKm5hRFSCHXFWizHrs+Lm6LvfBQahZcQlrvp
1+/aWtI9h14LURB9vkjHDH0lQqqJTSeo9ZW4JaqqdpBuEnpsVPrQqNynHCPOZeCqj5NTZQrotWZo
87JemorRC3txXqg5kFR7nA+3Xcxu4wJbrcPSdtw3vjSKTgnsBR4/WsXrEQRLkfFWpCAePLb8nwuT
1HK7MnXMVl/rEcJByhRFZDMsi+3d5SOOH3MOyU6vDKILxiHfsMspJx7Oa2VBfoX5tO32KyLJdtRd
e8AbPWV/l2ciydWFy0rGtUC3fjGiLxogNtoUs9BXtIZgX8trKsOuDvcsgEYT45qeX2RQ1IHQLCz4
EPO0z4hc7SsUnz9SA/b7TZn2m4ZFuipCuNbZm+tf8nbKXnmXN0FRfYgKe2M1/njz6RBjRpT3wPFw
MShEXPiImvVfsHmPqxVyhgHEPhZk0XsBYNi9uvqoWuBaDJT0dsjY+gTPBMe5TwUwCIrp0q3Drm4s
c9gzAUgSP9QOXvWePCA0clS8Lw+Tnb/fxXh6otDrBp2i/JxY9d+ian9rfVWjayUmufV9fM8rJ0bX
FeQFfcWtlIAbCcldNPEBRZtJKd9T9s+OL5pq36Hf+7+vp7UJqERRKjNi9sOh/EDQnYSVU7wR/ugJ
kWbrhS1MhAoIcmOOA3GkHLSPGy5dct8AFRk6VT8SLCDxaE0Arq5H1a+p2aGtlG4OcSBJM7mKF9ub
EYWritruoveV26deXFXVO6WVRszS/a9nL96WK4Ko8j7PlX6H8K1llKkzHT9xMshh09yHN5ZAJSaz
gopO4LBEPsBaHbh8qChis/PvVUGbA2VQmmjSt4p0jCXqoTUi+xfaGublGWnWbQVEtdtjI63DxGu9
1Gx2/R2OCiyJDkuUvm+874kzxQ1aRvscal2OUDHs52N//eK8fvLFQR6rUmOXT8JLtTLcNunEwtXA
VkcnihhjwyPQn+4zaJ4BPntmY/eyGiqbd9BcL9LNlAY37o9MC0WrX8Pr6LvUmNUaR44BainmYxOO
QVvDn7N0Ud1c6XHCl6L0f/tDfU1qkDDprQD/LJcOLlRw07BnoCypXWju1G+iDOkQGe8cWydjw/MW
rt7TUqGglDw285gagdHApjGRlmV+lnKmyoulcUtPv9f4iLH7/Y3gMfZvJTYLT56LDYdFqhzCa5Ns
Pwn8eu8W/SiqYE410Q6qv9qdQ2Y7nY9/o9kEqeVT4PLKC/nMUWikiTDpczqledNXbcVe7nNKpTgp
EDrZPqT6hMH85cAWl+Jf02uSy/JjSe6ZjEteN2h6p7roMGhjLs/5SpXoS0JdgNtDGSexy1vHlwyK
wqne0e1gLKUc4LvucVWKDaYsegZSyZuJXP1usImDxQQEMOH3UuoxD9Jbd7tNV96oHsW4IMFXuGHf
1LAzgUH5LDRVnN78yUXHOzu0VDrHS5NyxQU1DWcTFvr44vJLQplFi0phXLhD7H41kt2azhRlqnEj
F/LxaDtqwyMNB30mJKARP/IexEpsnGn6tksee1qQzJuQF2QtnjeLp3+4uR6Yd4l2zNw/FijK43Fa
1tpRWBU7z2O2R96cCBu7vi2DspduWkFSzFEzSL0dVWrcg7Q3eG7MyAOBT9D9pJcmTqrIHLfta8bH
yh6bM1/CrNJL3ZOYQITjvUcM8xFReiUsVfFLPnM4z4j5M6VefITw/YjR2rN1VygaC+zWbH6WNNlT
MbyC/kjv1aMpBduZYlpYylt4Z4r+gfQmn+2u3Cwwdy3MYLgVKDigESxqtDDdP/extRA0E57B+MUb
YXpvbKw0oUA2f1gltV/tmXei5+8NMfDb3Z+d3UlpghVhYInNuO0M425ZgEtdJS6AcZVMGW6rDjBM
QixcOW8CMWf1AmbVfgANaAwZpXR1KwuWOBgf8rmooRETCyDlThDAHks+JBgoB4dTGLG0QfDK0QIO
/4aHTRn6aIHU647lXwMsDZmOaRO1cFuTlkMZ/fxvyVJALyGoCN2sNCgUQ9d5EV5UHpQv/iJNeSe5
qFODAYAbMTaYSJwnjEjAHL/d5QrYlX4zUjkpzKltrcEjorDiuhASW2YDQH8XThMnSKr0myVW9TCN
IY7z2IAp3U6dVlecHNrvKqWUUAefRczE7oV+uZTBV/tQpFh4yV7sV3skRT129qfyBVetohi09Rtw
iACqdjDLT7PhzaKCIelryonXMddqViVDphF6Be6SaXEgKIWeTn7PmS2cYBks3SRfHS4zr8cTzWhE
y0jGGy23rhe/nSOUMWC4Z+ZajFDZFgvnfJQtIzkLW8s2ZU4foxNrzV9s4pk/42Taf5FTEspu+h/2
hOkoBuEOlxigC5h1oHrtF0XSCgqHzi9p29anevnnMQhEXByuxxTwyXGKAs4ZKqf0pTyF3YZZlYMa
FounH1W8yDQlA169UsDauXXyn/M1fN3OvaxGvy0c8imOofbyZ/9weFtARfWm1Wst0vYq0QB9B0Rs
yZfp9jI3V/PzMh0FMFWSoeHLgN34vIQ1XGPUC4Wn9JgEelSaAtTWgnbPnolX2xt9J2yuW9KMDhlu
LHgg9jdUH4Sd1ocS4W2bf1nQTXqh3U2vSSmXj51O/fP4zPZrWGG9wO04yIVZ6FkklyLIsV3emQu3
Amb8zW8FP2jw8Es7IJ13cha1aJGwj+6ix/H65FriGPR3OEibyBfm0hjMFCdy0q2LQEGoLRf8naN2
GvGWKmNTSQm5Mz8dSF8007FgUInPMSRy5Y0/diLx3jFHSeanaFEOZ+Mc8mnDWBocOLxYrUsdsJVY
h1pEqTNyfJWQmS8EieTDVuP5FcMXBm6hx78gG00zlnLgZ/kX0joQQnsDO+AIJ0Tqo7Fpa64OOmXN
7s/JIOCdIGwz1EE6dc7njyXzmK9X3EuzEdAsvKhds4mZ1+5qvm9iWqRb0IJ7fLAvWslXinyP9dfj
qEoZfEZHjPwGuKjo9Vwy6P95ujqm0jPTwlG/gmBinqBnehK0ulHFRTXOor/nq9ZIJNP18kfj+BjO
l+11VjWOy5a9TY7iNUPjEymG4sOqeFRALUSx0OTYD/lB3H0VLVJRQ88QswgZ52c5YjHB7IRQ+gVo
NVffiuTxqiWnJ9MQpSKhbSGS1Tn44tV6sg8O9i/xUTSrBf8D478ky+mzLwkYNjGctSwpS/CGxh1s
usgn6BUghhbSPycgUmt7O5k/bMnIzHe7UUBKk/ycnekfdvz0SKsQ4Z8UBfN2KI4KqiAFxUWEbkYv
JV3g9A5+6Vh1rGFJuCiNV25j0RBtM/ImMr+EDGscdITjH6y6THGGf6kNyvWNdxyPnIfjwEq356aF
WiTuUHT8V5J3xShnHUjzz+ScGcnQMrMnEp6+3y+JSpuDcaOZtWv5MUKb/+pxAjA09cXsREfXdk0V
9KXjWfjH9X1a5uEmFqjhr2NnDGcm9vIMB2q7GuLjWjJCFCkdc4GmdheYvHC/TGy12ZcgeRL8jYZ8
+H82iXzhLUHgKe2RDR6dHs8oQdh35G0a4ycx8eD1u4rfRmAfYKz9LnDA6Gxp90cRXJkaqLtS3fXK
Mc860IaT7bizAFfKHVHznlMG2lWe/vZQTTLsFToSmgSKxWNP7wsNZsUlwkXfWzJSSldAAacjVwE8
crwW8yPEGL6Wh73pKkF6ssDRjSukMgWtjueclQZYvy1SOawjfdvteTi2QKbzxqxdhbt606jNvxfe
FYbYiky0IGb28o0v9Koybr0MxMQaaXXCwntWbdRJJjbhxQuhkxUN9Z9BSs+qQOQ8REQl7q6CJcrb
a+lmWny9/z6LZbV2ih50yUDLTu8JpnsCgGdQIgK3cL+GP9qld1XY50w1rum7MefVxPtLw5sqPkJz
GnuVdwHdn6vzaMybTH6ARgPUFnK/1+57uJUMsZ7/H8CE9KE4cWKyPVIQrlXh9U8grjn9lyNPCoCl
8nCetQ65YLseYJtdeApoWzgPXJh95TkxsaghNtGVcdCd7uPcmWNKlIN8YX5auVxF0zVuIjW9gUng
PyJVBw56rZO1a4Cjfvd3shOAZr3JIOQC3avAJ+r9JwQ/CMNeWMqAeKQmEHlqnzHmDYbKjb5FAtJ/
UiB32VMRYAo3MC18cTgOrxxVqLmQl0oXK5P+JV8uisfMzZl6f7tKgjDmddr1pssx4mYZ5uh1Wojp
HbKgNbJ8o4f40Z474A3J1SdcwJU3I1c/BD1WGeLpsAPVjoaVCtzLuz3J82twwlye8qNZ8g71G0IW
PsGyY0xMLy0emrkogG36RrwGvFMcrklv6Nv0KmQlvQRr8LpwrdmFTaFMZTyE+h97IVeE+ar2L4Zi
LU2WwrICLTa0aH4gT6Dr8XeTQ9jOW4U8FsCvs2YI+iT/RUNaUH1lw7O4eIZZGMqTnXM9Pr+fxFfg
+Tm/dP8qHGSs+jqFQzcjuDGbAA0UTCzD/WmfJEJjzN4GiCbOISeqcOhS2G2DCsZa2AtirKU4Nh9I
ztLizcOpwYjFNCPGWn4LDpB95PvxyuMKRlXn6m7dmcWlRHhsAbsEyEmUG2jcjZxAx5uM75RfbTE9
eGwqt1cZ3WG9SKhGVm52HRHL7RNu72BUyw7kazyTQEYOp6Ay1sPB0Auxf24pytFN/3tKnMw/bCTy
2j9cCzCb/V5LBN6ZL7kBEsZx7k1ITbbnj+WIUl7GvlxEUamF4jw9c6KSKnyjjh7+WZKP6tSTke3F
BwHOOnwJATdmdB1F9lMgzaRLuCHGl4K4FsdBF/OQ2EjlAdIvNWjmO9GvdifdbzEizY5k7T1NlNYe
AiVQ8/HTNNHAcYaMESDK5wcb2MHc2AJVSs2QzosYO/ALolF071d+lNJa+Zv+xg/Epvp1WPgFlUBf
eNgksTWplmmymuSHqWnxXEr39LJgtbZH8unSC6X2S4YEY6zH9QHopIVWNUVnmltw0Yq9Df0vhgG/
7u1ARn7Sh8TWbgu0Rf7h0jsdvZd6iWXXFv6WLzmtpL9V19fCqbRUW9rDd1okIVMZZ00gcQEfB3bW
0SFGRY3GKfR/NMEi9PSbVs2dK5J59BdqCCnel+O4U298KyBQ6zxtXI6siPb3DWj26v8bkFVtfJrc
olEK7/Ey44uaXYbfEe5lpYikhlbvIk3QPKdfoZ9YcdbfFOEWU8R/YjymLrGnp0xstyBks4hQ9rib
F0SYJNNLevXmeVrJQL9Ofy0e/R7Yw5xAuDwrhw/ASG1nsCzDZZvIl5G8ioYHYZi2KbgQQJOKN/wD
FOHapLFIaTXID48Ho8low2nSAsrhykqyubNkekE3A8ne5B3eLjpSKiWs+M/lVXl3lF2K8D3aBI69
RbUcbJlTEOGCnSi2SU427T/pbRDv3f4ppw5H1VtmW8LT8ACsX6v1VXk+gzLC3RJz9/BEjyuJATqj
l2zF+tTEsKaIgWjER0I45zRADZ9lKiJJLzrzIi7S1L+ZWOXwi+TdISPnSv2MrD9NQlrlsV969Wxx
GWx6KVXffXR9UXZmJcZZ6vpPG2VbKrarmG/XyKqJEWH6eOAgEE+74IDm/2KHZMxetGmL4toXfjJG
IUIJa2XLlbzeWk7Rg+4WHpfBZ8Y4lsntljrFGm4ylIXtoHbN6I6VEhw7Uq1LVvgF1euuHKvl9zzM
BwSHcNmrcI7Xc9HnK71N2mLpa7M4W4QvSHa3V/+u07PZ10RYVHPvTN6ThC/15DKasXIryskF2hme
CwYL3b4pLBXG13uwU4Tm+5gl0bOggpr/SREq/yqKfPBSJY2deFWIWbYp5y+3Nkd5qN+M8Ju2nNrU
6S0qnlxOUWOSHT1eyDQapP3p8N5hNiUrls3WZs9hUmvl/BYYX+FSPH1tjmMTDWlVi2Sq7aRQMAjj
5sk/hIu5dqRCTH2xdJLWlDaYgAscEqZdVDy4Q9Xo6OtINabUQ2gm8dJeZZB4AyPBzclF+OWERVPa
dDyfykoSYlyRnaO/Zop5a24HxDrOPJqxx1P4mUI5DY461W+J0H71k8pyIhR8mXD70+fgN7aa1Hjg
oi3vGcGo+OQQn0iOyeG4A2YLi0YSfk6TmIeDpVdF4WGO7cagSVjMN61T+vahSc0ZAcnSvXEDUKPj
PtVb2aydBltLYUypVuDuJ9E46qEvtG/Qnl+JGv3iu+yeljsoqVr4w3ZUUDrK905RwuCrUeKfORK9
Uidq1GHk6/ejDkhsGKnO1AF1MdR3DtF4SNshvQCX2BA+keTHpImKMlFd3IybGtaWxQvGUHW5Iv2l
jVZM86ZWU0ps+3dYkSzD7bfx3ndOFD8Jt9yx30DgbJzxaGfrMaRtx0IJorxHOuzzqnIYiKBbti9/
rOY8nY2VX7XZU8WBONZjeDcHMen67iuBMGNx1FN4UXdQJn+MB6Ytw8+Qhxh9G3WdEl7tuK1nJuNw
c4FYZsoBsS+rqu+ahMcFlDK9aCGlhcKTU8Fhx9AZfy+BgJXCswEZJyrhEFW15oSXSUohtc1tOAvi
/ezMF3wCyuh489pp8+hzlsxvdPad4cUjArF7RphT8qkGKqbJI1/w84aySuJJnDw33oG2H5Dd/YWC
EDp+uVBB9XQNvc9uqsMglc6cD3yFFc7fHUy6dOMNMpmwDwODViN+ivIpIshQ33m1caJkluYdZfBB
x6rOfzkqQcMhK5ValUNb0iS/oUjFyLjtQ9JarJrxYNtZaKrqyDvQYeZ6eOkk+kiuL8rXnkdRHbMU
rBALFnUJDKda4Cbtr71Pm/4OlB2tTHXmLUHaQ/ezoiSJYuU9MnDm+8HKu8Su+TTjOuY1ZPQbyZan
1mggrxTxJsF0toE1uQ49Qsj59RV06YKNuyBsuJkhmODA5JDPm8++c/7U9VotfGVDP9jYDlEvYTE6
5HXeeW+9og4dcfX5IuI446SG14ra6SLzb0jJMOcX5Dbtmwa1NbbrHNAz7s2bmBm3Ys+y56AP/uia
rL9pvc7PaM38xtIpBlmcCxr0WJ4hhy5xCm7RA0QWDQRFH9NmIGObupu5afkJoZ583rbn04nrtSRp
yRXt7zIR7wIqQZdmy0ymGXdPBscmX0TA9S6vBvmXYFzk/AnS2f32W9ZsyH4GBPFckA8W4KYNXHRv
keWlkKG652OxWwE8FPyyP5Hh8nD1/JZpel3zj10QDGZQ3OWx5dSVVon+L0/Dd5MKP+LfNA00JWrY
FACCqxePLyb6mKueNqSHPNUmUY6s4w0AYj63A49XsCiqQwPx6Lmaj4qZB8cmvgJ+G4q9GIobNWrm
NdukQ1EzYZqsZhlWkosaW8wSoBlYOQINQSgqwVizj82rKGq4zZT0U4R4hvCeLLttCqszKd37WSZJ
Cmu1UdzYff53wUo8widvnO1hWLnd4gqOFuZ6sjQpe6IuPWy4mf1BlGQNVDZpIDJ+G+JQASGnphYh
6TeUM3H7/Owr7AnpG486DoWChgLFYGfNejAYIdrRxewr+Pk4uRFQOurLIkFW2tMCm5JZIhNPgvh4
CEHsDXcKn2thR4jS5FsSxpXhA9rlTzoniFQtF/Hh3mvvSsgLK6tRTs8CdBmR0590ZTzQyJlMYJrb
inJxLEIKy/DAkjaEOWHErl+Gb1dLq00fyyOLkiJCZlYghG3+ZvuvBRABOhsXmCCi+JFJGbmjeW8U
q54MX5mLsDvtbBL6ChNDwPYlpGBy+eXHxUYmEo90yguS89NEypJbDQcZXVJ0u8UVnXLb09Q2iZ7e
R2Upe/Vd8z1uPSvpe1nD/ZvSTAVtLU+iPA3/cI1h9VmNhRSnzKbJRtu5uC6F+wYRjpaXm1Wky1LL
KTvvJXfcBwgj2CdN1lmxx3XC/ZttCYQgAFK3AQsJzKE2L//J3IeMAA0skDUZbBN8GMhQ+iC2Mdnh
J7Rur8hZktXUjhahUzHgWeHDAmWgu6jRJLwMFuxoUfI0VrAafAqXywvwtMVu6s2YQFo0BU3TA2Fx
xLFrGjda6N/MXm39ABVKfNUKCSDrs1RXkga+jxhC/Vv5pd/PynTpf2pKV5xIeFTF/uRwPbZDuzyJ
MBlNWmAJLCoavODaTqwyIUAb/+/biBS+MFB9RW+XYL3Sc6CroyUwAwRNBNwED4syg8KfC1KqmDW6
W7vz6xUhiyZAY3mlEqNQii+XrAiplCP51NgsAjFcO0DJTVLTox4h0uZM2W73KCFQnr8xDj5WnT4Y
8XxIApKxhPflGlvGyXuiD+NpkELKHOmr7IW9q2xMyLJrR/5SldYHId5aECwnEmQOiLVfxc8Iso7N
WbyFNDqj66hj8wMB10PQeWKq1qA4yBqIaIiATVEFDZ+mvV01wTvO8UFftdHtfBsQ0aRsxqeo1AkW
vsg712khKrnH+hWST1igRtQPb2ISkqre9NDJEkAS+HYqkAUUanlFwIQiysqAFSU1hhelcx/xkcOY
SQj1MuV1oD1kDdY2EAXJZ6s8NEEqAnNRnVNEMn6WJ2X1l5ceGKpNpT5W2EnFNRTdMpi85hfTJ3XB
qQFZ9FO9RkVeU8wB8MC+2I/Tzr6VCqouHdOePkxA3IxJZuxLQVZNAQas7RW3eO66FLIWSUM4TTaI
o/rVS1lPv3dOXQz0TocWFrJoAmG0Btdtt1zT++NQCwxS6/NHJBYN9IKbvGXdKC6U+E2qPUDBKYyE
GAATVXhDxh0Y8HWXM+cEA9V6VBgUjIWXne/kEUSuxSYMAIr9Nx+8X4VEL7vOvWN3qlpuEtH4IBVy
v/3ydIvWdmYmdh+wwLbVyHs6zFABCflD7jFPdxru1rxcC8LoiRTuEbsvCMQ4tjjP37Ic39Cv68Xb
XtfrFMoFASckuCVFXesRjuSMpf4emk9MrMuV6MK9W/aW/s59kjumKemXqoNFl4lixi/Vy31GE5Dp
1DJWem6Bi80Jdwqve2DL6dyDm8bWl4tuA1rUzBFR/0vOnDWBMAMbzICd4bEqnV8nI6as/Ys/6wMo
MVp2SQyvNG2b04M5vUNH4p4gMwEsK+xdoIBNAYBHpIrkdbDpKhMTE4I250eD/Uy0ybMKbOlDlkan
xHNpS+SsVTRy8yIWWm0Y6zYA1+J1dOLbvvS0dFXdbOFGQGbpUrmZ/9Innb4v7b4tnWuqjssJSpGF
dZgfIyOxVIqyQgJFn/2xgmZDJMT6Oc8k+Hvm2/gLv00na55ubaYmTJPjvlSVbUN842VinHRqmiwS
k0xYoVXsW4b5iBxGVaOSWS+eneOMssFPd+hdxfcMJTrydYlTIKteHibPZQRMeC+PUgYpCvEumHh4
uM2dhmAUBt/f+BqsHuMq9QVzYbI3/+CBu9jH6E4yutFk4pSJ6Rg0K4Y0UKXfm7ivdWr9DCm8c88l
zpCzz5+3dK3DGNOegdFk07vM0HK0qHnqZCQE9iK56IGLAsj+DMclXGHuwvDS2y/mMExdYJBkVxqq
qb5SZHcyuKFGfh+O8wn76QBiZndFZob4vXPPwZIgJmhwMm3sIJ0ngttNsXkib7Ejg+I985Nf7LtU
k14RgR76LsdGTPkytNjYlK2UFjJUt5agLZjK1BbZ4jddGZ2Kvzas9wxvznx+a0i9TAjdjssSIhqV
6XJEqRcjWMv+DtlroM6sDi3JS7j9QkLtShlvT6MHA6EKolTfRsZQWh4S1ETN8WvKwFWs1Qu72dCK
hTnE3PbVrrxR0L5dMKLoey9I2pF04prxb8u7h77kAD7R8QsiE4hBVK8Rl8RVm+dmaDvcHgjRNcuw
HD6wrx3dsFAKw0rwaWSjp5FNb1sLU8uKzYlkKUYk30RhyUC9ULyUHBJ+H6Oee6VOCsbWMmlv2z5O
TR8qA5T/905knXXjApIPWjsPkWavOnhuZa/GJDZFnsmSO9zr8SYpedER3DsdMI4S0TipGJh6Pd5g
2vIPrFSeXT1rm/QhJdf/FSZTSB2fQ8/nN/U5akQSopf07B60tk5r0Dtz/j2IATNrJvo7zjo2kh91
P+IQPQZnb25wzQ9Cos/drQhdfLH/ZRy4hixB0Rqv0tAp+c4bULqy2tSD2KpvFrUEfS0zr3cCdJGx
P9MIDAXESZqXjCiCagRNikiG0Jcg6NT8LdbIupz1TchLnY3wCaYX9oygV4SELg7BGS1r25wrtI5k
kjfPypJ9S/iG2sabkLCoyaxkkxsdlApxiQJnBIOyhR83lD6sh8K2vN6kk1IXxJaQPT0I4a49GePP
Av1FBbflIBbt1AWUFMsXzY/2NtsB/VBNT3ja6/ejcELWdWj5SD8OcEgDQOLNMYjKzgEXPa4P1+CI
PnnvlURHbe7C1EMzZ7RaEQtrEPOO6BNk78YO2Ao5D0TCYRVljefejtzJkQK89loUDYigdOFTVKOq
v5BgUQAlv0hwcRAsj3XrromBNcruVZx5GQywlhzvH3Mru96gipstnqB8FU66RoVAY8nQSUadur+f
0DhclF53K0tcMWGXUbfkg4cDLDCdtQDWh7Uj18Yfs5IWG6G6NZ4OUEf3iVlL2qPj1tJ7fyUmHJAr
bQKvnYrdcl4P/camV1cFv1a/rdDWXJhWEW3Ht+Oq3TDAcWx6jergbHaUgrnf+N/QR/URbVYhxYp9
U5Ks4xriDLMLWrmbrfKNVSS0W3pjbt0JZBioem3XDbcnH/R3MEeRIFGYmgKX1dTYv5cO1LzJlLPX
R9Ri4TIynZJfbVBOwybnLJOYuNoY/4VZooJl/ci6A8S05lyRiruvyUtvraWA9Pwrr5Mzx7gfgYpn
jsV7INDbENxGdsTRBwwGsjWYxp6D/cwOIG3Ti7iWuZJKjvfAA+EBbhuiAKPlBP8aiNCucET912Sl
D6C+kZwr3wJ29Io8M21kHIPNSA8UZZhO51Z56dH2pMFy4EqnCRdsVvzfJW1aMrm8akgK468AJjfQ
wZ5X3lSRrNZkrOA3FzTBeX74SlOVtpNlSiZxzRxeQ4EmuhnYULeqzXeTU9VQps/n/TmtAL636kLD
FqC/VtKePxl7DnvWwpZ3xg20L62dpwbZH3PrRPES/brPQQi6OsHh7fQAk9wCIs4kgVAooZfLJ3l/
/igy6j0gFpvnHX22Y7l1Hvrj9ciUgz6lbCOHbJD2N+wARJL+Xt65FDxdg4BE7/Lw8/apHwrrOBzd
GFFyKPyNlnDfhT3WQClF1V1idOPfXkpeIsgsTa9YQLIiIwI4didHaY1243+S6P4LH8tFQHukQWPV
C+lO/kYf1tUjUK8Mk1tQxLYgmpH5eEI7u5vL7eROt2KLOk3Id9UlE+/vccdsulk2rRUF0puzhHSR
SGBCSg8Pdd++V4LjqMPhgD8qewL3ssd/wcLuhtJoRYbOZ67bDIz5LW1xRnwXQILFJqFedAHfEOvL
SiMsc0blhgRnK3duFuMu2TmjZbbkrYHPjOT+zb499QNEkoZGeOwov5ahEGFWqGAIQZsGiXdF8O61
yUQ75o9hEau/CLwhxUXW/bJAOu7R7/E10wsD2bN0//EC7Z9yJ4JTiI+HUO32oCCC1y5jJ+zMHdLA
AFZMuIhdqn/cRRoO70dDe8rA+lA3mogmnJn0zz68jlWjIHW75qGWM0++Ar0BB6e9ohWxwoF/1/aN
L+JC73XQbZPLc9P6F1+Bkzqe5ffixaNxHs4EuTEYIrMm5Ixf6Qqsh7t7RKutSlihKxkmfx2TxmII
6iSqW/IB+k55TLJ6syWPC77qnfaAs2CjBcOxQeyvdiV33XwOI4hDAv2E+uyeTkgsE87mQgQRXg+Q
tLmnaTfRZi8XY28Lre+lbOVFsyD+9QNzWIgv+ZMZSTLfwoNM74vcXhJT75EywVFZrqAjpWbk7T3F
b0N+iEW3yPwIUpRIurP447jUvRuAjddZ8OaVmyj+5NP6Zk2w6xIz+1esdHGZPSX+4b2UONP3E7sx
bV829DdxzoNXp2mEkj6/UwSIjVFzkXLpIjdbly+RCDC8kmtwgVmIAPLlTw+/i8F+6rVlAVajosMa
8MClFlEOIoBtc7NXGf/XbBhm7ts9OV4nArl1lgZwPiK9BFLWz1T0CJVESH7FKJ9iGSxl5QDbbuRx
Ji9bKu22Y7yo9aW/TPiPYvBONJPh6q7ee6GJviyljsR5QDbJyHjwz2/+8P0PGH0rLUYdA/sTDout
ADZXLizmd+zVYT9Ir6g2pYKXSZo/Ct+5QvozXh+uZ6LDn66FicYq8vFhzRa6mpuwICRAl8Nhe8B3
fYff7kjyi3MRjnl0OVrgPHAZ4wGnytCF+7RvFNbymuHNRL3Hc/yYrfqk9eeRNH92hUI3bR9c9LKm
fe88hX3budy6RyyqhBs+nUmcS2h8WNlO+IEJ9ohVcbzAUUxXRQftfzm54zYj9MqiPUPRUmDZeL8r
q6hV/2IwIwXay5c6Qv1iqALFbRhero76BMgZgaAhRWrNH08dOppixrwJz57j2sjBxfN+uxndKshL
YJw1GV7+QTG0wvDeaY5Gv4OuctY+fOfeCUFB/LvYyNEN1JKCMNDYKrpCXLC0NpQnAnggdoG/kn4O
1vjO/n5/1P4FamYpB/f2nbjFVa5ozPRYveXu2/4+s1GKHXpNxMn0T3Ywpsz+Lvmhj5Vfcb5f3cjg
3JsmB6vIMFExbC/riz+tTWwzyQ35cUylbMOvEDmPZK7Xt7snkkNnFKHWbRKephiv/aMchsplVdmX
dgJAbj/REpE/IzKrSitm90WKsRZP8OHbIfdHpQA9kNxbKma9y/ZNR1jfJIHahhsi81K19E5ghee4
40bI38QnRQtIrLM2+VkNhwJ3ZDMj9ppzonykBO7L/ShT6a4ddB5tD8wLfmbIdIAL4tXnqLAa00lj
sz4XXegUIkjEdgsEBAf4Ue5X5MARE6wXuDxDLx8hx45TbyPt7VV8y1xAmGMP0Z5l95bxfAjIWISQ
0HoXu1O98joL/iQr169ptTsG/pr3D65PFjLNNsQ08SEbLDvx4Cqx6045NNPtswPlKEBogdmzoQS2
oDp5JJx9hNcoxDH4tYA2+N4upeNW/1r9GOiUIPkrln3kaA1ZlDmixfT8fkL8WB2pZJk83geDD71p
IT6cLKUQg2Yjodir8cWchh69nzJcMGld8fMMxAva88pNV8sMhUmoRE8N132/s6EsTghv3tm8l6ah
xGK/HZRyV8sfoQGQJcchk4Lxck5VpFuQMmeuopmuPzTTz+7ouANB/Mh0Z1+TxC4yU6309woTeoJl
Px3XTcnTUjF/RzCFqYTnQoNVzZgWusaIwplDJy+nxlesOmO/fyN/cloPIt0UJbnFcZ5ueJWkyL27
1eX60v4iWr+prWvdLZP4WYpRxNU3kZ9jT85N5R1lY9k4nJ2i1IHz7efXdB4g6sNZ5PZh8ISdGqQ0
WjmJ8vIsQNzBGyE+CuyofqXrThMCt7LFjJBeXfrpx78Jz4WdCPGC/+Zr6C2agaLfe6niynUEWa5i
phkfWLFk8qoVw5LT9+VUHhb3RURVe7G24CMhgUuedfkiE8eHQl960bTkA/tGW8tyKSLge9Me3QcK
BWgLnZQ0NgXFhtUeV9GmMzZGTAl0zHMnaZxdbpy0DapPcx1lUVJBR0otMJMvQOiqm20qFGtk+ipy
sGR5l2Zr261cRof1bVg9MpClXvoqlcr9d5JSlVlCekC6f6Ji87FFq5jTKph1fIi0IHg9AmsMusrb
zl66V9ntvJ9PYBdZVZwUSqtVSzag7brpDOYHgqJE8AjoW3eM30wFvjfGVGkZdrx9h7cfvAhOzW5A
rLASZlAYua9rUzP16R7od7hjllU5nzl+q8gDVbtFV/+unuv0kJwocZo/Aq9jJAeEJhzdLzjZVbYd
C3/nRgibPGJIUxvs0+wKuWEeOji1wzcLNtnjw1tkfzr4DO/Pb9TNnrE11LDNj45JfcfbuwULU15c
NEClB259Mbbr5S0/rVM7cbCOTc8o1ODBfZEGpS4s5+CFiz5YXSgR/LRFEhSILVYMQSOZuftOVZYm
nQj1uZpDlYBEkAxsmR8r3iT33oZWvyHFGYVqQyiuPu4qlBUIp3kQTlNJPlSdiHTdVA9yDxCRHFCm
aZxYZ1gYqx6cz+quGECzZ7rIu0khwIv5hwd+RQDOdhc2aqC2YeBMu7eJFA8DCU8rxkxI/cC5qml7
ALb0nk4ygiEQgZ0kAs8c/SjDK8Dgi0JT+40aJf9bFBzEs4ojw/hWx4jYDLTGqekZ8DUOmsgF2ul5
yUnbFEFZpQR3KxhMzD5jqDh68w13R+ODLr5lq9je71NGuPYZ0jZpGBN+595QUVNSieV+AtDDaMEQ
LUIV6pNdjdWZ9Y2OMomg0xL4UweLWMkORXjLuRY/Bk0DdL42YCvlZJQMiJuaUhhKgMmKamzHBQzg
5a0iIpegyPz68fdaAEmjWnqsrWGfSn70iLRxTIUjzxpOsgTumPNPPF6f8K8eGtdhH5VAlkfogDvs
EaTQwrByIJRQ7++to9sANtQN4asV+TSZFzZRUcHIPBF1roiLA+NmuII8AuebK53mFBMLqPa7tu5f
1loZ02Ejjse0yhnMenu72LGVH+jOxsIoEd4tr3r1a1V0HkLPXPtrQ/KbLjPunDJGwprhcGDMyzsv
K71MwkglJIFIw2CrMQFiJJDr6d4NbTld81Huar4ob8iZXWPQwqdwyJefdZUHmDNbzC2k0SGD1yER
41GfXHD7zfIGj8GpF2jToiDW/eG8etW9WiAqRGmKGB8y2gPK4zi+ntWrZRUZ7skc6Ea4QuF/RobU
3GP1YmirXbF3LsxLkWfApysqN2zcVKype/TDvUkwDK5jFzKltA5KWRKezp0PmsJXBm+pADkvZmLO
6cs4jbnPuDR87pQgA3Y9DlpUfXVLkY3tzvWtjYZzOUQR6RY2Yh0UU/IxXyqO2XleyFy7oY3wYFoN
5iuzuOtALDYGxiVk2UH0CiVhJUHJbLp4rgipvbKXFcp4APR1QVY5GXNAKuAoGzNlzZ/lTUCScssw
q4qHkXjespLQLx9nsNEqI9kkAhFtXXpaBKa65R9uxx4IMjsbxclDNy7E3vFyiwKqeB29hUXlJ3XL
R+Cf0ydMiHJHdNGm5WJZdwgb5Rf+K0OYaz8u+7jvQ0eJC6QqplWjcHVDDh8W5jOV787aE90uGTCT
zonubqaKxZWgTMjFyqz7Xg978pHVHcReyWFwEQgPi7SvEaAV+LFqbYiHzZA5se98AldsXbeZ11tl
87rJYz4Ki5BIcI0f+3gGHnGpZ5s1Q2LLtHCzM6Nh/HD2beaJ0gRc920aGI+r+eRlubk73q0HmKhc
b38qRZCbZOVRc9wK44qrIhLMpwz3f+aG58olu4vXJbTYFrH8oLvr8wDFePtybqW4iEuqhe33sWH2
m4PmTcpPy2egDHij5Mu24REOBGVhoPe2qonV+Rkin4IHXdv0C+DKi/hBeCbmw0BeScMUamfJiMd6
mOTx4qif+kpPUh83StvlMeiLqVYgzPxZJpz1a939T2mTDRm57TRWteXvas+sFvOZBYfA4SA1U1mQ
w2Wr+W7Hlx3SYdccJmIvo0+J99JhbE2WxsGkvUGdeFrnYfDj7EZvsMlmCaPzsmf+dK1GcIy/nJTp
1Ld+iqCSCFkU/L0xSlyin8sqUn0iyyK2kPlJaPumN+L/RYYQ5mkvlrBOlNkRrikYXfBor61YkFzY
z4AzRBUXi4agLbJDFVnYQPmq2gFy5Y9yQIMWZmbjTlGYap8aUxv738LkH1XMPiMC/OqXfyvtPCCv
posulv5/G07cnhREgZPkDuGM0QdXCbsl2wXgtJMezshrTnHXFXFtG282IexFFpl5bdHcCb2Al1qL
nrbJqmwPJ4nXT4g0J1PN3NEtI+0nx4+GKVuNUwTgY1XQSUe6SrJyB4qaz4FF0IgmI/T/Y32AV9qQ
Zurv6yHGg1K9ls3FbG6XgAqBdTGyz5IO2gazVZXQvf7AcSoKw/Vp8SwJPfBgqlZ54EkGv+VndZXa
QpmfqDWMOqcU8p5CI3BVW5/bRMcr1PsQ120REvyV41LgiddWULoYBv4anYpa5JY6c/26Jkqp85Pu
ryV/uIckycQQqS8W0S7gLQ0WybXPbDUteUp1L7r0dcOimNXgQh2+XzO+BWzXqnTStiMXZb7Bj894
7l39uzgsq728BQQ8t75TKG5AB9xCtULn2r3A2QwzgSYS12d8BzQM3dHkRI7Gaed+sNXElzqrvyPG
xe5jV3OuW1VfKuI4KK1M8ocRoFzi8oZr3tImn3sG5b0LlKN5Ug3QNwSeF/2eTrT00Z+PJG2CZz7y
1N911/e1Z2ogR5qJekXMKGx3T6AoGt+SCrRHMYXhElHAcuvNmhALBTRtlceD4vO2dCyR/I0pll3v
QVxD/QF4inPVG5KJNJJxq8ZqPXzHUVbohlcz2bPpz6XUfx+zxU7tBlrvEq/Kd+L5sOBGfsrV8OMK
1TC+WKMSEi4EmJZPU/VjPmp+mHtAUWbze72nuasN4BKGoPHvYf9kqNIFqkLITxUmybJ1/SdbHk1s
3zGsLEfRB86TEII/xBNW8jIfXMGape21bcP6nifcM4qxlLEdXiGB3esy5RvjfST2pbcm8Hmkvl5I
0GP6AB39+bh4dr72kRXGuKETRfVYg5hVAaGphouGXqlLGSrGACz37yo/kguEai3eH69VBb3hSn+H
OKqfvbMAwFtN+QzFlgW+5wIMaSl4c++9JB+CxH/7E0BO/Z8TthVLuhQYOaNT5uRX/lHiV/UzPmCy
E1P0EN8rBpm+5yz62Ek+kxqQOnbfePSb6+pP31xCALyTjt0nTc0hgcpvtupnLJdvwPej7yeTOesA
9moXpt5By5e7Uqn0al5u0tzcLnkLLEkbBEefhj81YVx3aC0YSj/Xxtl68pEDejeEeIm2Pma/7bDj
fDNRYNB4U5e9FZB3aewb9QGF1NIU/8eZDdeKIqgD14tBib9hU4B9fS7CYoxHxqXvoW7BrvB8S36u
BSwhLtUpvXvhYq5FGui2vwpZ2agZX17I2QUIfpPOby5GHF8a59jTVH/HzFMWMcFxEU6lIl1TfvbU
cCY9LiM7pgZkTOheUCaA6V20GKqVXjm0jZ9U33275tWD1BNiJ8ZZNVOoWAb9ko9Dc/kHjzO3W56E
ggpUl1pDEGGN7iZCa9cGZo3UFt9DKoXq5OuEDHvj7a+yDcpWq7uhbAFSQzD0v60lYc5IpfwMymgm
n7YMyT6+4ajPhf4IyZr1awX5ZYFdosyfUS4q/+PMaVsbnu1/3dvbkm87v73GwUUHz7/fuigAmGZM
Qm2XMJDKh7Ci3MaGLrr7uWCwF5dn5BSIePjnxd31H40cDkC0bOTWmM9WA3EZ3tFBUUnN4f/I89ym
v6jb5/Ga2cI1Q9AmBZlEZwWGm4mqfJLFUcXJc+ih4c6yTuCfjByCq63tn1hO40Z23cWWRhGG1wgm
EIV9zpF9jjUC2RqNjzwf1mJOgAunAE5qxS/y0U36m2Nv6bI9lifEaW6MiUgv8Iv2F9D+BZSvZwFY
xGIy8cGnCjQ02uXPPNUMC86B02OkKMSQaHyaDmC0Au5wvgBD1CZoa3REs63cksPoXW+pnzWc0zKg
oPQttCRlOlkTLw+rFr0QrFH2oovfvlS8MMEMNcmVEHfpM9KBiWFMsSyFPqZLvIXsQjU1bVoh/9Ll
EqG8ESJ+5W6/YinL0excl6fQD33q3XjvAT8O8udcDKo9C9FcyoK2Sjd+qxL/ddaZg87kdcbkz5k7
ZacMy0u4bqM3Bz6/e/rxXbrOSH5q5rhrfKN0BF5T1os3S6YkxiXbDSjtWDVBNEssrU041qPIFKou
8sTPjG3e4bS4wk4z/RInvBE6NIr9PK5ZsLSo4y8CIqAqJsPFlysFG4J7lXTl8oZfhhmm05NlWzOn
JpOtlaET29R4NeNSLfKjWUqaf4mnuOU+TnFdzbqnNV0WMA3VHBPDvtx4AyclYWVKuHDMylw/Nnng
SJ3iP7hg4sKNJSRDtdj3uNQb76vcDmC1X3jXsfeAsfuYTMhKeVLq3tjv9byQSLtoLpHECSVKB3ig
LGF9mSpboJOKnFLtQdy75C3U1LGkUgUhytqdNW+Q9M0xXoGtjc6mOj4OfRKqiQoGYM/gpSgAqn18
i0Uh9Gp8iLp61J4NLfUTW9VpbzXDPA4B/cytb7PdW7q14BT67B4mwB5bM0/FW5DNNZisGIrzhfAv
jrBPgrb/XBYEWfVppOmVuLg9PTKXczQN65OUk9B2ChcZUa0e925MAvZocj4jqVx8pNllyMi0MYHm
+455yjcWy5tBKxmCXZHr//tDblB6oh7IRpoJnuXmuRYT+DC8NqW8mimMpRSIqb0W4TlcGJ6XIO+o
juOvTR4HxBjS+YwmTs2lKx03L4e2dMI2Od5rE1/ADbzejscds+wdvtkjAFYahsQ3wC5aM4ImRPo0
YIiX49FKzXBJYKNjBfdzj7WUOpAJvDtVXHnY5Oqpis135t4n9yY7wNIoKfREB2utgjQKjBzZ2bRP
eL/1Bv54w258VISAvna8yBw7qYuxapTQ2AAkDUToI/M1AVq8wz3NZurJEjzA0JicSdbkqCQNjFte
Q2GpguoJe0A9V2xoh5tQQGZouFoxBkT2DWOt/UGbIY8jMalabNfitjW1pqWJ7TKDCPzrlHkEEnOS
IC/NCUW97w1uCs+JMnzGMZS/Fuoxtq7T1eg06imFmU/o5hyHf80pwaWWB2xUI9nO+7+rcyHPrUo4
3j5JaR8w5j6kPAe/Px+AePURnulknyQ7OJHtFFZks/5OQOZ2PHvbLSoXDVqjfnStonHvcPrZloZU
FAgxUkCwXYsaAxpClmxrHFAfJFqBAjEZoX8pBjxr1kutyG+j6Gr9yg8K9bSfiqPpl4kaVvocxaUT
WRGeeem44rBCS9UtZBAS7ZCNtzS23NnWFKFTYIet0kmvsJUVkc0DIxHWBxVviIz7Q3qcXyqSOV3F
teGJ7y+4rGFBh79o+NbkPdqg0JQ6dz+lwRQNA3+rD79SuGtaArw9k3KzaKomO77KDb+hKes/+ik7
wJP3zidGqz7i5tNamkuxZhZjhNlASSDZpjDQceDLgmjGGx+HZAP6wQdhIC4JkpAZzCQC6UIOJLkD
FCTdEsdOUO58625HsmBYGt6eCK1X6Lb9V1SP9jcTZ7UNk/y17L/Q6UVgomsrBzC+PmOQ73DQzd0r
yYLgvDcYslBBVHLVopo+/Jgs7yeU4POlU2/PQqgwq1AbeLO/lkv2RJtGveaCtIlwMmyO3gtvNnlg
VFPnPNOL9P9ltLfkzsNB9qe1GMNTtZrV3IGY0CCNilCA7ZkJSxVio+tIXU8Jiy6LHaHxzdTbUDUl
Zw7nrZQnvYmv1T8q+0hJ66vRBUaZLfXJ6k5n/HU4wO+3OPhjGnKo1i2dK3SNXM5JLeY2Zkxt3cAA
IzU/zY4x3PlqqRSj9HtrOjMU838P1uaS+tWMXiUjfdo2CrWTxaaaYC0BMSpSNd2PYt70SZu4wbKB
+ig2zY1Jq/eLQek1RxLFwQmVRElO2nBjI1wdwTYH+McI7tlklU/coy8Vau4qRklQKEyr9xvbZuDf
RfB+2yX4yHoWCe6obqCarybL10Y2d2DJvZ7w+MEfg0uD3aR8icW84eDXLb/6utZruIByxCh10k8T
LBBwKclaH2CczAQwWU4t3ZD3hAWJbfxLi+uhUmqg1VgEIN17dlXeS/uUzC972fLYdC4yAzb+GKvj
A6jL2tuR9PxUV2HfMbnA9qTjVmxldXYzdrPsyq3gOcADQtincKmDEzIaJ/Z3qghPZ7blQfgJaiQc
7g8fX4OSVsvbJzHmW3fYAMovPLj3fJ7EpCHoo36yGfJ34Gh3aoS5r6p14Vxl38GqI7Ou99mgzZc5
gP2n2pOyTFcApeOTZeczDO2u8xBeOsn2tCPBjIhSd0hhx1gn+k4TCtf2EUT+JzXYdob5le6767v2
23+Yd5+k6sSiBLnFvouW/Wxo53ns45nY1PqLgqI/t+eI3FCzrg9pWxKZO6AGmtvDRyWXeqvFKaPx
HiSnn1OTjZVpugKmIFL6+knUO75qHygSMrlTzaRPaciukBkbc66FCZI/qYm/Il/NO3y3f32/UkdC
zu5iAy5EOtIln8YLMOpMCoTSBzTmYwu9CGwMWxTS/NSb1uM4kRAVZGBzjoMXftbKK4tF0qzwH4O3
a2GYdXevdmD0aLALNI9yvQtECDaHYHcZdin1dDK/ncyM+65vD48gThCbuy7E+YZjXrL4Zshloqe9
I13hJA1wjkXuGMcd0Fgxq0nlgtkrTiZ60Ii2ionyH6ylZn6m0v5/b0x+E6D2X5Sg4MIijnCGtZVf
IwZfwLNWhgrJOJ8GPPbTgvmc98O+Q9YFwjuUQy769KaGCJGBBtd8GZlMXERpj7772ywfQHMAl6Yt
L2zdDP4tEl0iBY27fjpHCadBYvk+hvPwLo8T1DxwkfRi5QlB7Ts6wH14EYvy0WkxWtAXXb6NLFe0
UGESrc/GJhwvlCnwdEsMqWmV/L6Cw+FnO9gKaD5XMP2CSPjd96FM43V4KP7buM1Dd9CKEb1SYyfs
c5iSQorhwo1MA4LWM3GF4iZjUQcxzkMRYRqsWg4Twu9IfeeOGuekSFlp07s1HMNsV7FexKmmZJtJ
m3yhI4dqi9l4fRsPjVR4UWbEnFbCaLWwk1TNVa2KXBMXC4Hdo6xos8IfH4FIVrGuE772RdktV40r
JPcrfkVxqgavKH61ob8lWtcr8UyecCnjuBmrxdExxuAwIAIme2pzKWBGYXZK0wjjbgxbw921EaBT
NvGIdV9MXc9NfnPk9eEbTjC1QEhzQ8R/ebQLZpSS6b2znxNyZNCw9LIW9Bq8kGXztCEueRKrJgan
wgRqjqU6UN45n4Vq09AN4N5N6zJaPSrNgBGrYD/9k2TAsnfstOiP/jwamw+DO1NF4nbzT+83UZgH
QPbu4qFcvZKeVUiPqjOUtDCONEZfExbQtHQfZUt8cGW4W9E8+Bdg4UzHnPHD1LUievPjpWSFg1cV
b3q/U/r4g2D73FCGMnqoRWskaUaS3HCOpIHQx4B1g4SN9jJx9sVLlxp4LBI6eoZGgXYc0m+8n84X
X3LEatck9m8Fj54rN2r67FS9+dUFLlgiZp0CZ95JQ9h3LFlsR5JO6TpESqTAGWNWsh+JP8lDCQAz
YGYGeKisCPz5DpN/t1rv/nvjc/UbpDqr1hiSXQuEQ1+vQguyuqqpYy6q8e0h7YpCg51Uuhfr7jBD
BHpe2XLqakPw4rZWuzKmzUvJfS+klbtMPK0V1HD6UIPUZbR78INDL6NCG6WZ34IoqQ3JNS6Z31Vt
UVx7XsTlO1C1Spr7fTLv32bCWKUYYuQbApdvBkHUlTXEFq/KWy+YB+Bca2uqWJsTaKAN+oga8X0x
vDX1hd+7pyo8CSvfvoq8itlnuaImbh9PVLFJdH4Ayr2lGrqOZmRV4+TfhmDtblHqZzx07qeup4no
dZIEnvZ0VpSLPc3LpMp4Fxcv+prsOjmJPVW9wjTYom39lTNzCz7FERuunHocNLnCSZh7rfyh8RsL
8mXNPsTc5lunuqeqKXAH/e3wDUqIzrTLZ0D8hhn8xc8x7jQ6yI4qCk9R+9ZUoRScewADKA1p2Qrv
QM9+rNYkci1IUlBkEoe+aFzv94KOOyDa/TWDmN/65bunnWiIIb0g57VgIfE5vFzkhxyzXA++Cj14
sSbluQI0bG6//b537kg1fwXKEf4yIOKOPqsgyYgtwNmCwdT+VNCAeDVjtCck4SuneA4b16/DNIDl
kcmLmLY/j1zS6oWx2dx++vyZUXWNuRP2N5bXSMwdTdQgFpyqMzkJ19pxwtC4k3elyCaay4ZYO6sN
yau+9mNgqquh6rfPFrszmkkMMZwGLUIS1WxZo28P+qCXrubLxF6W+5s/mHL/6YgLoyqTsRowfDcB
LpOOpq+s6/aMXIP/h+CaGqK3uHGY1erWk8PBL71AQx56kYPQZi+GhD3DWeJLPCnHX2SQtOyPrMun
XIcuvdvQ1yzqNo9XrO74qKAI3fec51eSY/LYRxoTssA67EVYpp6jc5e7YgM+t/j3S6asS71FfVzO
crxBCAHSIgmccgkGzHYLT34Xq2WYphbWsdpCsFKj7ViY6mXrvG2JFqu/HkkNxBys74gOhU2LTt8h
OW2+ozevzewevztjBoyqFl9EhTKwA7ACFBUkUDnHMyrZ/fWUllMNuHmVw3YGBt7cV9BwdndfivPH
SvHQvZXAbPb3Yuh655r/82gS9Lz6ALRcF63otbByc7XXt+jTYwxXDHQv3ETps1GzJT9dKSe3Vim7
ASei1gLL310pJaPi2CEuWt/V0Ks9wCQ8WMRoPwIcq2d3nyMDrKJ2XpIGMdXbAG2/6pEv/z/t+9zV
2X4H37ChhY81NyH3/sVsYoh0RqAIC7i3Yn/dBF0wQetWXhqKwhMD4LVJxaGVToqGUMXwcOIemLg+
WUolcy/7Za2Jfl0RdrZk+X2dQ0FqYJrGxOUAVVGnQvlvwmGPGKBZtwL3a2TBCF6yTBCotSNtBuCc
iSUq6riRXD22kx/jQyCsXrzgkFGzV/0TOX+xRo/8OF0OcMomuUVyO26m6+nVwFZjcotT3R01iy5V
2KvEE+PqRJdTzyNEUyGnJ+JJQK0IbjAwEOEga28FwAGQeV1KNv24B+tMYtb4RARamxXbPxP9ZyMo
byG/0pTDl1L3fC0THlF943mtv9otkPCQCC88rgKkVCIKwueV2betvZAWvUANX8eTIcB3c9PkKm58
pACjLlQUqRghkkjI/wZ5J/6LquXR62lTfz07B7AcbV607e4vAjPqixwJ4UCFeOJemcHNWDrpCicF
i/+rjU/+1I1dhlXNI10U34yLEpc+1KY5i4HiHYKkiARSGPYXMVAeEUwk1iXTqP9yJLH23lmeWaeo
qLboF5KUF3rzOW0tpTi2msb3dJQ/Yqb5uDAFgkgimWhUUQkxC0/Xa1DoV3QmcyDtG4aLzB4d+Tod
boc2rorMeTynuYb7gN1OM12YoYIUz4ug50wo8JaI15etKiUyXywX6u8F8NAxnumKC3OTd7KUtItK
bMNN6to+ZE43AqZvyZ5JJg9EH69Tl+5n15XRc8ClE588CKGGaIJsHqGLFsZDlfvrLsXELFB6USVB
4+GoF4PozQ5/Iu6j1/gQHBTD/3r8LDYkpVt4pi/9RN9yBxwQgwGrFUaeEyqF+O/2bZAusTwEVMxS
ybJX4zSZC8YG6nqhdt+ue1YAWnL2ONJHUA4yGR/nHFjiDVevCOI0VohkYU/naUOuoMqKtdK8tDJd
2F0dZM9vbI6iLCq7jUOI2FxPkvHRkPlvitRXyvvv8mEjFCl8DnGK7X5SH/CgTZyTPXAAShnq31n9
7CiGzGnAB6Wi1QQ/P/Cbc1dzv5RPHJEYnJeo+pqJ8VdO3gg7Ya/vvMkD7JTu4ejuxm76d1FF9KEx
l978/HdkA+nwWUps7O0eIC+4TF8D/FTNOU5C6sRG6mWTFvexIWWjNl/ZtW6Y667XEPq6CE3qxqbu
dWmjARt1iW/s60T9m/z0vy6feANznjZYRTYCfS4XqSj4Dm6kiglu5zbdmul6Hmswm2ihxHMOkfau
4IpFXV6LoK1WxONcHDLTZWPFNJhk0UB6yq0jZVciBouurww38NcrHBrvo0dwci6/89b/IDLYpY3E
OpoGimuS5MHiRtojyIZfpOU3V+8B2v5wPeDtHt0IVAAvz0VCVVEhXn21opkIAOGJfrH/DS9LpV3n
Goe0Xd80X2MN0nbdj4II4z2Qe4xcbCMddOtRaQYcdkD32jdpynNDievbISSnnGrT4Vx82nazQWvA
GaKhdDPXmGnez1lGbft7PCQBa0BzXjygiXt0QmVQ1agNeeNZq8O72dOCCu+tj4LQ5pfrKRTMw0TB
GWGXB3gLLPX78lSU1myfxXPkY4TN3FgvLqPVdn02vqrknRMviZ/YHiAi5AXzQUplqP3vxTRNnVuv
TPzvLnNodIiRunHiYkLGINIJgozaXw5FyavInuTKmd81sbXNT0qdZSrKtY0njx9bxsite1m5qNiI
0GaGoLTtL4uAU+tXGUmSYGAXiQuklkLchSoXCACLlzhTsXu+t3vjVZ3BWyriMRZLgV80euBC7AHV
ZjA34ZIqz1nm2DBNkcj3rRACRO7wuL3CfmZicVLqPLFqlTVc9rccwGXGVVAOAIRy2qiSMXuIzI0q
Z0M86YtSJcqYB0eedYIQ/bqcCBVZu6hpMFjqqTXf579z9nwmwWhdBA+d9MHdc9th3H1ropcaanFL
iawRjh3vuPuyPW7i/bztW1tC+SfOs8FWNR1CE1geqkWdHsC2Ro9Fb9GfhjKkTYahj1qqlI5I1C7f
YLivNFAtNwYBHtiyL+yNvKAUWkCQl5/WI/+lEecVkDG5E8fO1/1rYPVNYdwjwIzHHnA+WqQDcdvE
DFkfN2rOidxsKByhqp/vAbAoxrXjwVFOC/WXW+P2nAiILMHedVM1FiDMA0iKa00otPYPQyk5T3mm
ZkA1F8oTKQ2DPnJpY+7omdE3SWxhZBs1EM8zLGqEOd9ucJ1WNLYOKpUrpOicyxmLy+Ul+ZOaCcKj
QCoK8L25fjENaCnxB9RFzYNH5AZawsunm1JLlRTSGOTScyRaLXYe4U2Mz4/ytMEng/QkvfZrIylV
HkxRlAmZjz4T7REgB6c/kaclFWKjhAb259S0EMcWTuNE4tnzZQvSlcpFOn2XST4ma9NjWq0e96M0
JtpW0NBUyJmqZ3EB8KQtS/53AQkgnfTFNzqh/iNLyrnXsZxHQCw5fdkbaH02VE8AgcIHQwHLazL3
z3i32vfa1BeGH8XETFTYNhTnwhOSAtxA9ypBr5iHzBSom0YTr7XaAJR5JdbnYyzd6Nk1wdi0xdfe
AkGX17AKuszyralGsghWiH9cPrkJ0ypphGjYXPn++QyRs+SsmAAuEL3Uee9bZlmzEGOkSy6H3fuO
9FovgbREBg3eUmgGdzjBTUk8sMa8OPw6H79703netouVicnHawmNYAGM6C0DmRd/foj6h7R6J1p0
+1l3Sx9fQbIyPXfrfygr2fo1VJPCNfXcoaPJbGOrhD1WUnw/cjGCrE/krWOlW0vi8X+chcClepmL
6rqfA+gz1xowTM78Y21i4gUQLNXTCtsbbIxArjTeVG1e8zo5I9RDVrAsxGlMMtImm03Hg1Sx+7xP
qvQEMLyMq6zfnlALaUK4OT5mE5VhVzaAo9QTbi7+uiDP3OzToqx9C1mFojeSaPYzelL1+WV94lmF
rYEawegmCkYWbz7/v6lgRh2eLzxBMZ/J1QKTtWW9s5GXCJFIVy2EPdWSSmyHvGy7cW+uNGjnqm6d
TPbSGDuc/qyoYeefGd7eq9PCKvVRi4eWydSWYtNWF2ZNW883HcPwu2Ks+gjPa6IMFXHJUmdIeZ/l
LXymQz38ll3rk/PqUIShpJZap/d/2F+K6AMVTscISxr7BGxY0N4EENGMcmCROzG92iqNJF1Nhd3U
6g6Yl44Ov2nVLKPXVovsgPkymFkcKyYsJajL0rLnenjOXX5Tl8Nv0Jfq6aG3NB+S5loNzl7zkjkR
9Gr3LVN+3BMxUfmODiRXkV2Tcy5k40AS4mu+pVtjlx1uKF+DU8D1KxJtzDXybmdex9F4rfZJoeg7
OVI1SHJayU/bmrAvB9yHCQ5t/9nIOeikeW87WgZUT6iIOWpMXZjNoa+yNeBtG244eQuVaEIYJ96y
kBmCPbWmYDTB4thoVzHstLAzjTYLFocKz4TEyBgmVz0OPbBhtSPANzX1PPxCJyZ7mqx2ASZbD3C/
DGRIr9TmuCycULDi+4rx+Q/HbL6DUD93QEdhJeIYF1oMa94wB/WiOMyLPu+NOB+SGBnDEHJQC+zs
/71KmzY50EgFr5O67w0j3ogD6ote2bwY4DsbeHTg9DU25HzfD9TcpRK5IuZ8D/4oc8QQHtoO40t4
XHnx6BURavDOE640QSo+tHAQ47AdK6NZky3A5jQ+TlCu6LiiTX5ng3nxmjf7C9tJzWF7zgCd+3BV
mxjuHBNYYNvGE/hdrKYPpbV/b/ltlWvmZItxIDBmAdLlCpIFBFZwsJcu/84LQTodxSWQLiIMIxGb
9SvlX+o+Rr66CoklxC0VtugAqSPe+p4FPBo9EUTR3rieAnb+OPiW+TNh2kF+HnbrkSSYe/P7Esaj
qSsIpsNJT1AKi/Ur9K2Hxli2jwLl6/KE8yq2qd1CkbfBKHOSToiuc/FNuxyBd08lpUec3F83dBJJ
FJAYPcd4MQFrQsv2zcTY6G7/WQEoINM/wRfkf+0e1awOR16i7Sh5o2gKulV0tFdeovT5f9uN1ysc
/8PLWQoMFH6XkAkduHklj5A6hJPlPDQPAqOWuyRiXMH9BjdGzS8yhDYrJ3nMXYzUUnkiaKrLwIh6
SE1JyqwwhzJpQYEyCC9QJ0ApGJ8hLn7EiLaToUyPH3W4Hp78yHmgSrxBsOpA76qZI6XA9PcuvLHu
r8l6cW68p1+bHvG2q2yMEBfnYUZwV9mevTLW01EOFkCLX9NNkZ2e0QHKxcPzhhXBWdEbHRpOO2rI
XzcYK66OU+D43w8Hj37gQG+kHpTnInAd7eb0jr/TjcJSfOlqkYO45FmaiHFuRb5X6POSRBS5nTes
qea4Bsn9U0JyaBKzmraaIBdEAXxeAGtjTuZz4tgHUnfiUSh4a0EENfjkkfZaqF4N6OkYK9ZsQTP7
VCM22rTH54L4MA+VAiMMjBATsAplsWiySFakuuBCdpPEabyefD7OS9Zx9ibn2DEmn2oBhN7p/Eh+
+vecfAzxuug+ADzw7gJd9UDQSd7x5oDo1E/zVgSrcdff5OJHzSrML0+x4m2vVb1s1th4j4duK87N
EoNHywywmFTa1vxvPg4VKTJqsqRYZYnadRdUE/PY0MtJO8LElTdbNE8SDNoqebA6snJ5NAatWhdI
fhdJFJYLnyuPyOCcXE7iDK/V25IviinpzCLOripfSW/OHv+Ot3pKJoqDioWzbZfwnMX+OPAtpka3
7nBBHAqXLN2hdkFMkcNIxQBgmLAuYA8U9wN01O/uLJ8RVmFVIjh1LiGKftRiu59y9lvqNnWEOnD5
nncOCXlIpIPYArsx2I8iqcqvb1HTiV+ctv0nKuZSkxrfevPlzwzDe6h8zaeGi5tDHxj1fpSIJgfZ
sy/zw+Kut/BZnoI6al/dXxMomPKwdh1di07sv3e02kRXM7kYNlTxJCaviaD6tw5ibyG+6sOXPbUy
di8sKcnCs8sQuI7M+NLQ+MJ3Cfj5o56eLPTOo1ROC0aO4k/dje41kgP+QD4jONdF9PEn19at8NwQ
ABwxs9uj0b2SxSQis4/+Tne8XY0GKy0adWAWVqiCr7ie19cwOS8wxptwWW9PCquPOtNDhkp2hegZ
N66ZgAOPjK7Zl2Sc+t1NyQLJhEo/fgaU0E5RA0MjK4jaWfinBEQwfg9KMZmmevnGD4ayBdyCnjTl
TEz+Ar8Ruo4/GtYssXjfyPhyNJrI50t4qRuNpbjdNky+S1PEWvgGKrw49wcY9KZE106bBIZkmK4b
tNb8ytpzfpJ3Edp6eTQ3SSqMz7BpPXEK4PDcy01Y/Z2jij1Hg1C+vYFFmNJEgo52jz01o873oO/G
20UybcA+1hDOw6sn/i+A9/wrV1/l+XA0QJLAAxInlPE1kjw1PwUIxKBKFbz9lN0qH+sw7CaTQSQ+
iJT/569mcmn86QlUGTFUmlFIudDkqE1sSTZ7/Zpt+3jPcRxTSrYg0pKPR0iS1AQs/WO8C5yduMu7
ZkTs9B7cPXkEqQgCKY4T+muF1ai2VYywegDd0x+xdGDg65iWxsnHQdFpoMcH31En/2YHbqiPq8//
MwzQ26Y809F+DUD+D11/viMyzi577o97m7W6/JMLvKXVUQb8vN40FvbwHuTWoojH8xGSJQMTzFS1
h7TC4GDl3hzWm+jkmh9aVSXDr1uSM9I7fYR0H8553iKXOkkbe3uq/PTC2ZLnxk1eCD/pm6j1xQul
CoAiBCU6gEWyVJLtTWmwedYwDCpQkDrTTFLSTW5rqh10z6wnoxbwPFlX+IhxVoCyJSxyaHshRrlw
2pb2eeYkC1VaS+mPk/udogBy/Bq2uWuEirHDG7HvXXxBoW6eu/KIWsc/shAIOO7EgLHaLmV/OGU0
yZMwPQ628dg56I639/A5V7mroHgsNSHR42f/VXVqgAH8dz6IQLgjMQl/y+MZdWGc097C3336mmZd
PZH7jecchCOkckEC8v8vfxhYEWufUZ+3vcZW5w2kMl2u8GyyO42TUmX+NNuqGGe94v09D7L5t2s0
yqIZfqjehZOljSJNi2njmbYTw/h8HL58YzRnIVCIqLFrCe9Heb5z2QuMpb2s6j6UNxDL3cnCCCnv
2FE+f19WBk4JGOX4ZHcyt7JA2Tb5XDqKZ8Oi+Cbu3buwkFTCyYLQhb8pEfoUv65hwLcYHDsmHkAc
bgaUP9GvyI3Lo+rAfI0bCcUK8/S7JXXdTcQ579A4RgFPMwrYWcOU5wSJSm9QSHytNDm7teYpFfbJ
RY/PBHWXOGuiTR5D50m5ImAWWOMSFRxMqFYIWJ8KxgzvqS9EIkPmPR/kCOSXbOcDaV7RNTVjhT75
pEkcK6NK4yv7oarG9ySZ0ZioqpNB2BanUA5OHkoMTjvAX5uhT9tQdAtWkuuL1gxzSVWJNHO2C/6K
qzyPLKnx1YbYLNG0JjVepc4yjRKIa5fHtnBLvYHPag2Dc2s8FdLCMRrhbuyMR7+ysKrg1YSQcsKy
Nff+aU+UPhkO97Eg6lOXu8VIJacyTi/pldrEEkxyNf/Xkq7CkJ3xO4nvc2uIEykg11Laek9vydx7
pGPif5jYBnbnouEwmXesIqdPmri6m+dUEBfpaXZynLlGoYgB4Vx6v8lBVq6mBV6ww+CegeWDPMsH
qlIxekkU+fOXnvD8JugUv2nqPsfde4yvPYKKSpncJgb0hxCzt1NIYPJcmHBmgXWld59bDVcCwyQB
vqh7kXh0i8EPH4S71S8FadsnR8Wx8zePnMeuwfGLv9iw0fgYe2PBZ4n7UUYk8kE8xaJkoKQRLz58
9/ADioVzmqOkgCF1rilWdRkzr26pnUNl+E5NHoU01mhG4kJH9rPGdU4fy39RTnE+5ZxsdoaURBJT
+uRT8oqChuOJp2yBcilhba0Co/1nXR3em2STHL6u1pLQElFyfQFkaPcx61/wc9MrDms5/1mlps99
/SZ1056Gi3pw5WNjAErtgmZQEI9czVrSJ2LferuRLwM9JyneSA/3iGKrHVNMwFTfga2ZFzfx3VIN
UHk2avZJ1SqzxQbpgLKXNFKyFphNS2pmByS6LK610Z6jUfPs2sojskLdgFMxcZsQ7iWCsGTMHEja
noz/Va1q3to/jmlu84rTS4MCy/hVKOE8S2vCv0TYLPX7HXMBOwjCXramQ6c6ej6dIhPLN1c95ueE
If2Y4dZhVoXouyu2oHu1hnGZkt0IdrVd7n40kfE7GCvoMRyupBjwBbgZgi6jwbNwyHAYeht5O3Nh
KzlHdDPOv/J4Ksf3jHvNJHaJF/mbg+IXrBvxjmaBQRIS44MqoVA3vCTe0bTaEUDyVUDFySxA020m
xGTYocPXIVph9GYJ0fN8oVt9mGKegK54jILoC/Zh7Abtnc+stF3/41im4td0uPcompX/MbSmB02G
65dqLMKX7PLhNVphzeRq8fI/mTUR/vwFIlTn5lmd0YywX2oEisabEb2EFLfqnAxj0KRQ4ptA5SeW
EYKAS8opVEmKo7ATXURAOVHTm7C2n2wfWwNFMdamqfBpun8XAn6DRq+ryMckVrKgGK8l5D1WaV9D
cB/Xrmq6xMVbSjB/ySZ1KuGFvE4nq8v4cvLdfgMuvUK2WFew2RqPNEVt6Tiv7z6mT2vjkPS+zXhw
cUYElYsdheGl88OPb5nzXnCsiXcc6h3FhyYQaHUieorwewfkYv5JRNHMj9Gw1nE6HT2MsF5zWeI0
z3UpOMJ8M0jJ6882YAiUNQuuH8x4+CmvdGg+XvyLlMvhE+kxCFlWH+lmRdGYyxpaXhCtOJKq7dfa
K37w4s7JfdE64bc+r+NxCGcCCVE9h4idFJzdsurNgMXydLsOm37RAYCuJOacVmvIX351oaSSwweo
KqjjDh4la99Q8YUp2ObCOzfUyyaF50KGlMOaT1+KBxdu7V1z9cFQ0tKbK+Thz+Y6rimzlEDGnKgt
zxN0xQ1hO8HoI+Oyaiiz9Wpvj6ko46u344OD4FqTK4jXZnfTgpOYIUW9Wzzir6c0AwreB3RK5Z2m
boMfLBru9ofCheqR5BmMhYP3MtY7UzB1j6yj529c6jhPIpZHqSJDcwL8DGYBmLMXcE7YrmS5NrqG
W3OTk+Bp1c4xLyyz/bWLXKVrmxJ9vJlJuIlKrv+da5DPTFCVuokeao7XexknDOMbDASNbi7yMOlD
yaSoNcXH+O7AxvyYtyiuQEnguLuxykHt1BdlQPKQq98D4AI8LOOtUG2vteveEz/vFhOuNtGNKssj
FZluHzpKzFPAdjYmJBEaB1BcNiIM7wkgGAurVfmLFYKg2F5TgYsRKHWaYR6jLIdH9tWN4cAFBMfe
2MlCQPKGpJ/tuY723FD6hVtZIdLxu5EOTVqWOhFTAI8ci75qfXaZkJRzuHA4jgjPtOad6UKUsFLM
CvfgI7jWHN12cTJdLkjB4Pia8OhuzyWmzDbRkVBPJbPxNU465AKv213q6tirw0rd5rPEXt9iVAEy
ONKaD71hudST1biBQeyTwuv7UjaDGp46vceD0bz97AuYV95udZoaSGigcBy994UBk40iHUpQY+ZR
r3k4ovNkCCgAxA91MOBADNa8bo/Jyuzz8a8IlbmWnJ5XhTwGMaO8uNBvqAYUSiOjGsvf97UhFthC
Wbe9SzSW8S/Xvzx0FzWGz2ARE8elWqEwkdH4idy30xZLDZ9ShvkDRaAOtSu63tpQqsEnyuVlUtxG
W5TzQ8EInXCfls/IlGVlko9UCdbOrSZD6o9+3yGwlGjT6Jm6M2IB4Ew0aPcol4/dxtp6sFzNTqRQ
4DFL/x0RMDa+RjCFQR4302kBDTnKqHMA4JmiEEFnGx0NK3GJn8VAJuket6IrNZAn+jzDPFgitAXL
A3KCBh3T17fwi6uh7pOAbYvt6pA5Dq/5ZYkL2G8myqGi4SQlO85LA1evZk1fvgX0BDNJQJyXXhhZ
5l5XEc0BTucoe2qMrfH3/8bgq1IF7P0e54YnEJ8TfGcx3NrfZHJi6ON8br+nvzhj4HG2vwLg7uPM
/1asf7Yq4FlRnl7I0AsL7mP9l1mDMDO3nfOYf3oNHMC+FE1XItSQazioTlNKH86R3l6WyKKqtR0b
190HiawEslrfHmKxy9uGBvmyUGgd1XGfj6HAAYsh1Abl11AESc8jhbm5lMxJt8mIdf5A3M3ZXa4C
NYrUm/sEmcX6JggcbF8zSK5fGGoYGmMWbjLj59ZdoH3wlrBJk5i8iJO5pv6HL9DLhQou/eahdlzK
Pinmcd8Xwqf80kNn82WPAghw0VN8uxrT78qbhZd+Sm+1a9Az5lQ0armSQ/OHgto2zJ7k3ZeoX7yr
rIZrptE9VsdxF7kTlxnpj6BcCaPW3ZlDFwiBMEDG9RvPSq16UklMxoUW8v6Rsjq51OTe5/G+NJ05
7yKdvhWgFsjO6H5DQ6kZZAO7hS6WcENRG9eRE98Q4aCz7e8VnQP457EZpErtE99LAIPYX9A+GUgA
4vnAyT0MqAzU1btA6fNM401umQC9qV/OVuqZQky63f+wy2t5BJw33GcMY8ek0JvQ9lISSh78XZAa
zLADZGpOCxj8sI+Y1t2yVUDQJSZtJhL0+Amq5a1XKSxgaxC/nHFJdJ4O0448E1NZhPkIcFEoOXh/
s0sk9ilefO/Ek0/FEvirT6xXABkbnDjPsN1gWhiR7MHAoMG+pWR8dvtjTCmuEaECKkITh5EahQii
2lv3AlP8lXT+P4Y4c8SNpnoy8FhzDGnyPWdxC4f5GhrLaACGEIz2307ecT9sGRiEvEdfLc473FN8
jhyYoVftcuEubWSRc181zdsAolM4yY7QbS7Y2iSEoB0fO8bAZzzk02HN96u2fSgtTtX3zhdAMl9u
O8a3sxQH/8BPGEsdKNQYvQihO/gojJqSj0pyrcxYJYdNBlNq7Fc6t9HRxlFdornyrBxeaNRM4kZK
u8yrVrAIsKMqVqR0+WGH4YJMDNuaACMnc5q/MBpGW/VAbLmoIuzUg1wAXMkXIg+Gg1qGhg1jSo8s
6p9VyiCQSP8WD1pUBq1r4+YnNmpEG3D2ZAj1ZoRHReG4GS3+EGH2S6ijCc+s3gTP9MVMp9H7xuzv
Dwzami9PjIjwOyL3H+/4w6qcB3YZXeSa0/96z+QCe2B3JDNelKe0YYD3+Ok4YgXh9YmSqzste2X5
YGzjR7I6wcOccDfBakq8uqDOjbU503o0px0pCxcKBvuFEmrcWTexLQzyerly+GXIk2slr/pzlo98
oDob9GvIItKF8y33JYoIRXPisclsCAJdPuA4RKizdIxIOFmFoL/M77MV5VTGjS3GQ6O3XmtECxfM
wSe51QrFILkeMLzN8jFRiVWEGhwVoMLXx86amxADRZk4g4x0uEk4mpCR8Mr1Uhh5beeN3pteb+4q
T1is7oqN/DOF0Ue9S6rndjWcmXqZ6h4W5AW0NBjw04Zolgs54QjImqPhGvbqlYK2ydvPoa9copM4
Ub2Jxjf3QEd10LeXUtv9Oe5NkKFqc3qW6Ze6pD0iH/U10kGUZ6YvOBoC59DHwpSQ6kBC/gj+3/cw
zgVRUguyLbf3vvikznwel5TfwskjmEIHvBBolqIeCbIs8wlaCzuucf/TlB4/FXI1Zlggtf+jl+M1
endejLgUR0AiO+iFZ722NlpqhPuwwcyNiIxIxtEjDwJ+bT+WByPTaNUDT+eqJMDpKgaEmjZOi9M4
9G5zcbeamvO7C2dN58Tcm1J4kW4kN5mL6WlkYHjnOH8zPep4KQNdeeK0VKEhAPPVnsYob1cBc/bR
ygbmJ19YsFaL3dIVCUVm1TXyzKlgsm6QdBJh9EUPhvjl88vqGDpBUU+6On6okioa9e0SR3hO9fuV
1j0gl49TOsvxCSnJjYMh+wEv0wUZP2LVae8kS7BISMAHdIw1RtFdsdK5wWxalCv0vdB2f2/S1YBt
/Hh/nBG98rReDi3TSXWoyXW1kY2hfKzZjq6yfpxSRvoUSozGf56RZZABO7fBmUjJmbCodWcCE77f
Ge0mJmWOq+OlX1mT0rhZRusBLn1bpLdztduXjkqdkFTN8NpjF1Lcuccme6kAtWBtdYMqgz/EOoNT
IFJbBUjyip3aTbeKuR0l2rVirG5X++sYE5zi4F6V19NiHE5kQLwavGRUpIn2VoerodKv7QeXepM7
bjTnxOmaYZkfv9pxGaEu9/fm9OAR7LUL/xR0BBkRfa+rbU8fXY5AqVcDPv3qI40FHSKz7uY/OiQe
Z5TjrL+o2kcR85kzorDDcqfd6lRYOWX6WYlopnrYlCC/KeHtdI9eV0CR3RxwCH67m+Djy+FuD90L
zodTPUJ/0nTjN/sRG2GrqAq91Szx/v1icINJo4kQ3ki1guSS5ijg+4WsMgDo82BnreP9+WFAefI7
ERRLFkfAYdIVgD8jsp7Dvd/3xYj518tLcE5swEjLWeFYk0OEmSHG1fK0tZidjRj/qr11DtSuneJ6
oKfS8kzvYUqCacl7kYIruMorZw5aUGtWEpslSxC0egfVUrBKl9qqX46ns/8fF8BJK/qOf/2Zmljc
1D1z0Eo+oSwb06mC38BoOw++QS32kLWDj8U74DyDCccNu+D9Z2kV0DgywTNM4B2rQ6pkdW44LDQG
cVLwVs1K4xnZ+UYjFzMc1wLHYrdC75MGf1UyFvW/u89NGF0q4Dt7IvPmT0ELESzgWwM1byk3tzmp
NbiM53aueIiVf8GQs7sQPuPiO3Wne/jzWWyMBgk5cp/C/3tALHOt4yY554QrtIpL49P+zcx+yiMc
DvIpUcAtYqLJyBAaRAx9WK1vyP/pxOXlKKOAzCjuMnSKd4gxOWGS1fL8lpLaVtFT6xP0NoDvXMcr
0y8xloPhxceVpQA1qRZw5hNrDvHvqaVhnzU1vkkyP7az2Y8W0iVkuFdNtlYJpddttVCP4ZEmO867
PHXoQ0+thhrtihJwHnEgKF2su7g2RvmfjVU8Qk5C6T0+y5RsNk1pt8qf0wvRjNDsNZBlcENKPU/u
YcNlwfzTRsMYq/RhiD46r0vglZ2JfskNlsbRXP6+sD0sDlLuVrR1wDm3B6mvhFYg8O/KciYkO89q
j0ZwsnL7B9ZWJQIDwfN8cvNxTFD+lMWtibKImCfesKZXynnAS/89H+jdPRnCodkFLK9podvg6bUp
VK7xgA+uwh8ukTNU08KjD31aqLMrYFK9X5Xg3OnQJI4qsq+5AnIF2V3akwtQWdUY2twepZOaS98Q
z+FJ7cYbYOjgoNsj3P/Slq0cyuLsF36q1CLHXqGk4uSNLXmsirv923xNWYu1qCj012L0Eoeoejys
puYG5IOBzYdBi6KTXfvnyyynRU/jXgvO/TlNooEgN7yXdBb5xi0lxPX4cZPIvz0FpQNldvwNGwwG
sfqQgCcjDlQrjNnA+t23xsvzZ9WzaN9qEinhOyWPdveO1wKPYvKJ+Kwyo0/4zBo1XS7SpBwk7oNv
0QD3Ix6wI88PQoiXG3ZmnrrwdPvuGjpVMm/SMqDABxzFW6+eRoY+pL9LPQjThg8fCdAASsRaXu+N
XeZGUZ9GtAUTaMDINcsm92R8VLsxu/aTSHdEmBpIGWfvQTs5lQN4fVndshfSpXX4iuzjkhggPJoZ
8DwGnjx1P75wYqXlWYEI3JtlKex5jltnuD0HhSCIMH3y8YyekbRdyrfUSh7fVLXINN2f9cGfkunQ
mlTE5DUYbW7bAJ3iRyhKh8YAZ/s69oFZmKls3PuQKD7FXrBOEx4LfI1Z3VtZ2LCyPybYIZmDaI8Z
Sv6M/Sq6vjUB4vWCiKmkumCl5tKzHLy0mnKuBfekWlZtesexweoIQm/f5Y977vtA9SgwKtJWMiyJ
aeqE9LK5L9ROOKX5tAYGxV7k5nS0xNu7hyFYu3Uy41/ZFFspgNiEle36R7w2QIkFWFiM+/4MShpD
tZRljbFF1Vvm9eovRVwS7qFdjnEX+e7WcarJzlAq15qqeUXnuxix96W5Do2FZJbrBa48f+7GJm2+
Ii32J2itG8JTL0MV45LUa5r1xeK0G2dthG1XXmPJXaE+AXZWVB3Y5lJqtDjmiTqB9w9HwVyXy+h4
0Cxi9q2LcPKq3dOUkeZYYukTVPBtyUcoerhEHoGoaFkRVyr+K8dQY8BnOa85uW5x/FmhN67xo/G0
ynk46s6m7AMmTEsJCn0r/IPjRz3sN/zwptHF2O7VjKgippkk1PmEsr2sVg0ypUsdvMss7jB6oB4l
tz/Hn0FWvI1tqgn1Yr6Az4YOENTcDHfZnDQ1jkrLFDhqkQfteSQwA7ye4AbyIQNccu+5ovl3bWmM
qOp7vtgTxj9/n1Dme+XurOJWj8sqlg3jXz7LkN4W4LzLYR5gRgmq7tl+1SebWLpmgPfj1yAdv1zA
iMHxrM6vkuG7B65I9S3EcGjb+PlEFPpofymYPNi4nraBYBoO3NGwU44N6km1fcT9BiY0AItumP1x
8uWZCmozeQOVQaV+lmNnrBmWeg68BULTIxeJP22gxwdbZ9ko0flwqAnfis9ckorH9St0WBv6sK4o
97xdlqaKWwl0tN9Sv/lo+PUkA8jjezWC8wpCxBvYn5iHW6VTGJqhXPRqZc8iMhjAYTTVVulD5FoA
CB8Yim5Do6MaepnDQtbZpHy4J6+uWiQz3gLxfzFyr+Z8SfHabBMYdyBBTmflqlR9pKV06ODR9eom
90c3HUBvujtbAUFUEvQlZvOirlVdvlMDu1cq9w4IeIUJf8ETNfYRYPP/jsoMg/uAPTGaoxvIjyET
ynEqSCETwiQm5gnVig6TGvyN/BEKSnXdqFwloxJ4DAtzi0uICIxkXQJRsWQuXW6TNkxnYapov/XR
4dGVU68IHyaEwzFtYxU//FFHIntzPJAN6WIKc5enTdgh4FA3nlf01DFcK5V4wwXDTi0eijGBlHV7
yG8G2pSNpnulJwOStmmWc6vRUkRjZ802UDz4/bgoUgsvuVgOkzqwHwZ1qeMGMfD7BgnPIYWxUTbf
BnzJLjs7wXvlvO78g3uVu4aspmBN33Kg8/owKgErJMRL/y9X+fUh3WlGzkOIhHbpgVQgvkAVJ11e
uZbllzhjFdFOPYncRqcbDjgVyChY7y/ZQUG/IlxgN9UUcIOaCSCQ/CqcskyyjqOwgHxF0Z8vJy8P
8OwK1P7WR+DYDmrevvlEXoq7A13FFW87xKGgUiE94XHOiu1c9y3ofpFfSEP9W/Qk0PN5kiwW+VDK
400g6kX50bwqxGIEMaz8GXR3tOAMK33u37Mukyu3ZzVgRgs0ZFrtqTs1VPtBFEYqCkhlKhm5y5Li
erhC9vHxAkdb5XXGL/zcTjjsESKFI9gmDP3mTxvyT+zF8A5XyH7ijSu9YLfshpdeziUS8/FHnJKh
9TAAJCgswNLS8XtTC8xRibD+V1def3l31JkUWI/x9hHqM1DOALHGOFNbO971XwBOQsZZ32DtMtOG
NHCnIOqeJfdFjEIXz0bc/T1p8wv1x4VJ+COSUkqfCA7Ps2aubT0c4+WMBIuxchK9ndj6GmXBBdAK
zoZajUtGMmsmrYM56Fbmo5AEaN+DfAMCRr+HPnGFWx6uK7H02xLAIs91DFG3ChQnmekl0Ffa7aSQ
Pxi3gRahic66500bTLZPvhz6tfygp9ELZCWL2s1gmoEbOM8RhD4KpTYyGRnugIb3i0Ct0f1a9Wx/
8BE0neT7vKG2RjyNXTgpkfKvFpGD/+LFS9vFnpLY/W8GgGfcnQIMKEEoPzS9Ui07Av0+2qTxeqFB
lgNedBjgR7PAvDbrGeZcsJ6TgSDOrEEDrTGeoyUxSoQl7tSFfGmnD8VjolKmMausxtTVVGceTSdG
wGxk0kRQY1KI+XdQmC0GnIIzbAgM4/8OaGTI7Jj7aLvveDUGs/eJjZo8yDXNBN2yqWWklDLYVeNR
M5phX+WWCniGUM8s1QVH8wJBmEXdgf7iR1ss05eLz1+KvPUTeKZFnsiJSo5rwJb6D1PF5NblojdI
qhZtxAP97+hoMLQH0mn/Z0+6ww5zLhOg+XtCVQQhX4SRWaUtbvyKOmXLFVkUrmvvDYXfPYD0sd7B
3oRUAUY/3blwbK+LbojQfMnFhYb+VGcULX6v+HvYH0lzyixFStxol5kMYjdQ6HPjlK9n+fxv02Di
5NtBxzyq5TRTD1cYTzSWgztAhNnMeh8UP1jtMWYHbdUc4JIc1gYhd9xNiys1C9Mx13cO4B5UAzUZ
TPK4At0SlkykuTJF+My1zW8sTAMLvJRAPPbLOk2BiOCeLU+0WKE/WqrVRMX24oLf03kOtfE9HGa/
Npy7JGRvScD83MW8M1dkvxbsU+2gs7tbNCDr+rJljLuworFjvQzSc9A+N3mSMhBmczf3VLEiI0yW
1NwQwcgKKTG1AvVJdAiPsTI/kUpiObWug/qyDPWgfflr8yimjOZE8ss5vU/6YiC3fxgRYSVlHSVD
LvH4TOwNyBX70GorPQwhRQkTOSKiRLE+delkBpoO2BslvNo020vz6Vibd3+g+FlsUehFBOkUpYBA
utm+K/IuS1KbavH5Vvp3FIG8dNgFQTotkzOg89tg/jF/1kOOb1DnfEomFJK4ArKrn6ezkZSgSkgG
KTDY9G68wcRhOre8+XiZCdcpxq3RRzJCTx2lGz2NwMfDf+PHzh+5cjgm1ID1csnsFJqRzM9aWUQn
POVHrGYZIhfUIm9Vb81b7ZTkXbVdhfrhr1wRoV3TvXiZDlKdDZo9LgiUw/oSZQO31zAQZvxkSq6Z
0OPhVIbVRRxB2ixmnxYiFMKpmAuw7QoQizSMCsEHrXNMff5t1i9SUXKlkrMmqHpK25+BcHTuXb1N
fF1LGvgWCx1rbT3q6AU9QvBnxUYixVoPpAL8dO6F5RroENWngHIlF5ZIzrqh2dxihIAjFkM6Y9ix
oPH7ys152ABUjCn/roqy2pagvPx7I1wL9jneLW+5Oj7DqVbgN/3tAJfoPg78pV7vRq6Y7lUszSvp
A/XRV5+FXLI11ULbh2n0Skz2IsmbkZSqj8bCqQv9k7zLS6WsHveh8FL6y2994+oYF+arjYFm8+Lu
hCC0XNKMvqloDwcR/A694RgZorbAvV1b8MUc6nfMISZlW1bJQ1APQMNuljPFu9r+tPaYoub5ANQm
jFTGUlWDV+pisXGTmnn3t+GIPVxPcjBlLsBDNuT375Ig6yB+Q8mUIEYy2jw9gjZduwso8kPTsWee
FbwMlGgJ7X8fSA4MLRGiXn5Y8+f5UBHjUpoa4CogBNGglbNVvmIW511kTcOMYw8E68QtH+C1ZVrM
bcxjwlLf97uzDPePEowwYzRu+27F0hOura53aSHsydFMz98PFrE4mowDlXTQZBD36e91oClctDT2
TPzZHCV2VJ+MxOba6thN8t4nZ0v5g5b71SXaRIbT7iBYExhZDCbCP7QiiXJMFmy8WoOYW4W09tJv
KIyhxgedOI1LIMdYrVOlMzIHBlTPe3V2/+o3tjt2tZDt02VGZwGCvuRRmePHvXrD88KFZOOK/nCF
PWR7YOz1vFUXq4HOMUfS4jxelcvCQ07WakUbExCvP1jAxOeX7PtM42CT4fMbll9FAzhDhkBt6rlk
8Mb2wn0g2G2jcf7DPOoJKjUjbdIvJSG1nIkTnXTdxE6qa1r7uyoPDaCbUw8nGmtyI37OSkuASt5J
52t9juR4E1ZIp7lJZpmkvPKoKpEefUIQ/9C2QPRMVqC9S4E19+LxYZ6BkP3B/1MhxJz8F7pwT6/0
0ejpj/5evEN4Vy5qhlYaWH3erX+YZnCTXEj0vQR5k/G9QbRw0RH46T6D7x4v+MMONf9SKKvU9LV+
edIoSoq/EtDoCbWcPLDoZARM9bkvGQzKUom3BxB5U7+NjMFn9/qQQIvbu+OZ3QQdMpCoSStoFrdj
sGOPgKJjHTsj+zJaw3hIHtiyeOLD5rAPoWgTdT1ofauEgbl8tVrpdUe3OXzSJCisCuK1KazCLxeo
PRraHUCycSttaePD+eh6umazIpr70ZG8F4SQx+WhIxZrheY/4lNG6r7hXD4xbBlKVFEPBqY9QIj1
66fas/N4l/pQH25wMX6BLnDDQ/lAtkCaPqYUGSscnZyTMlLbM+ss70B1vO6SJSGUwE13CPiQyYbh
GqvuXDfjQyXZqtsCwuWHLIexChAUvJZNFBoix33WfJ/g220kySll2ah9vAiQhs/Vhu+xysL/ajzi
ud/XRGR5rDz9J5LnpF2lZyk+TPwiQ+hjxFlKLN8jn0oXQPxVvG33CyoBk8EtwUquuzxkPyUSXYtB
+t5amkWyUbIc9897RAE2pXOrND3UPAeQ+OjpKlkFBaFfHISUTwdwD6G4KJjByViifqamCVaabt9U
C3W5vwfoegd73fEknYc1eL3VDCve9nJwYsj1/1jQwwbojh54wodKHSM+RX8Ovn8WWieRGwi5GGLT
s+/Zr7YWQ2rcMo8FiRIlr0JXrnyuBwQEGYIk0asvs3p9j7c1gid5pZD+ITv+sIJffzv9qlB8kpxu
D/rNaSBDXBrwSX13ID9bQz6YoGalt/TsydcTmRW0+EJuvKwvUKMDU/knQAjDDyQAAAX97Gc+Yvfe
RHx6glHliPHr+5+lWqlacJnvRWsmr7yiKd8gM4Nlk0Y/d6J8FymgLmcx6CADkqEg0vXawxQX+exV
pIlKxxI+j1No/EA97p0gst532ZhRaT4rB32YnxIWhxkvJCVbAGFmYAxSg90AcT9ALjg0Wd0PbnEU
gZ1eQ2yCsaRDsEli5Et5XKx+X75T+dMNLqsSVIvhgvej1ennGqzb0Qhu7dECoLPrw4x83Oqt8SZG
9betHxUSuxZ3L/JxS249WvIGHJSvMFiT+BkEfZAKxCanjF+SLvil2pJDYtEfRdAi8mjpjaoMfIBS
Xn2YrsDu4z8elzAeDpHfZ58UPQOSfhgH3snXQd5+p9n28wzJoiY7hLoP9DRYctxQn+iYQQz6Wheg
NlSfkJ9T/ErVfqW2iCIsq2fRUHf29/zLTFVMk1SqKRwtrCaJyledcjP6Q7vhiGgSOqHhooAuOMks
FHVmQ2UKv3it5lfVBx4KPEByWPEXBs1VE7UocrI3UZx4UD88tHR0JZ7Ml3cwhKV9Kqwxlg3vsJqY
2La2+o8eAPwt6/HMjhHOkdWf4TabBrrd4WB8h+JuUqfI4YcBEEIVR+h5HwD2SwJ90AnkNJ/F9YDo
5RcsUg4oWFTNGPn7ckHOtTHI70PpSDRhU7yNX5qOtPMWYG9GbFzQy45VVYRsp/E4PaEe0dXR6RxG
/pnt2XhRuBOKg1g6dDlSDRCUVQd89LbGxI9jYb1XR6SuMxoS4DFk4aQeKr14BXJWXSBysq7ovqCI
B+CM+90zyNupUCVuloKoJDv1RKL/f6WXhJawvKAVzShoeVQVKmkCbAxxLMPk2XSo5n/mfS+eM/kT
tul2nN8aibvCVQLw/GuTjlHqrDAD/A2KQ3C8VExHXqOFrYGTVTWunkd4Sf+JtO+yhI9wOi05fosw
2IMxKCvCvM/pFtFTdFZH43e8u+qunyVzQ+hauoHlSQ5gVyR668O1rMYaF6zZryaDVpAIRnvLEwiY
oBrBu/I6hQS3UFRky7OLHxo7TFFzvyAZKpo76Y5RPJRUOuXMILmKNwrOQXHcj4A29969kzyTIXV6
OIUIRbGzzEvhhv/qwFoDmjm00LU/P8zQ6GJ+IjZqrqqdKOsO5b7sR5yFht4V9iXkIR5G2myjS7XG
lPxOXu6Vc2oDdH6sQKyyRRHaquGqon0ivWQ9ADaIFWnOpiVFe4IyRLODJIoCSd4XqUasBRb7JfUr
O9ewHo4CORrHaRxrMOFeLVF9YjE500+AXVr0bwDAUINDmb3piECAq5GoLkxN3KVwdghM78Dej5IQ
N2AVXIkMKZsiXXU/e9ru/7NrTfVSVZTAaI4wvJYVVwodeR1kErcW1l7oRVB+aCizg18T60iNLkOO
dkdf37k1ZF8OjP7MT+9RRCOqJOTexTvNMxSezT+n7/yuEiGycgA0h6vL3B56qCMIQtSpQrNtO/Td
ZP8/NSixF2E39xSQB1Pd7rxRz8G/mHFDmouvcCrXy8jHeSY+hjyCzi4TL7986MwvvtJhzaAcwr22
vSp/DaeQ5jKRYvh1poKP7V5MLVL6KWv8z13aNFbADOqYH5HpglF4qB8KpxhjCEIWnHM99JzdcJIs
bg85R57b7uv+41F7YPU++tEP/5Vp1e8UXd2LKq7Q237osIDAve/gdtPmUR/xbimRpxitU0QS41ZQ
cvx2VNwiEsFb8jCJ1AkYekawwNhAc9Z6d1CDJlpibI/CKifjzgJeDppMMMu/wNQwQfNHnDGh6DxT
IVni8pjVQZlIHFch7RuF1lTUH3u6mwtTLd9jfKySqLFat/VCNA9XdhxGCE1x6QDF8LTexihhV4Mx
xUC+WZLwpS9mAhl+ERaC2cpEr9V69eoUtwbkZQkEXw9GHbkGYsK7LOJml4lqBiVeQvmBH+8hIx42
QBS8AU7PXPxAaYee7qM2Ct/whtXjjHmYe+pNF+3DYfq57NxjZvJ5+2bAY14XThhUHVHWnwrMNR1n
4UWuWr6x9A7I+D0ah3v95paTemXSnd3guDGjKjOw27/+ojVFPHrHd3iF7g0Ofh2aREm8IVCXKBbK
wlVGB9gI7rBJy+A+VvKm3sxL5mlbeUeA8Q67IqU3wmKr2Y0GAGu6wwtDvDq9LC81mGsYZHZUWuwz
wCzp0lD9zec1zQ73PzHN9YudtxshKSzefLwl39loBujy1tOEQbMaONqwASKU54RLRROss0M3iEl1
HxHM6DbBLhOg/7e+EWIjpRbXce0EW1Pfe6IbTj/pXpyoIKInrRP2P/cPoThU9tZ1WHGkL/vW9ZxP
e6AUSN5/7/V3L6L/g71ndnU9/ZJm02tolGvBIDBcyBPrj10CHuzg1eD+J14nYTVL6/Y+6qdEwNt1
DIU0AXWBkWmQJnr79IJmT9nXpyJXv4frgQfq8G+rnW5R9gXv0DOdU81U4a/5NuQB0eZxcqNOTHJK
ztC7AR0ua7GWB515flGqHQRvqlJy2bmmUae/zBgXCvHArObOZ0Oxm4gj9x+TlpvAxqGsNdwzyvTB
neZar1YqLvFYcXjbYsrt1roWyLxkqw8f4k1XZCoWqMOMvBQ/NNXZSDLQBO9akGddHxUHiZHcU3Cg
crSWkg1RnofMA3FR7xtHNwPkz9lVBcDSMOG5bFLwq8icuETBJ691ITAZN/BEbpxc7q1xVt594BJV
y8Ec5kGy/9oow7xXS+MP90xVqipkGvxupwJQpQlPOEagm0IDh3kNcZzAiZN/vb01anLvrWC6tD3n
PIVkb8tE3HAjhRLpbLVX59DbeehItjW3n+JbH0ivPANXe4JfFkDKTbc279yyKObsfG+u4Qqt13wC
OSHBRbSGeDzHTqZcVFJzLDRDISGVJuh8b0D96Cx9RMrnOEyxA8gynbIUvLodV4wZQ6sgIUaz8lj2
h1IzaAMtiaQksypwEnjon4wNU/3ly4J0NdBdcWkD6ZO0mGXvpvppqwqGKOJDDhe7r3BYe4aBfGGi
qKD0/rvlKoPfPx85/JP2/LiL1/DO5yg9Al44gmPvzAtbwJxrPMveOvXStE6ytEIcEOfcD+c1zTrQ
GsJyWcTM/9jmcGBxX+gbmwR4N8YpYZwkDrlNmm7UO1O+XoZUa/6BqOo63qTGxuHnpM5bN3BfMOdl
2o1Na3u69DEtVfRnooI9/wMl0Hc1Lfuitd6W2EbuzcN5ESDf/q0/+6yriPyN/q6ZmPT9JaPD1Qdd
aUGqKTM+OVmeZYr9Pz0Z3kmqRI1ZtLEUr7ttej1ni1hdArh2g/4AaNHZ6mDQsysKEJDqM+HwPflH
OftnOWtSNhVUE7NyMu6b5s7SXVcYEMr6F1jiqijqbv9LnpD7Y2TcTmvLTKwTV6NXUx56LadUxhGE
fwJaFsfcik1D9su64Dc00MubrblOyebuSHYToZKNCRRtSyh08S7/SLGK710E8NI2wFlbjnIEQ2Yr
Ondk+qYLHkuioJR2sEmH542w0Jhi+Djb6TQ5C3voHUyEeLcQra86kUcq4NKJcd8xppap0NnHSZoj
BGavuUcKUkP/syzB4Nle/0jGFFTlE1NbHZ1ff94JCRrkUVWPXR85pvebcksBvJ6l597PclkHv2AB
MLtQU+Gq2SA5EYUruyaJNx6Z5uoIWq60Yj1/wCW3Lv3Etki34w0XU573KrhbOkJkUk/YLzjp1YKT
sbCBUol+RZuD7RXh7mLt0Yn/VUOtPWfkROgn6sUOafCC6zD8Du7WVKQ6jPoLvBOd9nneVf48HYPK
5jZTrxvNfbQpx4ZhNN1iz6dMhSIJHpAJWepBEEOR3QovJDDE4tMjLmorBMQm6ErdL4h5yP5UnQx6
5R59eLKSQWI2b4YXzqOCFdgPwm1/UrU5Ksknr8g7PL/RY54dwVVwspQtO6XfSlQ4S4695nBgVQGq
17CKt0BjkXh3UgQVjbeRR8m/lTrkgHNYjJwzUyOgQJi37/Fu4Z1NuGhpHCRWbaubfDEeFOHAu2eU
t7Bzd08VzNVRm0j6Dh+T6YQWJjGm5LtqQEUWis+nne0fUTJX2ULwEerT0gE8Ss4lpCeRtXx9IaLe
/CTecMiRmNtWGCJreyXIvLOD773xztDB9lad9iOXCe/HF+HjLHrVan3RvQJ0JDQJyoxncvwDZIWT
wAY/rH6IaWc1GOY51Y/Pd9Jutx4vTS9MAhGvYbOiZ4s/8V4NLFJQlqg5FMAm/FFv9ctyzQkTOArZ
dCziZE7NoRoElvc+iLwfDXSur4h09wKDvbQj6JB8VaN6GLCOlpDVJJ+33ovY3Tiog4+KA+iN7tPP
vHkIIvp7pq00mtGbVPILRG7of7AJPgipHDyTeAJRX+9Wz56mRF7TSQmHW/1vqAlI4lUyV9v1bjud
T4dp7KDl+/jL7sERWIB2cc0UIxBgIiOdXm/ncpU30LmeIKg07r2WOh9PsokQViF8Pxq+vhljKDty
bDEHI0egV5wRnusAH+dyjDwqXjC9fWqrZXjuL5xZdnaXfUMVAJTdf5TqOYnuHHKbNRzzC6H8I4ax
WjUD7K6bRcLDX+bi5f+DSRBG0/N+IpsFXrrDk1o+LP0PNq63zjO7gVn36UAkA1vSbvKyRcjzjxp2
d7o0OlxocBnMKIr4/hCX573dpcnrIqStTjoDhtm6TmSMN9cBxL+QGpnX+9koHtloT+EYDyrcvWZ2
d+C3/bR8ZAbDyM4ECskBe3y6FqxqCI05NfIbw4Q+7koCIDiwLLSnGf14z5C+rfQNbaM3Fp+41oIv
vpqftqkiMq8LWLIMI6Icvwp7dljFnuhJg0jgYyPFAzwcFtVvCMqvSNC0RuVcDENZh98lrX+fQ9jY
aXr/qvjwpeQzQY5DIpPIhKofLkUYlwOx6Uw2oBd0ODU2C9FOeQT4JZHQbG573SSGiuLzXHhTwdCB
ykYPBj1kuhYt+7JzCPfZh7mmIhYvzLbq01YA1HbL06pknN2XdXbxlbZzQdrbtA61BCFH+KJRFwZi
3oKRSldfRMu3olAecjQgMufioYdzzLx3wGacexWkprtQ93dFNaFjvFo6fddApa3mHxsAN0Ua7Spx
Yon8uYzKWs3bqPdc7KszxTuPhh2sXkj2vYmwVKo6t2fyR0BpvmCsdOFYLU0fRu3BNg0WZrvIVnIJ
1LH+iFee5qKh1/vInQz1YPxEo3zIFUBQ1Ep5NIKYrbQRwqGR4Y+RsP75bhlxdksr9oJ9S6JGzFTd
VM+Ej5UYTkUEG9nKN1yJHBZOxJqGmdNj+Vcruwrxed9r7XTSI0AGfk4dHl1xk4OL0g5sreyBTNG1
efQDfuJfmQ59miUbFBaoszBIp0RBbW80vi+Txd1OhLCsqRQ/eFIlhG5ZJLOruDWWKEVqJlwA2lKN
3eDEX6VPAv73tOCGcwvt6kSjuazj9LFxFQRJgVtNYXKfxlrFgjJpTTlT0FoR7AE713niL1JBUI24
1FN5tQJ9ogzFDPjcDLmKU8J50zFtqCS2v29tetGb7axDwhJuZ1lDqdAXVdMyPnjhQBwNTmVm6skL
3/p6xsq9e7JW37zh84Fc8sBr6qWfGi1xdZAOLyFRTIssz3c+4u5mxPwHKNEQbEGgX1O1ggaVwNvn
rfB8QW+11yIKNq85KSF1dxx6CXD4a+C5U/0ZbQXkDxhH+8wcYhpHTpvJzYyaYsVlewcJyTtTqj8v
RT81lWOPSawjVYgQYqjE2rizDlCFxvCOK9772/DuBA8AVjYR0ljjYKL2JE+YmL/7VIwSJ9YmBeR9
6wlIbRghHEJRdY5saK89QXKg95Gv/VrUAHFfr2VKpJWGCAtCpGg7pnyvg3lrMtv/IUvBeQGpg/YR
+ayu6IScjNQJR7xmhrrPGSQOEWVQjaOiHgWtoLCCh8n0dY1ojRRObOyRF9I5C+12ZiQvWiQm6uhz
qAkdljLBz2Ni7LQHU++5hImB8gPqKms7jtkstxMfi/lrmQcoiQ3G8Z+gPouRM6Y3tYOg0LsJsvp3
xt/mcKDMfVgWtvhxIJu0nUnpnDqxkTM0qLawpUbrwGayq9pRFqUCwzVB8dn7Tp/S7Q10AgdKPRVY
EK8dHe7HtydHdCwPCNZ6kj7WADmfg0akER6stRHxTwpKZs7OYlN1cpCYereUeqbQYMl3sfmwZce6
QOtyxkD/SiQAOykIZftnJwU5ISyVtE92ZfaCBqm2K+mPRchrT7+wInTGxe33pU32BhTFK0Gt7BKS
+Vj3M0CjMSTAYoVlBkaHQGtq3VbLF+Pm9FMV/Q26owvKZFQNqbeDJFlrPW4V88HKwoZhFu66HbqS
EmOsHm41ChEie7w1ujzJEv32hvdzNVrPzTX3/QbifRHiFxfurSPIk/6fnzrQQN5NLoaAMexol6mr
1c70d4CnAPFbS0iS5VtlBv5SU01TvJ+9CH8bigos4tf2if1VRg4ef0nsGfDK4nxQaOG/4ZixbQsT
MqhKC2DajyqUwlM/74uX4NkkPK6tlZEGPireZZK5TaINpPdXRLUlctcVDHb5gFQDLNhgA+s+XXJj
+1/bQUu5lTdh3/E6NANEADsVyBDjMetWKDpVxoyu2FZ6c9/3IH2rNeZMbsfhMcCMpVxTOMoH34Vz
QRLLdxVGZqlzJGBIEb6ZR8+73JnvHkSRHoMAgUPpv445+wGV4LwW6Z90IYxQZQine8YwRwkVg3iS
Dl6pyTFoJV559yKpCOGmcIQU1/BfFDoezUchyMUfqE3oOKT1eo3SWCvqZdLKtgvnamPpTRG6REoW
pfpkeA4vJOC41aisesMZtGmnduJsuG4p3No9NQfzNQZJ3PJCefVRVw7LbvMHbEZdm1myWXh5fwOU
AevPTYh2+M2eHGS1lx+PlB6W1K7hhSkTfh0zNWsLgGPu8Wkujb3BBSR+HW7TaT5o2urW3zz+K41Q
9cURXcs6e0LO1cnl3z9K+9TMLIBkH/dlr7xHz+ir6yKEeUOC5XcN4owDetglT2ote9WLCp9Qov3F
CuInZANVE45x9ubivJRRUGesD4VX2ypGQcmMws6dvk4At9AunsGJtLzCM0IiIXNdO2XWu3PE6kW2
48zutFdHVKp8xxhmZOvbw7kS/tw96WM4IbBJSrUQc32E/gC+JAz9vby8NeE/RdJyj8IVuihySik6
sLpgSZZHJtr4ZDLq11br5f44eC/8H3TTNcg6HkGoHjl8jvcwwgq8sswfYYjZw9AMTD3qHgTRicEB
iFGQIH4QE6W18KvMY0p3gFIuaeXYAX3eG1D0OpszR/GBZ3W6ZEvdbdbgXFsxnQHJstP1rT6x4106
3BeSgxOizYe9zwvo1F9ktMUSudLKg8/cMXNUz0d4G4l95+/qUB1lKJrvMy3fdpnXQeiHxN5CbZFW
sQoKGSgPvG0PRgRNikO7hsh6kASkrqZjTOVvYMt24y6wWTXh0gsUWcaqHMt/zT8g6lXlLoNCnrPC
TQgZdQlpSsaWCMxn8G4HtmkVWk1tsT0J5OtP3oOO3JABZ5YVDrqXoa3F7Dr+N/aePQPFQZY8LuLB
hJT+SBR7zXf7pN19Lubo1oaK+8DZ6qVbuI2UXWVIvpMEElBPnKSJscbLeUBKCZKM1H1/x3EOAzBW
X3+uiXVnYICu/6OsuqJPW2zuA1KE6Y1uoOB64N9zhGPM05JydgKOn8m9LK91ORfhzlOLGwWArNgc
eIrQ42wchH0xxWweTX4iZToz5LmLlFugYxlK+XgqDSEkeEhiz8UAsQElm5N4dmk4d3Uovj8/njuq
UEifzBsFU1uUgbUNTfcNffMgQ2I4aCgIscJQYiC3Zs26UFIXftqGXbQhYLLg78lY3GEZzR1YpNGG
NrL/b6AliPZnZVuNjxNmLkymjYfwOODV0rvv2HfoKTUhCVQx8ekuQ/mtQEMn4lh6iX4LiQtdU9De
RPqQtO32qT59OIBeYbOO/IvJUws/OpMtUhglTkAyV+S5PGzw0jnsgeAQFer0xK5puQjdrVZdXTXo
bh3iBhGxugae9uxhN8wKkpkFMfR2QMqLaerdZWpFEFPfJiJXwU9wRYcfGSiGCWn53PVupdS5/JWE
kH8xZ+k77iT7seHJL3L/J2U0CKwDOE27ZZpHyZt1bXLjSANoueLAlrH3BZXPMthhzYrjRLwdFOQ1
cTVJIcKMNenlPpDS3Q0MiMTGMAJflUwtZ/styc7Ck0+gS7yinMA+ObFG3LJ3JlgrQ6wsbJ1YXLhy
XptE47Or0CIG+IDpWpHscUhcczMKtyeeRIyH7cb4vKLL8h3pGYCe3t949we2A096tVR5Hjg9fpZF
vJnLMiIGngQu0yznOZMjElvDfGjbJOxyDVhEg3WQZYB6XZAPdCedN+yVXsC1g1xkArbYtZJyjgQG
aAEMTynv+i3CPQtUDVs9gSzYzw79FqLWAjn8RD3brwdk9FZ+6Dnq9dx0BQjgbc8zvkGqDXozlq2A
lsm+IJeXksat0KM3m9M/hlybp7jjCI1FVu04G/IGEQRLPJOx/97ZosHXRgoSoLwTMZIZcZMZVJYB
g5DFkuT6n3p1A99RMP14rKTRD8wOo8YCpk9MB8XMmp5wrlAShiFOE8IkvnoU1JTqFPsJUYJCfcfO
E76j5qbnfnb1A0iFXEkvwyWGGuMoffjQm3nKXocfqAWD7jUKXXGazw5kUdLxcfUzKKQ1tVUzQqVD
GOt8ewvhD2D+CrMDSfEpUrHdFUjcGqQneIMlkHAWQoIVGTQntfVx0v1rv7yizWE04OHBxrN9OCqo
J7ejKqtybCn73lQtW08c9kvYWrV13cOgcyDKWwNXEO3Gowkj3PK+mklOvccLKpVSiIRSjzHtuKzt
XjrzFrvHA2JHAUgI/lUgBcSgWUWEnzY7fqeUvU5166v+N9e6f/EiFq2u87I3+PW/oqamRYR/+djn
RGmNrFFktjMjGdJGo++DkIUeKOIX+ilWxIa/CTh6AIfvRyEJ5rd7jRGF5klaOHIJUUWNpIVWBouF
N22d9u9DV/dguyJ1o+Eb6Ng6DZbfKtpIz1GIYIkfegNqAr3qtZ3EBy59N8ZDo6ChH5Xv+3kTG+ck
aGpSmwi7HPP+h+lVZAg7IZtdIjs7VlDkF+L/ydhX5E5WmjMdG//mx/d1v9aZNi6G4qHIIDVsDtDQ
NH2oaNsDVANUOUTMLOnqSN1iCVyGgDj2ayQ7ibN4l8t24fNj+SsJ03xFyKWGsasC2WJXGVq7LwuV
Q/pXVHgwvwccitsADwMkneGuYiTJttAnJYDtiDAqycWLSKWUGihha5HNUq06uowEtQfAIqra7fav
2pu/IuIu6Wbfh1/i+kTngKAzijAhQSqb3X3/Zl56VKJJoFPKBeG71ubgr+68pWNOe9YPFWgG+aAk
vb/DkkTuhbdVke35rMasYTtNcTIhiRLK12nz/ikmlxOdibNsZFf/NEr4xs1JXOEgi6aZC87q9iTF
z67b+0twjZk1xolDwQ5ixs9R7iCVyURMpZqoVTqiH/kLnUD7HX7Ns48pnZDApnqlSEkqVYYdf9du
kPRJC7iQG6A9z5Mj6IIRLLeupshNcCDsGx/SYdINTwYPkrR+mKHFYkzB9UZXTKmF4b2mJEShBtIg
iJ8sb6zZTd+af9JuJ3WppEcjhkEbFy7wflh/tIR2YqeVb41zGJGXQqJIrDpED59K//n369wbD6gT
azonl6Y9zwip4LzOBe269tvZu6gIzB+RyYVGHRex5LtByWuHzIqZTooJ2euKfhYh1VYb0+poe9OB
TT4LCl3AnH6Y8PgINVHR6ruA6eLVZTDw3ZJ5L6VHegumbeTc66rcJ9C2wzLmEI2vh5tvUdtTcjXf
6DiRA7bAi/FaQ7NyOSfR1++o94+FBIym4ngqdCdF9QgH4Ug3KkNu6SG247/jMN3cEgz78tIHtQeP
XzIt2SlyeyNubcOpFBij3AaLIm9Czl2pRfhzM/+KjiCmktWsSRO0yhXp3xLP35sJ9KCk5h5006qy
ZjKHzrsEtPHerjah47NIegvnhe+T435BgJR9qPk8awVQKnI48LJNeTIVClbIauUXYAV/CpS1H5/7
2kkaFQGbzRZ3l6GxZWdKzdxVYXBEsh154GUmCUv0MzGvl+dNkqrTL1w0gPyoXIclLuQ37b76XuoT
+6txzcxQ85R4ysJhzh/ztRzNOWLGAQm29WdiCN4MEj7LCxx4i4x6UWZep2OOOdVbOT2L63W9VV65
o6xJ5d2HUt2AomZEVAghFPL52dip09ZcuT1yfmGOuFXhvUoUR4RUTPwJJN6yotogP3XkKOoinruY
u7NhqYaPTaHevAqiouhlEwCFd3ZlgaEerNE8+g+HOwBIGOF/KWZWx5nRReouj8vp9yfPJF9GXkGa
NpT9RrttCalo6X2ExiUSr65Wh/LFDpXX0Jmqzg/ttDk5xkiW9fl7ryd1wYs6ba4Xn5vNAyNL8Die
rmqAvb9MfHav6olUf4/mzmF47+qyibZT+Sw8fh3hUvi0QMQp2NJZDXQemGmK2KJnjrApOFViRExT
I+Jx5a7JhVJWo42b+DTcGL/9Ujg3aR34W10J5VgX2bZpTipFzppxyA4EEsTQKimG5fhG+qtPaDYO
pyyDYzf8m+1XnTDVTXg90xlC1eUZvn4qOVIYyN+YnfJsCvGJRQ3mzrwXKgwFIt7pjavCCEEjzsVy
WF2ngVpiin2GLKrMjzxNLLOu1YYNij+6MqMqF4xiVfauS6XV+MWRAHah3lfMr6gYWvWRZP36s043
o8RcsgdXy3OW4jIsgPt+IdjOeH2Ux1l1MhhIqOdf5Am6DtdCzBeu0dYHO1K6aMvLg8cYxVsfxQHZ
61DJCGyckGGqp0Y+sH+xKc64i2CPFsOkEcB+MOX7Sq3Js1EvyH87s915xX4zU/lAUEzzlUuPwIK3
fvrLtlXeRnF3Kt2Lww9gwV9KP8pM+Y1HMsK5ZySoibohQ1Ucv+ILIZgySGz8iYIDAVBesafPnU/h
h7zLvQCiKvzNLEMmLDBNNd02DcBzYypThUFUJsb9kM6AnGhMRU6NH1fSZx9dewjIeo8BO0hrPI+r
hZ2QMx+fjZod1fRKJdI7Fn8k3xYQZcWQZRlNMbif1A8nOgKLw6vWCBCjbjZzoaf5y9JHumoYoyXn
pKDdVeiunGbpP0qkFbE5dAjUMFisTG2xt6yyxmHYlxRDnitJCvs3Y6seb1681GsVWycnTZmZX63J
LzTOao41uE/+Jk/uc10OnijH7WSlmarzMdrs6nHI3pAODl2p2A6T1aABzERRinliCMBw/Y/P+77u
yNBemZuPF8CoE8modCdobNwnYqHGCIuTna/dmdzTOtXCVm+90q64KLQ2RmczShc4d0adAkfRS3zw
PGZPsuknObH2ICJItqDeQ935SK1OftA25afTrBApQTxv+dxS5oWK5b/No5M38AcVku6RFMtWTQvF
9jPH++ny2HBKsy5WtQPJMdK6klTQGxguD6aoVUuZ6FgbALrMTHjy5pYekhmEwTmJxAmN9Vcxo+/A
zVTqHF+0jl1pv5ZU1YR0eIqO1fMSEoOFFln31gLZ5FEX8g4V/t1023AS699IU7ffsJZ+qInrZpt0
FlKHva98y+5j3wQ5rBy1tV6gEdXxn9ho7tP9la9oexX2Y1Tk61IZAPM7kruB+347xe0LzRVksK85
JLsx5dj8TX8P2MDpxWV2Q7YqvJwMHSMrKNzs/RqLS2I9q9DP2gO8YzNfS6NzcTGGGp7/lnwS8dET
uIcdYVBQrFWRLKBKDMwmF2s66oC5FSyR1EuLwU9p0IRt+tlZRsCCDqdeKk3bpmU3uJ6Uw3C/3M6C
rgqhbCQOZWRI4KLx3fsF/M9i6/RZ2S0dkUr9cAGb8svxGtq4wXy3xboghu72/Yhoh9gEN6ltcZYG
oPkbpNAg21dauYg2WDIiuiTjS9bXYENYshdp1C0yhSgsllzmxoAJmQi3Tv3GsE7LJ/VlKuqRtpdz
E1P3jdU9F6B0nXWdekZVh8WxTN+4uDuMKK2T1XoZ1vkP1Z0LcVPJiJd+U+7TkG9ddGuq+gr96r8Q
bI6g00qRqovIxp6mW55v+MCz4GeOWzvBG6KuCUwUzf7TpfrAYUlP/pYTai4ZcEJJs4eCbyeJ4AhN
DUi0vLr4AH/wnGobEn+Mam2TuudFOVNZX46WZ4m/boBz8ypYmuNUkLbxdDpQRih58xF/XoQHNZkg
rk262umo10Knurwd77GwTSeEbeCFlNe93OnUHTELPpBViMeyj3c7FzufAeicn8p7kqztSPUWt9Yl
PZ93VE/CnvLjVSsdEkqpdPKQyvvE7V9yUmqF9aTXbIYI11TN7cjWcoq9H5jKTVJYb7I/5gm4N3ng
E2BE2GxxY35JdagtJEc37un7jpafjjgsWuLMA6RnPsX96M2Aua1bVln4xqxPdQ7nfeyzFcYRasTN
p6Y9qY23CYB0pm9R6OjS1P+dojVC0eIH3Ak78oqVZjbjqTxSfL5YL/+u3TjZlw2pjQ3AyRd3T80D
jjefhn5uQi3zL9K3DqBTvLsGFKN2jkPaGrj9IQ3dOKqO6X8E6wWqTSe+vRDHpZN46q1+n3cfv3DX
5DNcX3VMZ7DTqAmizNuIpODMRi0Z1gLc7074WhS9l2kMgBu2f51cAPgXRyGEgnLWFz9PklgF8c9D
CXERfoJ67QWNszAxZvK2DZoDeS9C3HzXfvyl3Im/WTHziPSTDnRewdLcHZlBD0/QFA+Wm5Fs54/e
12PovaD71UIuYW17VsBmc3RgY/v8bApZyS5xncUFghcjl8pucCxV+qCIydKH52zWeldDG1aFfloE
zK3avnS1TamRHJ828rcoyAmyPD5RlokFZcVIZcAjTLhN9b9T1FtoFs+c6TjA8RtckJ93V/8+Sgtt
rS+M65APWZJoSC9TE1Vws1mMo9CCdVG/XPwdujqt1bGfJmS4y1dzn5Xxmu/PSR+TPvLHSWHUum7E
KoG8ywSOU4B2FnS54rzD+Cq7e0fUtb56UiO/AgM+rvcIwtawCQxJQ0y/TAGZtRK137n286+zKplG
36dILahuVyIcAx2mu66CoPEWSqBaLyduMy08B2gtMpK8Gnw+sB1omvcfXcuo6oo4HqJUXxA0n25a
cJTAgYzMBlKt854gaT7twShc2Esmb+SbAmvXF90Vj+ciA5wkHYozmIC+M0rpEtUj0qB1TKFJPm9j
OqVMAA2QA4PPEqKBc8UkK8WHz5LapU9lc8HOYR4p2fpwoUzH1vmOuiweSa5bjyXjPwklrQwCfAPF
M7iWs2cBkGNf9LY8nuwHZAP7CcKCBs5TjOkDTLdVehjHhPVhYEPvvRjrUkoCd54Qz/KySlsO+OtR
hDDuRuiKXqRIglN5pahK6ZEaJF7Sm9t+o4hVfEUV4Q1e72P3c8aHYUnECjKaxC3ecPhwKl+0ziJg
NgIZrRk4adJFp3/P6Nr6B8YwAHQFecSukaFVWCVi4tUYmQLQx5xBBsqkFQMH0fa8A1kZBjdaliKD
ymmccCkMw1fv6HfStsaDc5FNRJ5yec1sc2MXWBSpDG+AQJhAGxW3dX1v3uyaNfEiLt+W18iM8EuZ
33Ml0YrWdyc2QtHoNn0PxqBt7IhyMBfjMYTtlNEUPCDjpZCbntebAzyumsNTC05BpWLUAviAJ0AX
XUSglUVN7LCZBEd4c2Yz6vHOEfoWv2Wf/M0xpEOuzAh15xGHQNIZk0k4RSJToHmFf6KgleeBr3Xv
cVsk1E/Cq/ovXqXHMSjxYpjoeH7zwLZigI1ZlbR3Df8lu688snNqdDudT7fY5jXC8ZFAJYx7ar4w
ad+e8AySwwXTKEV0bz4p0NqpAZrHAw+qTJrZm3TZbzfgloDYXYhfgMPYf4o2sGPJwYWZRz2F6f81
3lRVBvj6DShnpEhNwXFjBO08h/JT63npD544bjsG+ndPAiPnnFUzIZ8WQ+Lg4exL9JQ7KuDJljsv
6hDLuMyx2OOiw/DyNAy3xtZz4RcR+63X7rfYnQYjFJTHATiNsD9uPW2v0BROTCO/Q79CI9+oC9Rn
yHyNRqioldzVN42ihwkLCVLc5HuuT9x/AjSFe61N0sefX9pwX07D4+E7fQDQBAYED++W1uezD5nk
RgUOLqCVPMU9tP6YfbLvOmoBl3FWMmOo/yiZO2wLE3jMnINVrphe6HBhxzUO5/DwQ4zpoKzIqOYy
pY72FNeQP1BTTmWu8Eb/QtadGJ85euBITBa9MNEsl+BfnF2JRQwBjHeSi1lVtmitTDNliKs5qgqN
sHox76lb4nYNwLAj6j7N5ES4eXM+A0pVT9TyO3jQvdeJVuiD9MDUAhRaycklOvSzzHILMP9ynhIO
taOwwa9CWkXGUZtHhj2aBpLZ9ONRskkd0+VBqe84ou2NZHpvmwvUhCU/FzlQttTz+lzcQ1TDxlV7
gOE/26TN/D4AqaC507ODyJPuKYT/NAIyeApYld7mKNGriFMRYktiaEOvLrju8cjap0/u3Er7hteT
u00F8kxHy1D4nliMyrIL1YYP3csJZJ7ZFUswIeeChcR7CXXzms3qh8JhoNRoq7ZA53e7g/pbtl3h
5hXl8m2+TdZZve3MXmfCd9G5OWwmMrOAUcyDKLmAZikAs9OAyMQRC2Nzpct/0RL1ZYiY5xdAf8jB
SZpYHUK2+Fwobx+xMmQnDxP8k7AwZJSJEPChpCNSoSHeh7rA5Hp4NUqDWaSXx6l1nIrE0TZQpZV1
NgmU4xn1TybHTvcmtl/zRKP2KEA2TG22XqRIx0yzUXt9nVDdHnRLqmdwAXmuSuT/TwPhyiwNybPG
bLFZ7yn831YQ+6xMhq2d9m6b7LTu28/va2tvK/crpF4+hDRwhRxQWD74A2PiLTnJ44Ly4CYrB12X
i1BJEnnSvg0xdZ87W1sNi0hK9q8JjLd3e/y3OdU2R+ZArpO9jn/j5zcw849BLD9j6Xr+Y4xiojl4
k4dDazvOr9mZo+FsnyF79D4zSgTH9Ft7V87JujFicz5B4tgSsMQE4ds9wtUPRREK8m5L6NWMUcUp
6NQTnlSRJDETqqP7VQReEteuedpUEzBMwAxHZ3CmK/1S6QT5LhSqvp7q16wMGW2uE8MXbG9ffu4I
V0udUwJNUBCmQvrUnvRvMfzb68QFH18vrwaXKIOWV7l2CfbvZ8iDu7Ugt0zEDdZ+/+dSO12+OlXj
qMcqNt9uiWQG8yGwp6jwJchAFbDNZknsSUM/Uu+irWJK9qWLg7pxFb8UBJrp2+Kwt0lzTe+c4x/I
TCAiugAZSgHbgrHAlYfExe7b2BKw0S6w0Rr3f3Z2MfluSSz9Z0Z3iqWrRiBqp2f/LXKlcmbXJWqD
dN1E8CUD2Gg/xQHCrKFFO6DiLNk2a7ePcwpeD56gGQoEsR5x2y9IYdnnUZHtlT80hEOOwuDxFK5p
9yRnsJp0QzanVreiOsdUoMSqIra+/IL92qSak4/7XoESDmB8cYQ4lKv7jG2dQqtVfgXKysxlieIK
hC5GuoG3uF5IrZmOsXHRFloz9akfoYYBtupkSTjUmlke9vMPY6pk8hWEMouEjG+93KSDKcGfR+fK
UVcKqEKMKq1/EyFbGLPMifNVRWei+5mJh4jqMaKE3/15sWscXk3Nt4+Z/8265ScdGcLRQvIjJ/cf
mephMxW87MuBeJLnlgcEio7cLJUa6B5ZsEJqmOV/oNNrogPMnObckoV9KzuWGi+bL+mZXK28ngq1
Avzx0ym8HG4JbCXkWVThvSF5uoSb9D8kZXgB+Ox1rwGi4YNPizZ418PS8gce5OAnLNl0S0mNJe89
OetSh8e6B/OLSzhwL486aAlJtgS5ohU9/vUUHXkcZIu7NgB5QkJ1UT0CzTGoTVZQirw2MqgIp0jU
wypVWLULHJz53k8apQQsn9NNcxOf5a6FHLagwvWvYvcurU6gr0jA5hGyoAO48Bs4JdU0mdbwXgiE
BGmv2DGncILoqGHTi7MEyx6zSjbNpTRWC6Lwu+wp0jf2G92ZYaoEZltnKCUrbI5vc/WmnCXc1MxL
NjtqsoREPj6W/CR+3yqhsYvxK+Ze6Mg0JkNtLjXu2UlvqEnglplvM13rMgv/vgn/7f0Vv/wEI5R0
U/wrk5VVnXodmTs//tAvM+wS7MGjRuhTzGvxhRcQgQtnSDO/7aRcFp9njRxvHY9h7CVwL9n4ehYF
Mlf03peIUUCrfKoT+VgXX7U+7xkg90XlqL0lEdm62meIgMnhEfEAQ2PpkIU6FeyO26uqf612BWUL
xfRE1Q608EtMnVQEivPY3slCKggzgnvBbaAPDaCHIzpBKW8nbL8jOxb1PGY7ssxbp9b5OQJr8tG3
QxFmiCsPGL8I9eSjnnI5kiymSUlKfKfnn5XZsMhVcKlnJ1kOC6w2EAKUDdI9yCLGfQyoIGnd1P7+
MffMVQXXl/syi7TQoF/r5kIFDumTmOdjZnHMzPFhEoxz4QFxWjHTbs+NCRG+GWqh4eKFLHIg7b7p
vnUCPV/Yg3ZRWV4zcfJh5aDl6BTn4hN0Ts21Tpx7xWXNL6DhuHtZNFdoVztTm3MbZm2XHVxU384g
s653Iy4v6gjbcxfyQ6mVII8dXiBF2CxYC4NjCP3i9iSfnDVaIWaeNJCrDod8g7KlII+au1Z1XxYc
kTlOys5juvDkAFlG9GK5kdlxagiHBpW1z6Lz3TtUXBt3LNTDuPALFDbYXoWksdhP74rNMnqpgRTZ
xk3TP5I4Mpm9chKGazUX5Wh33axgeDyCa0HREpJ/AJw1dLfenR7tJPt44U1R0z7K8qj/8go9Ftm2
vYmLk9H4vQzdB8kyw5uN+F3znex6Ro6mLinA6UMM7bAzdzO/MFNpFAM7Gx+MLQqRJK7VwJr78+NE
+MRTv7rOnvwCnyRkxqbnzys3PXPhlFNB1jMb1Vsu+E1DE9RJJIb2+mqmCag5P0xgsaG6kFpfH2K4
t1FRaP9rMGclbx2xekKnj6qjYbSk6szfV7DVMLR5uFv0YrOC5xsPlTK94n37RJ1wu9H0nomIYrtT
vhiKRcA57fdV1S+qxl8XCXaKejL8vPFw4h1hJG2Ff2C+zIf4TpnhjAZXuresPf3ErghFa3Py37cD
dCY1LCndw0bTwd3weQYQo37I/CG7CbRz2vtBKZOyWV4vPDLhNGis61u4A7blI3Byi0utR1jgMSzN
F0vsWhrwz2OEy2c6gLvE+h4FQyNKO0TMjCZkgou67SjCZYD1qcyBRQESWlS77IBNDAoZw/b9+xe6
DxW5sDEa/p6VxKiYyOclqq0QC92qLNhMVflP2BNtRwSYUdHAaUxxIXsYPiglq08Zn4tDRs2yYXAH
4dQItzdpjtQR5QI7nxMWlmPw8SRlzOzgY9QKakBZ8uq53oQFxUuFjFTR4xmNPMhwXatR2KgCY3EJ
RX3+6zhiEodu09uujW6RzO0dnY3lxvQ3ijrPqcaH7oW3J+feHGb6q3pj9J2r16TFAmWJgQcAJ2Mq
ApytIZSotFmv12c60qnAhr1eqaShVqdGQmD/nyBL6KcW8zAMcjHkMd1Pg5/WCrLIaVVO49Sgs0Uw
YCJyqn8Sv6JjLpeXzpz8Q5rgIvUPPuCCsQK1VVHq0Cj9kU4DQx9v0lnNSaXWdN7ZLJqFcL3Abgau
xWpy520aDgBKigajp5dHh0LxQVI+LK6fEwELDjxTaipkgglQ6L4OGhS79AeWRsb0/KkA1eHfKiLb
9v+WK+QBRg5AskVI1Ps6S/jT1MvgjUvFRd+sF/C8h8TkGBWpkS+cRkzdYu7xtb1dOSGuCeO6xBLv
3DaE1ShDeRUAOvEG54dEULgvuunWN2mStZugL/EdLYKWES68s+TAqK/IIDuFiOWucZvyldmTAMu9
3a4aCbRSflq40vi9/c3W8u26jB9Xwjvwo2M3FpIjP4aZVGI7aFxGVQKrC6uAgHH7TaOoP9e9FqTa
rrzujWLPwuuO5MjmWoWGOM8dGoL1F+0unPjO9JB5oQjbQcxMCff0VqoOaPdH0SKCqZl6L2IleFDc
tmB5cwZEHcyqA9GKz3vMmHUyb2bIDQ45lsiPqR+CyZxhi0s3gjK22s6ncj1gzJY95WYvEHX9d8Hz
Y8dzJPn2Px3R3ChRBpUOX/as6HMSp4GQNtPPUPrBcRGBOg3+i1nzbv2BtCtKhNCxsLw2bHnSIHsl
QCLSDxMI9iLQkWRiDvQXJOc+Q1VVZn1l/KrJlKQGCn7MXxK1Lu6k+w76cyPWBvTcdi3uVgp8+Ni+
dgbUcxEvVYJlfPNptUvcOOPxiEhMF76G18a8Gjm0W70lLabdNhn12ND6Z2Cjy+Ovrt9i2oFWbt5p
QmslKa/YaFli4ctSVHsiHx9DVSscpz7ag3jK6bxAU+hg3TAJfiKj4P+OMaMiT1/CmbM2Bffqt1TK
p+lHGu5NJkqOwb9MirHvYcjSFRhS/SL4xSiMtWqWnFdRbq7jkgy5gmmfcm/tPSsT1k4vZ+we4OjB
nLLG5V1sghwdMyr6517oxYzspKKjr4yYiBGqZlzJcb3x56EYgQrp9MsmPGM3eQfeHHiCm1ymELVk
VKN1HkVYmwBxHEHonQeU8xt1i8rromK/dVBKvNP2EeSSdPta8cLeyNwdI10h9hd43OenYuuzg8Lt
QLubJnvg6YIsE0ndQAPQr5uDcTQfrdItDqmTWxkdYbevybY3P9YyiZBuNETtay6p0wdvU79kYBCh
ZFuT+aMbZOEzbqfYax+KlYdcFSm+/8QKs4Ty6LzQkGRxNpelW1u7ABuVpTBGe30EJTuzhiNyohA6
WVb0pSD0G/td4/sDAcbJ7bXCej+LNf5ktAbsePzKVh+l5nfLPA4Bc3tACbPUKg1hDwSH6aflYy+k
7PgAkea3Hz+YwzWORkOEZVl0VJODgaB7Eazi/rtlvqCYQDF+8eznSWvlm6nfIep+wTUoSY7DORGt
de3OumeyQTcKFtJ37b1IuR4uxXQ3g+c2Ajvovsw0s0IeiUpOwnu0SFBlnJYqKSlCA9AmErlzx0R/
/Zy1AOT38lpwZFUGqhF1S6fZjf+68vIov1EHOEnndGfbskW3taaGhekDXqZ1EKTbv0xPr0HPWF8y
veYslEoVZ2QBVYOH7FQB6pH/lGs6dWeGqi4Ub17Hn8ZF3N80T6QtHvdeMSJEWWIkeY1aAZ4Ig0lR
l5uFco3gvrV8Ed187vqxwnFqhxpdQCUsP9F7sJd+fBP6g0TWMusWOoU2qVHq2od6vD2ar/+7w1KR
dY4Z5tbBT4LWLJclkzBc63eZj5b0NrwhSu4u040Puz4/P/5Gto/EVwA59QvhMK3nxNulp10+hXAv
Wsl88qv1IY6xnekcegkrusPgObxncjp2udlOhnJ0Fk9rfrpFj0O8fSmT7+XiHRnBUshBd7TASq0Y
ZAP6Nw+7iZJVZGqzjiZwsxQbhLpEcZj1JPlWsTfOQb13kJUkyYq4+yOM7EjRehSKfzeN68hbNFfW
SawIXGjniGzjFzLFSekqRqnWYkQdLnaMhEXMy436uQUZNS5lHcjh5VIpPEz6yXV23pbvHgPeD5X8
Q7ws6qy0eePOcPGF+kO5K1riqH2s0LYKKPCdssJKg8DpidKMKQ3FcdFZTiZpTxFroAWFe9DwdutC
mKZhBEQAaFzDXIJOslmgOZhcktgIup+vza7yNpdAZd1h+fP0a1EETHUirAN/ll5dHK+KYF2lXbeI
j8Ca8shKTwmRINsL91eYnyTiCAfXIZhXzASkdPzhGE91KGJsZFxSlrgLHyZvCGXwZbHaGxdhq4jK
Pir5zLpj/sgWebDSFinutl0vXOBHm/3EWK4AmxoqMnxP6hw5xS0NvcoqNNrpqmmOlAQenodJ1wXi
OAphLvpl63QNexS2xuSWU2YNChyzRk6NLf1ySlVjHrNIJC28ZPnowsX0IBOk8DcyM2z+QF7OHlv0
kVWplG5r9moGjLQ2lhrw2FMI1MylCFma0+N2ysap7kMpBrDZmnrkSOi2pXWODDSLt0uv3A09YCQi
XjuS4FKJSQ0reb61NeBoh4KvswmEkBGQSyaM17vaSkvIT2TpNLjSjvFXUTrdUqmmTPDNJeoxmOwJ
gy5OMCMvg3vB6RNKlOLxuR6zVcUSBcEJMvqp24yVyIX6beajmQxMGXxQRbKSykGzdKyb1lod/R/j
yldXaLRTRoEb4nsF1e06S/zOKJ4ZebWpQuCP6N4jbFVN612OuLuy3IHVnH1I2kqEkDndEE03FFJf
nbQKIuxglrhUII7RWRTYiwwTWfpQ25DJMjDT+ESOAWEF+1xlJSePtmPwW+s95NdUZD1vT7XRlQLM
Bls6RX70W4hKNgeflrSBgCLsm5dwU+oLozkIXvkcsmmaFBvtaE5IfeuA78LzpZB96OZDHOYjTfme
gS4PwF/q8Lpxth8A92ImPP1EHTp9JVF1S3zWzkZishxMImYzsQ813rthCWvJnZGU5GCae0NtIq51
Wsg/rZ5kRSweLqAZTvwQeOkXKzcON6MlK9meS9E+B+kSqjgOVMg64Gl/+aqXRuDtUDCGWyY2IgTs
r9IAhQBBJir0lW1HjZBzLqgLsGdiVkBHHftapx9CQ65wQHZaM4WyOzHqYjT3OWs/eUaXZACi8/ko
3dsQCT1i047rLZwyTVylajachpzS8sChhHRZTAJlcIPyVh8zbJsBlGF1wqVqiAPjpGkAta+YhZ9u
6xulkoX4BIqq5rvenIRxMJiW+qTniFISwXmTSG+H1wYw8FlZXh/1k85kqb4itL6R9YUKiTdKDuYO
Rp3b7hZ1G3ObFZL2+V++OzeoZqolWelgIqhVzo7oyd8+EV2dbfaqiLugWalztvfEKPSuT7gYUX0L
SAFt8+QOZriyjUtLVCzs7k+6mPeJseCEnwSBbzgPW7X+bq39SK7PFbHhQKNzeLonnzh0gjyfPAVe
3oKxO0wny8Gu9wp0OHBsd4Zzid2IcY8jmPeyYnva4YQk6rfSlof4l8L7ab3Md2+viH+c3IaeH96S
Rm6gGBQAHEZOnp1KlMHj2FN23och7OW0x6qWbtS62VrMU10myq/seh53ERCOmQX/ebmC1dpsOsBQ
5Q9RDb3LYFc2JgPmfyxIuoqwoqKP/ACQHA3Axa2747h6gAc7o+e4pjJC6kqnVqFblo+5+Ov/1v4j
VISZYCAzkpayhaMkFEJjIbB2rybouOxx3luM2wi9SJuT+MQrf56TaWOu4fcDFJBEQo28wtiPdTSf
n1Ysw6N/+ssPG5LBhLxZ4xWw8g/gKTPpno93shvRb/t0ECvVy/Be+5fD3o24SjaGSWwyUwf2zxeV
qlA7bQ7G00o16Yj8UnTIONikPYSLe7/tbVY5JUpBWaJSG6grpY/0fTfb/O7pAKH65LguQgtv8m4h
qzW11ikyPkytlob97zvZadYxnFUk3/IiMIJpDOXBZe4Dze1QwGJil+fs5tTuDIaxQYL3S9GOI27y
MHjGoIlw9PznekR161TBFO1pFmMKObRLGWEqMg7EO6LEwSJLJh/dd9cRJmuvyfXAdQbFFyDmLh7l
wbGqBMYJtPUuUlmS8D9niwDSbbFRNPwLwHKZXmd/cGBrY3RRaeO3gJNgcv4HEJZJHbq7oUkX3KR9
W3QjktA1cM0aJiWnVh7fiehdFPo3rlTBE9C6WDvPQMxGl75WTOzW6gNOMQgnJ3+9FrrdWtmjVI1e
qsRSPu8XvCKAfbu5uggI8YKchq6paeIrjJRZcfA403ISF/jR3Vx4q+9+0P7SfLstUnX1WH7yv3Co
RJhyspSe2eXqOmMq8XkuoHX2b+LztsrMbX6HfOIcJvp6jfJSukd7yWK92XtcRpM4M/xiP0eLv+X5
gsnoK23dWCHhjwhnIW/X+5DgNIDXXTPcUYTFeuRSCnydseWad99TrnX8uPMkp6vvULJeqmEhyPKU
JiBrQPaGv3+RVzRWLKjsKLwurm1LqdhvRwqLsziYB94paquKfzaOu83FJafQREbmF1qDzQTgD1jL
6wtF+JrhJZiXry0r8JUaWDRGcwIrMVg6QSlWEOM0NvYbseMBGSo17dZ/usWltSiMn4rU4oZRK74N
kjt7DPTtyWdWqeCHWAzBtZXGAzSdpWz9k85NHmQZ9J6pgXbi8yfWhvE+fycGFkjnnlLM2BD7EiHy
aXt+3KGrxs3lkyiPgqTibnPHs3qTka4ElySPsjCia72Z/m6Hwl7q5gjvCCdRoA8hGgDCPCwtsJBM
4LJTOl2cUwy6iCBw5AgeuKsF0Taccd0DyKN8iO2lfVPrxK0wAwZIok0HAGOc4hY19imSBb64GO3f
t5Z+CkHGuKzo42nWTngLMdBKMR/7bw8LvHpkpmF+6QgkgD+6bNHFcTYi2kYFzzUooxSfa3MTbKQ9
rpCjxt1aFM7ye5Ae/VYden3eM8LfKWwz+IOU13AvHXc6SwBR1rJhtBILBktn98Qidm8FtTVVN+p9
MEVtSF0QFk+txTRgt71wXIznTsBOzzVGNfUcJy+Bez5e45VyCF/zwdliIxCQkm2gl4HpMq+tzvaz
OHA3dpPixphhypsrfxnglyQ+w9cBDfPQLohVNqj7vrx0+qecrUTS/iHMoh9KdbumNYfOX23++ipH
6/x4PdKoxXZlTpQxoGqUTq6JimfK9dh+wOZpno4qjARrkNxdDV4ilADCednCynnFxgSVUR0APXFU
yiOnY4B9f8LSE3sD5wa0ScW2yb72MRUnw/dC5ha5/1kQRycCnf4HL9QvbTzmBYrrkLAiEpcn6mLB
uxqtMwCq6Uu/rewhtJ0M0eg7W5ByV5zrQE92Jk93s+u+OrJFRr+Rxwsn/PeQZiKMEWgssa5k4Iak
gEpcupgaMUdkl8YEzDF+/3XEul5i21K/RkDkHkKZ8YOQER6YwyqZzUbN4/gObmsnzchLHWTs5+c3
QaYXFZprPso7Cb3cyui7uuN3Ua2Jyqao+R2r6qumsdJYPr7hjyCQeSyliJmjktET/czrW9uvjCmt
kaZUxhCXa+yBM80PfVLOZo0qptI2G52LXn+AoDrSIWbqgcZlV/2Hfh32WhJfSUJEZDg8Snv2dOZj
UdXbQf6d9UmneJmfhEdRbw3GzTICMJNwrX0RFY2TMU11L4jKsP/9Wcv3TeUDtHqOws5ftOSuhhf6
vTSVudhuACD4s6ySzR9iVKQcQrKXPYA5Lt6S4uUnImlhE9R84Djt6Hjc9mwjHMroHxPWIZQKzAns
UzQB7plMzf/FcBYvDhuouDbaEgJjHgWeYaCBHhi0SHfjI8LXzr7n/c3ZrBbm7Y3MncQLfgFz5Eaq
gSJqjGkYarHzB8EZy8285tc0Xh+z/HnncL8lTjKP8+Hyos/s2y8Q8tZk9HSlnd+of+3T9xQvaCt5
i8/lIWbsvQuvfrpF/+DqVSwLCq5c4fSCaipocPBHeC9HiAWFOo5wSy2Bu1KcDDTJHW4iNWzUTkzg
zgqjU3zTItWgGZbBwLr5FgF6+48tSctqlFvFENOO8KukPtH/cx1N5iAj8s6+v5LbNr/I9IDKc65q
lcjku9Z9Q9gVp7D/kO5kmgW/XxXjkv8dnqXsUuORkdRi/193ujN6o5jCwrTjVy8GdtrvmwqaS6i/
nLB5MX6DACT6hAQSFmUDyR9TSatM2OvPSSV7xA++QiYnvocQxD0O3PWgk18xv2k4/vDJeUlex3Yo
v7ySjb3BtkDylKzxmHnsyxiuImrf85C329nFMrbd3luZ1lplhuYw6qGwnzY1ped93rSK3OzUSvag
dSy3ciinSAG4Yo0bZGjWGilXzU42c9cg9S6jkCI6MoElwrVGkXG5COIfXIyh+tDN8CwW5TlwZicc
oRpcaTXTsn7QtkqRxuvS00Qp6XoT1XE9C4n6LqWjJEbpoQSjQh2SRtaQ/UzVdQ6wrn93F6Fs7ybo
zNNgXsb1dLc6Iv4AcGrp6UtPYcoJV0mEHzR2muGPanm3y9nH8PZs0OvQXNfacAFh9fIylOa1Bfy7
6aUfSEF9YiDajYnfKcFMTOI5z+32/Vpg1TmKNULPqlhbCLT+OxZX+QYV4xfkTyTXVyduJEyeHxdA
qdpoOfAmkHDZsnZbPg/QkD2AWTGkWLJXwqWqaAJKUl8F4/bN7owKWEPJJK+H+JcrXZE1sY7uwmfO
VKtYFADS3xZE6BMpFimm6EgO+pmt45x/xXD9JsiDalBVBRIcbOaYOzhQtNNbjm5wHgF4/b13n1j0
EdcjMRlfHkWLfQfI5w8a46XMVrFSqVp6LRldgMs36rc5IY3LopzJiYdEYSHxMhSzUZcnlA7O8lbq
AnbIhBuQw0TRrTFqPGda+uWuyWFSCUFEvFZygZdlSGVRkczbBTQ2msE9PPCi/rUQpL5ZL3zCal4k
NrfaG2uDSOrxtMsfpxwsYVDM4ZjoMghQI8jixV7W0KrwKrelJsBlU1+R1fmsXYyUahCBTS+3o0RI
gng+iBZM+cDiLCKzMIwnsCMJ7xaqun0ywIAB0dzqLYl3f1hLWDrdoFqbGUWE1C6SpVxmkilQ1uFc
7qAWIgNeE8vcJxQA66D5nvUy1CrRIq21wG84Qja7ETiQNqMR0uWABDBQvSmz5nt2uK5eaz9Xx2gH
+GFJdutXY8f3U7sxG+J1Okh0ziiD8t4dwsIOJ1kiB9zVEQsS7M+KHy+YjVGQAyYHWgSuoY8EdfTU
WjNdiJBeZqq4QlyA5A1TCxLKDSvVdaR+UObRIkCBlVarVgYw3i/NW/V0oPT/2UeSM53CCn9bgS0c
Dz5Twn9AczXcMlkHraRGAssZ+SrJgpeiyOODSoW33HFI6tnOsUdvdBZMakLvH2tNgOhP1DmeRfGS
zO+qTEyVG/wDuqC+EuA2k2DMsfer7VpZHTCbVxYZ3vEQjxPdpl2UjEJ9Syxuo6U168c1Nl1in0xl
35m5CSYitTSjnXDCsB46z/uMH2fsHM+W7PEPhxUJYtrrYrerA/ew74IUsblbKmdgBImJ9Wfcmlgj
RBvpQIQNWQW4DpWi5uPTsCadQR2/j97DtdOLAE/fz583RdH2JJp/WgnTyhs9bx0kNawURtWtY9QB
rs81381YkW8QQ8PKZ2g+pBK1ZXrJZ96oHjONWMrXDcLY4C6FMsuer3JZxwyE3i/xVTcwLbvnMoTe
wijTFrj1HWbOIgv2vXq9LglXbfJH2iksUKHDjUxz+YOiQXvSfOiFAVsdEgwS6SldZ623jxrK9jT0
dgsH2NbXR/lQe6C7eIJ71m3qjeJv3LqU9Xe9ZPgHdrZ+ZVPWri5GHZujkRUC7UUp50IU1CfUg9xZ
qkUp/UA/rqEW5o71cAgMDX8ObhniQXhcnBTi1QDAyej3uCv0q4+Xgt6SoHdHbziQTs7c+E2zt2eV
KrJ5ASe0wtiqjuJ28Qd32JT62zr0VIZdSRgZkKk0JrkwosLMBaVRyU7FlcRZNPRZLBSTBAqobDHv
xwCF5rhJSKlfZA5uVwL2VOCwDOCVk4W1Ws1fhPt6ORxleaESlTmpgZyDvWtv9rUJxf4L6gJDyjeE
rXx/uVTzdzf4aI1HRhL2h3LOgg2s4JcN1if4222k0zXhp6wDUjPBCk3N3GHdHPUqf9p9EMZc0nQ9
A3b4yUaI2Vx6b/R1mY16KcZ34x4aGsRu4F+f5b/euPTFcJYuMvAbZBDBgq9QCooLCGWQQ2a9wXcm
i6bQ1Rtu7vSOA98qS07RbrQmBCQo+geqR1jejMS0b5dI80tGwisWQx76W5EotXl3YqrcxyxQz398
duuAwllUwkRMbukQ5QAE7fPVOTIfdSwVfAZ3KkR8kbiijn1BvSGUZTxadPSUs+OCcHHRiaBZPiGN
r16JuCtu88e5wGL4GPjH1BOv8QgVip6IeuH0KBCfimetRSFjOpNy+7j1BzkbrXfSTdjIU3h7/nJE
OgNrF7vL2AWg0RSqJub7l6kS/A5fjS2+I3ptGG9mB7A8pm0Is1s+d7QWQOcbnq/YVNGkdGPNSd9O
f28FQEmpOTiP0QjBJ0SurNOmNvi07FazPGiOAPAHK8j6Gv3nuDgk6I5hsNtlLTa4hL+QPjexMVkU
Dqdj/Om0/s6vj9hZhLUB6qizsmC5Na2KGjZAivOreOO3M7kf92lGeSHbTYIzQkvfd8SOZaC39vkI
Ltd171MDyXN6hNSPeZiyifRQ/fXKJqpVlXbC93q0VrsKAcmRjqi5IsJs50CTvVo2ImDtEhrWAHgo
21tlRST/10MCr91M51h4lM3LSa0cxcInBsRwV76NvvgpjN3T4GEmR/phcbSiuvLSfGYtisDn2Ei4
oFM1Uh97Fs6Z6y+HzJ3U+9dD1S4E8NHRmR9DlX2P7J7LQ2uP6k0J+g2/lFiYxRRhui8iRvosO7VO
g9upEhGwDe2oBUk1qrNhIONjgyjiDIqYiG1ACvS/m4iWfiv2+Sr+HZW2Q0BGviryUlVWlRdGLViS
ZmV2ZPw1Z7w5ouidGSBBlWFgHpvfME0RtwJX+w2Lli1izlqMh52c6CUW7juCYo4hR7TONsnFwwpT
8DUn5WWKpKFO502mEuXb3NedWHHsjkvpl1eqxRutdpE210vXB6/DdljpLUUaQj5x8fFt4lXonG/k
mtQ8zegAm1xJ6u63IA0rwk4eOObjMZPvryq1wUmkhxZ3aSG4MUzKTC0U6ADN9vQ9qQM4RszLzyL/
+09YyfHw/y9EG/jEnTsGjkrv54CrB1+zZCiQhCD23Wk9wZLiDKquZzMGGW1Vn5w/N5bit3HBK66k
yKEw3cN8rljN/jUuNF/0q9PhEEVJ4m3qtG/NVjJqAWVH1JRHiJmqY9oNrPtFiYXqhfVq0xVguuLM
V+5rvVUpw+tn5F8en1aYZ4/o+wwd0vE6O8CUr+Ty09AAJUrzhumcXOlwlQAC4Ej/OwGkpCGK4rF6
MHLWTsvRr//rKtL88WWdwoDQaNmrEhl/bfuAcUMK8fihjCFELpby5oehLzZlN/Yx69hhCjDnS+R7
N0We6Cn39pu4vyjPCPw0JT3x82T8imTGt78hrXUfbU6fYEbRL8B4XVg6ZcDmLs+lOU5NXuoTIdaL
x1s8taQrkOWLvTf9kQ5cmq35fWXQ34oLlEyCGZA7mImtshHxwaYVubKNEU5Kvt/bqBX9JXNsSN6T
D2gpBmvrPj7ufvu7v3KZlIejhhQdqa5Vgn45iHU+u/BjWJStBULYBrLWhA9mTXrsAyatJ1xIHt5W
X9vmd14/hBDP1khKdu0Yq2dOMcfkOD/W2JvUxLWS9pOqIanS0AHzxDFXXUappdqZusDp/CY1/oTt
zVRyRVFHqh2coqS2XhJHiPcBTQ8MnLlLKpt4u3IXLvl2ATKj01lNHQ5lH4sysxICjG8JSnXNtBGW
GfqXEymCdIQktLW3yiVAh7Zvf9JnBR9/u1Zxe/PaTRic+tqTNKOJf+gLetAo1CeIgk0a0s1/XjsR
kgb6okIqcxctPu0W2u8umvGUp+O4r9/6semmmIaC+IVYINPyYxSJ6QMGuG1WaJ5LaBA1SoFfSNw0
Sr2Nvx05/RFBvD2oFF0WeJ2FJayJ/z04TazBYAPGw/u3vU2v58FufhnYUdUBsa38PcYVxcGxUfhN
l1q7YwG/+zm1ydfdiDtBS5a4O96be4+8p0EF8M0DXdHygtIHOOxdDZF8ah8NExxynTY85heudAdL
8vQDqYtadnTVxKylOi40I+39KAU68UweB0rP2BsqeRBQI5xzB0BYiudM2819ROTqjEgwcwXMNYaW
PvwvqrwgeiQuVX/FQMLRzqxNtsC90oiOUe0TgM3pyYEB7GTPPQQm5+d4owA8ktpWQHIF3MK7w/0C
6HV2lcFChRa1W4dduj9unNlICzkLjr0XjHnBw9ptezuKZB7iBr9GN89OKEtrbkVm4I4O495gRcsb
7F0kato27bj+HojPell4mrs35brW0sy4nBMXXlUmiZJC2/m5ivAwnXMl+iPxEKAUFBYMjFM+h46j
y+pMhUdOV5lHehgPrwC3GQRf1DMt/3FxbSHyqVAktSzOfkYD+F5nr5PCAarYLZmH8dLs3onRg3KV
F2QG4/ERnsGpY3xOtjiCQGU5pGLykZv3N9So2ipIoPgd1SG0VKUo7iMaBNNNjcrebIWF/J/q+RlH
+dRauoXIsuFrT/tepxrLyH5ytYlnUsezfb+pH463nPLBTE0p2Kw9MAyT/IQkt3c3CzpWrsuhKKuF
t+aSOqKcA2Fsz4nn8Xb6A281Fv/sjh67gMo9jjujchrfWtY5cqj4q7sYCXayVdSY3xIhghSl9/cP
oaKconnYNo7a011RpFcxJmmXqmT0vpFm5Tr+SFWgneXcligkvbY9bhXzA8YEBJZ6xn8mZgHH9Z+r
P+W/qEREL+wqB6eDeNxlgm1ZPSazSx0kpvzNtvkVSnlXoPgGgmFrPhalhIXA0K3hFD7gEb4oyaCS
rpumTKYryWcy8vcaSUjPer1fBYjW97g8Jwtuui92Zwhn5XQYjg11t69OHMFW2CNbjFRtvajy/09z
SniVw1JmfXMEYpgpnYLMT8KZIMb6iXFcQUwU2tTY52lmXTnpZifcO9yBAoRNzeceXfxlXRoitums
Ure3AOzyhLslRLsemGZMWfKzZ3SSVT6zmbF/J1K4ckoLwhxw5l8xLtAp6vzxae/wFftazkUck6ib
ZvJBSvfG7N9ZncmSj/juaIH9SaQgEKg/Lze+wpHFYzxGwUSxVHdUVmL1ngD0L+GlRqldFbKuICET
AhOk/fBq+THNf2CeOhHylOqCKbBEpr9UnwPcJJcwYIB051u2LV8ykNl5CV4ACv7gZ+QYiwzJHdxG
JTcyS4SNJbcakjIe6kdnYhvtEUh+G4GxkN08pKIaJ76Qd7SI91wBPRhaW0Tw88oI+HsG/DRKjwm2
/eemAVAvhBSDkDzbp0SG2T+kkKkbXG0utI95RLBkrCK8zYcm6ihrnZkRIGJfStWfRBW5ptnzm3ch
D71BMxGESmX6w2FS5qDHVkla5uXQ9yMtNfjmuHzNnfW/R6lZfdZI13FrIoRrYduLE0fHNL/MogbH
LcfpgaK/LQSkslgirR5TJKnP6gUrGCgm8kfuBPJo6oGBUyFF68TbZL8Tq/o1WkWjV8OqJWOSlVZp
fRmkWtdD2pwpo0YhkDxsbVtoZA33pkyHjQuh2CDfeg0ktJhF9692oiWA0/Y2/5KmKFszJarzLNLQ
eX4KJwoAwKp9bYclR7Ryh6FPkoXDD+HeiUXXGwC38b/UFnyMiXIUcAfAUKq65q3AbbPh2QBqRN49
JM6tqTLNEcuo/5tWivmCeX9quNAt0G7lG9/ca68lDP0zcYUWDqjW5UQ1qbqC+qmjyRYVgU1r+7gG
JqKbrRlHZor9tuXtbL3+NACVS6qrgdt+Fg6g2PmDgzpCocfjJwP+m5CZZIYzVEfhbAzQHLhsiLbs
F9TPLQ0/zsBrwlhS4i7b7xiD/9ZUd5Pu+43DNfCzecxeOyeNh83tO2RSmHNIoFNvwEqu1lZEMFGH
1VKrmfmNmrH7bss7ZeXOXD3rSh1rv5X4BcK2dwuwmwEnOZOQYhu05DFHlOqq5QWIzms1Msto/bUZ
HdUf+d5wOrJu0Ot4VZiB/Qgq73biD9T4xE/N1rvftCpNA7MjCkvlaVhd/s6bKJefxfQ92DW/efK+
fbuOcWJ3VPNv1LrrSJ1+CrlJ9WPsmgoWKj82BG5Z/0WioKk3Vneaz/reAZNbHcj+xkICAXQFSrCK
8chnlZyDSv4kvr1Toh4WQ9YLVIEsr9pScR3yvjjfBuy17ntvu3W2WW7HE48cDMSRvUuT7D5fAxy3
xmTjlL75zP1/JT8s8szyPGt1kLFGzk1mPU9EFqca97J+iLQhZwlcnDOXMzMkzWpvQu0NFavQnP5Z
G1lJ9Fas9ENtyREUws9Jx5tr3R2erqMxN4IsWfFO3uYScx0J21riyldPCGzS529ppxCiF2DCZD0L
C8watDilXLqOO27iiz3TuCaByGNU4zx1bXAochSydvYerIeOlLRsXNxQndUXDvPPB9qY+xxbQ3g7
p4Gku0i4f7/A9l47lbzlWUZYLAWpnkKTdiwwLnL7qWBcfvTBIq1HnfwYIGe9dAQPhhCubMLL92g7
MdtYDoS5AUcpTbYPtnFlcy+3hhQku174ICE17e+Kr+diDsoe7g+NbPNZMIAN45kPN41lrdAWZ2Ze
o4fTAQ9HZjOEB4vu2vwRcAYlp/z9Yo5aidijLKTiVJwRmUgnilLZp2p+VO+amB+OYUPxJyIDkF2R
4a/rplKM3uVce3xL1PH6jGSWglK9Hq5oI/t9YPiSOTFIA8brDQHSQ2bS1wC6feZkA84a99ToBpUZ
4qN2r+PPu6JY+qG9gbDA35oj/Q8UN7aLmDCwsdND8Xh8oR9unwNhJlVn7PQb91/+T0j07uCrcFgm
Duupg51F6IvJ56NA9HKt0sVMfonLNFE1C3yJC+6wmE8l8gulnAH7sO8C2QsQFABNt3WtlBHAPj/q
xvx1XO3CJ4BK6KePk0u6uV7ArflwNEaT9QA3QLhlj5RogxpfmCleZpLCgUVjv8rVtCdCwYXK5VkP
ibySsV0Fiab0Jv28XfZ7z2oXpxmGVFFQ/p4cyEcknPvhdeOjcvI3LFK1mMBSx3GpYFUCSPU43ZBS
U8Nb1cV5ZYd9CbO36gBZk5VBLL/xo1ujeathglbw2DyS1C0lA4YpJIKVL/9GKraDPPclRdl0k1bU
7/iboNaXw/pvagl942k9Nk2mrs0dXVI6R91ZcBTnP20uhj4n2ktQnmV9AAMZpiC/eseX2TTF+Rm2
UL2FfNpVl/hz1ZGe74bdW96ojeBBeQSqgrfxdxPaifRneeq9pcRgJjURCrGYxgXBMd5hEWDb1gyh
KrWEAXRk8Ngc7Rvvqr+8UEziyP5PM0AT8mDfqU+dNgnhhNQNQwjodKpN0+hy17GM70G8Iavzn5g2
yXbmL2Jby03gdlrG/NPlz0KczCC8jaPWmzpQhn/ZQe0jPHjd9hovVS6/Aq0VZhBqwXSbRGr7uE5b
bbFh0homWYfaqf+Cx4u+kggTomMFJLbKjIS4NAEEWZpoHldgbOinD5b4NCWdyoftcBuIwjBuG9oC
e/OSpl6GTvYkZbPt8w+J4aFReLfnXPtdJo3sw/ssO4kS34cmWIn2IhkVBSWps/aMhMpYVAxMTCgJ
YdcLML66S3hBW+K4/xLR9ov/7ID+4cePIoA2UzoJE3Ic4NDCsSXBDgzOK7K+aP6GdWMzCJzEgMUM
1FTiDpZK9Sm2E1NFpzNOgbaQGpmEHyhTv7GPNFGPzOcw2bEx6jaQO8c+71jTANuOjm+MZ0rFlTTo
zE7Tj5PSNawy9UPwckf2QjqMKxIJIoAPOF0d4AAUQ6jdNDyzwIldiiBIKecZ/+1n5Dph6VzPea7b
d2z2cbXyTeNOEi5pGyYinMuQyJoDkzucfvDU4DkXxzgOuOLBf7VpPh69HL/P4Tcu17br8Ofd5cZm
bm8ylJmRoNa/2fwGNoEmnddlBUZei8E8T31PurmcPi7wFMLS2LFBG4J9ZAIMvDiVc4oRj6LZEfNy
jBF+BmrWcrc/RgZQ7bbREkQOORAa+h8EsYmy/wHzZlZx6m+TJPI9TNP4wTpSI4H3MFC8zK5vAbOh
rOv6JhlVpe0SWqUvrrg4hPVL6o2CPz54fPp8SMPtM0ULZdWRM2RoljLizf6CmHnPZS8dElFMy3Z5
zoKmKqcBc4iXFnI5U1JPzOQaLFpx2y0+bjQsMBnzJvPcR5L+uMCxxjmn+imZCee77NM0bVkG3NqS
jvLbeY31p8wKmzh4fWMhKr0KFVYOHqc0k7pjTeX03tDZ5ylSXagSWJ/T2iEo3iX6QGg0pKuyr37A
pWUoWHxmUAVVcmUZWD2RsDMmgmWvZiAitMHX9GTlsz37K2UhQ/DMOYx0FUyGbzn4yNDg1SGw8H1S
+ygKsVtnHzue7pppWHG/9jXwsHSUCwJfPM8Kdn1zOvVB0Dm0PY62ORK8LUAhgDZ3UhSCfKOHi3UI
wNfPB6mpaPnhSX9h1cGCjoeiEDy1m10e84XLtJY8/BY6H2SqTxGoQcBNuFv09B1D4lomKz2S/TYC
dmWEMODWxu1zGfOs7L8UVSDI20JvkYc5Mu7H0j1m/dHeDKndnAQ5Y+cgldTuwZPD0MRqb3mCyryw
4vDmt01QqBLxn/Iyhn56wMmfImPzvg2/5VtKUcyZh+hCYIIYfItmnUixU5wWB541WwZ3ghiC7nhF
AEppMSoGiEcxaft9kTovvfheE+AnRI/MbMMdjOh9ljmNqfgv7i/Xzi51+8/jDJL1OFW21e+LWeH8
fyS0dYb2OnWv1bWsS/P8wY2t9TheB4Nd0ctetktryqTYS2AqlZGArXi3hftFXdP3TO5+RzxlBfqq
wSjLcc6jdr/kbehW7bZfo9CYoFKo5w8s7ch/UPfe0s1W5P2VN2rFXujFfhGYhzfk8AdrA6/aax6+
fJmypkjG4p2VlGkxT3GBeZZ0mcHAYrcjc1MloCazM93NSlnqvnn4r+CLwZ/QIEVsome9XYGNgQRO
O4DW2TXALq9/vf5n3C7CtaMN9hr+fjhuKv8ttcfAFyIkaZEhCQrebkzRMABbkY258GOuzojm76Ze
afMe5QtS8EqY5Bg21yAfam4E/k4QIEnGZABsQXLmI6K+6DkaMs30lgHjoUQWKePaFuAqjaMfhL5o
rNMfxxCo7tIaoXTvCktJ/OwiWZ9g2xZGEXFjR8AmFUrWV6DC4gzLTByXRK0hOUOd2e/r8ZqRUxKs
Kr1Ieo9PoHaGkwPNIo2u2Fi/8W6wZEHsXSPCzFFhe5AYsItsSX4+WemUJD3vORAgjr5XEd+DYWys
xUHDqlJeSHkwqzNnRHO85uehRInKF+6xvJLucf/iLQ0tlFM3MD1uMzVPcbDS81YkWIyy0xtF/euB
UQkBEpWz3QF1yOvqcJRWEKEEyJZxlajyQQNNtgyMdb+QEtIVfCFpZ/KurCsKN6DnmeMbf7uG10UA
ZcFicuYC3rrI6PwRXIOr4MjkT8GSDHoUpz438OkOVaxd8pSGR5L4JLkPJE+xP/2YMzYB2TFD+1tt
WkRiosqlhmHxaCzPyh5ylP7JyU/0cwoKwLIclWvEHIuoiY0uwNJc185EdRKfU94Re69b1KO5PDIz
P0f3tJo014nMD9gwA0NLC6Dl97jp8sy27a8MDcdZv5yI4mmHdZnCPGMbnd3zrT2aGsuhai95bSbV
5iRM+88IyhsdkWwqvq0BNd1vdxT9BcATRH8qsmg34tXJ9Ya9wABRdSBUhnhSeQHya/dqbppfDxQ2
rej9JX2gzbeqyZo1ui6f+hoHSXTruy0QWKaumlYz5g9FgvWDREBe0lr/F8edbfHeimpiJiIZWPmI
06XYmWkxWQhFylbIqqjlkFQGyA7H4zlNC3kkNb2FsEuNuvs3L+46PGjWC1l4HBQexY+M3k8yJTUd
PG0NIUwuhzUg+OpJSVtEf/oAFULCigR8Nwli48aOnnkpsolx1d2N9U39qNgTZJwoigoaHRJ4Mn7b
pTBhLa6inBZ4H4Hdy1hLtnB2UEbcg+hRl3uWCBUXyJX3yyBAvqDLebkn8kA6JoSOV93QcPz4TxQk
lpfjiOxsKMR56LROLD0ACEUJWFB93PdTcC4tx14S3XQbdNmDKD77tpJLf6DnfmtPWBk30/+sHup7
0Qv16QGoJgOp8Ven4p1hdXFSbWQON9Ygixixf55JymzuYFWCTwDURCn0nFDdjGTWY0lJgHNid1ix
KkfpDlQvhDM1YEYbCeCLLs56pyEzaNNUo+o2Gcjwa2pC2deHIFKw7cqbk+mIQ8Ew2J8ksM9FNVzC
/9jpEiG/6DmgFYknARDLEh5u8E9HyUOde+YSL3svRcewXVV2lFVBFrmnj7RoPDIEpmqDmK2ZhnJR
dDbncYBQVZZurVQR2ieMuH14LG5yyS+PVKKW1f+9kTt0JVA6n47j2aYRdQNq3b3nO6L9hjrT8Aba
jHbEFIIqvDom5i2/GwkBKFxbSNDxuKnPm6ggJTSEzX1xFtlS4G6eX7fvBhPKBpFNQwwgEEOxQwo7
WsO3UIL29i+QQwNrru2ZMsGCr5hW6haSZLOwuqgcSmVMXXvLDmViHKwbkR9uphRgiehZVoFnHskC
Ci1RErnovB7K+tANWewKyWAa8hgPqSUTqCiam7NPxEz0R0KdhQRG7mWdhUQ4Xx6TvIpMDbqdS+DS
ucsdPDull16TT5dxo8i577sCfiZEFd/gQqSHU9+1RkFyCFQqRQ/TpLnTXeEcVoh1X3JqWN6hSWvO
O9cis8746OhL8+5hMmgYEhYA4rIDxNoyGyEoOU5gpb9Q+tzrxGSz943ol7xngNh8Z9bU8FbKQSwu
7lbrUJtZkNFUvOmfXy3OoANvSFpWwvquLhG+mIoogFljTgM1PZFs8+bIy4JWbeo/C30ChjLWzJxs
Ze+JfLilHyPD4Z9/A6uyC6mXbnWCyR2qu+z2zA0o2ngekzzOz2xB7SfW0UhBpTHwTQ//LtSPcyqZ
Ll5d/vaatIs1Pbxz7UVw6R+9xGpyLBLSOstTfHZRotOjFPZrgnrSNyLLP0TrmMQcbEzzh9GJCL8O
kmWXetu/QduWdT8Yvl5t6jcToxbYUd08iNdoKsgSEFk1g7iRpAaWg8T0Ozurr6QJwa+5+eN3VP51
Y9oS86DZ78Chu7pVEiylf3MSqkk8uvJy9hyQQwFGLxYfb6moZ8IZTPYoqlsavhKqlu622sb7+ZQt
o7QJwDe1FxK6cYI35pCJVJv4jCF7m42+vbnA9SP6v6O7ZKtImWwRRepuK29f2aF5CtdtcHfkayt3
naHwgKlZohKXMDRHNd0FmW+862gLDq7uF5CPwFIXjVqBc4So2Tc5CpWnuCTgOy3j11/YpHaQA2yO
s/kfw45xCmfqXhhIFKbCx9bHR7LA++Lfq2Vl9bc8Qki4FeNqpbTjqpc4mxiF+WtmC2jh2+7lKt69
Ovg/eTw7AqZFBPieh+ioC6vnDXU3KUgWkCe1rvyl30FCPiVkWHYj6zrVP9U4AoJZA5jwOFhNSMoo
T3VyhLOSPMUS8jjweayzEYMxVCRsbH+4xmfs8UhCQDUrw94jqzSBbC6TeNtSaRKbisjXgMIzy1DT
i4qMSJh1jXzLtQOfXdGCpICG4G/PvBcjXR36fo5vNMUNNjmu92MdXrlcnIjiggCh4h5un3OuT7oj
3IUbLFCArDbD1CzjXFzOTvOSZeus8poXC/+Ibfl2bQ2iQBa+bn4xkIvHLhisllthHT4JH5EVaUcW
xR9uGWN2o8iRUBRJV9IumSERDgvansrgvVoqqq0KZMyRjsr4gedkZav7cOBq4wCcI7jW/cCP9rLU
SJBHPHlr8z1yJVObD0G/w8tmhwp6OIb/ckKVwjOqVedhteETUaJ3HzKubm4k5e+xwSodSPKJhH8a
SS3YUKCkjvcYQXAYp9Zacq4DPT+2+oNWFvOias7/9BawFJYVBiGmBUrfBfBTve7C24Y0McjRb9z1
CXzJsckNZiZTYT3HZQ6XBBk4aJwkJgfXkUMQZkau6JfL0W/7ehtaDxsJHvEX+ZMD+Hag1tJ0yLlc
ltexUQ5wE5aSCoTEMtOZlzWxiwpZUuCveVuuq+Dy6edaasIEAJgELjYurNGQhqFQYqyP9XBk/jMI
PplMhNX1xFaOEAXelSobK9IVcP6otC9T6II4muUOYHwln6Go1rltmnQzHOV27zVsJuTTQn+Qca9N
JxAOhtAZTCK/J798AXKpIvULZLv3mEFO1qWQfVwtfdFCFiWBmuRDbwRVdVuwKR4q8yAdGM93HpfF
X4pfogc6D0h6HJCXKfzohBQ/SydNsaI14j/R1lQHXeg5h/Qxvm0Yx++JVEFbSK5ieeJW7rFz4fBT
79M7lcMgyDO7sUujahkRBJhx0SIwKTIXIxUW5O8cG1W6mHFasVSQat8sZOxi+3R/fsEJ4CcBOaf+
lY3WYbYlLR1AupbmVIHNrhROCDQQ2NxjdTWm3oaMR9bhi5QVe2D7X7ZMHTGNVMe11jWyQVqRH8sR
DevIyMtnZDoQldnTkPa38ECTaLRPI79ugib1uAm7vOviI9xpeP+Zx4fK5tM0rSU6cocpCBPrny2g
LwyAerIZZE83/ns3nygAihGTMhynTUGFt+SJNCarFdy2ExTfThhjl90U1VcFu9yY2hrUnAfMAYv6
3vWuyPs1Mg8mFS1jg/2zcGMZRVekyuzBQSbLMNxPuIDJId0pKx+XWJI5oTTX6DIzGheIm9lf8WuE
f33l6kNyTAmSxMmYHbNYHm/JxxDu9M0XYxLug1Rfj9rFPvgcqlxHtGGficTMwIcXZe3rwp2deDoY
afBG4H0z06NqUZQy6zc9DWIMNPz5ASJ6DGOazkBOc4dAheVC7+iojgciGxEYjJ8o4L40WZs0U+6H
h4YylzxHxuDDPZktMmKs5pxx0RY7cbrJwrYcJ53s+7mTUOkJWPP59zoCNs5Z6p/0KCfciqrGoh2n
TZfipcgc0BViLraWxBKHsShrtbk4YU6MJ+E6rDaH3Ls3cfV8n/Q0QF7NfjNutIuzYPLCoIoZ6RMz
OBqe1AosVk+PYhLsTGRHB/8e70ellcfALsSPjLtYpXEZcrYAFcKWXHd+rqXEM7PWk6sNP/PoIHX1
v2ob/DNtRHwo9AU0/EOJlu7uJ2+29hhNkxLWDTLQjLB3tQdr6OG4Mk15f3ffG4cvcb2HSPyjl1uL
yjMb2DD9FdaAbMEBaKryUe4uFfSOWLgFZ71dKqGbOKtH8hIWDGvt555yJP3BAmY6Fyq9mUSDnImo
bPEhk616qopKJazTLGdEGxQn0A1GetiiwNKmt3ilQ8L4PpEgckpfPd2qev4zXdgktNiukklHm4nL
E3FRxMQcuZovBdmgXVCjFZtSHRhfDkEse4bnVU3eLfVA2YC+E1h1fx1pE3P0On7vxegcOMdMaab5
eaJsH7x8LjXNrCxaTXLDjUaFLkEr0KrUizr9eRxSEAL6asPTMaMbZEZ6lOdj6eT/ylrzEfRX7FpJ
UvD9JxdzkIvn94Lscsk7m90L0P/AYzqj5zpeEvI9l2iwcac+dDt+uR35C+5XmOdhp7yCGNIedoHt
FqVRv2PjQW6bObOFGKVpcUJ5vmFKGlAmeSN2/FIF7CSHQKx/Jd0ib/c8e4NuQhwUgCP3xnwMKmeL
c62eVndwWjHdGnk5DNj8wBHUXp8+HrcLSGeIlSD8t6m875mvJhU5rLx7OguKZ02KS68gpmRCh/c3
ihunpTtgGll9tx+1o/rnLmZbLl3l+NdZfYGFJS2o4cscFIJOG4qVv9Ht9pf6MdwzJT5Dx7IufJBO
8AX+kLhK0V5Uuj8wPOuf+bbUXb314XspLCk1Z14XQRebfnC8rI4wgVQdEZqZ+fSoXNsH0Br6voGv
W6fwma6yOLiQh85Eppy1kJ++sKPD9/7earYKUs1w8YmrVGyW4/YsC/KDc045479ruKIOoSLRTTgW
pQ+0K8VuxagTFwd/WYy0834tyT/NtCP8UxQPVxAdgfog4plnIbKS7IiekcHsXnNnMnkKC7cKdxF0
3hZs6jz3R1eOzvYFBeYPbCiX4fQcnkx/RFcoVHXjjUlxYhWHO3TNv6v+B+a66lKpNhVvIQLKuSo4
OOdZ9Ytn3f6qqTAyZsvdacWfdcItF+jyQ9Yx7cKdiqSFwG3EAuuFrcjs8mtpUyGAhz7FDQfmsUoM
rcl3tyCB7RzBnotCLjZnovVLnVC3eVTqGm/owhnIbonOvdRtO5ekmjac+ZgpOqbRjf0Jfh8CkZ4i
ALiS7c8qx6TgAQ8onV2iB1/ceBoYLKoKAXEjFshMnGW++FbWgr3qKj2y8bHzDPfV1i3Pozke3Y9M
OC2RutCmchjJeEFtoSqdIpBVcSZcLJtJU5reLLgolold188A8/jGn8eD9SM++PxNT3+51xqWH1eE
2InCPt02vaZwhcIpnjWyEvobOjLsHz45uf2vdpjAfnmd1DMIYjWYnxZrQZo6X8gkHSBB+JZRXVNn
fEw/bq0+Ke2e1Xt+UAuxQYS53ipbg5O22bmA2Z9FNVbUs+F3lwuhWaKeNvAhFh3aRZShLFjCcr92
Wm2u9bqc826OoMPg7HYthY4/QCkAGcgpPC2lcRuPaOc71UxdS92oIHqVfOqg6GRT2/GavFIAYkQH
WaJ+JSvzKRbKR1hn1gHlxuXtv2quyeZMy5gu81w/6oPJ9ymaUZszg33bGLpEYpwhxsQ/GGmhhfDr
QXcYRe0tfJ6N78btBNR97+QkoBXn6fnW/MrfrAIo6Xqfj5zofbx+bNPsuTauspKk7sKkGrdZZiBY
K9qg9D7/F0aftnQpQW3ITEliZpqesYD2xDSl8BWuFLNdt0PCAWB4mvUdWUwLi/C3DCbFkTDE3dzW
aFqwrmDkzNFmV1GPZlVYyflfj1WKO6H5VXlKRyP72U6ucEkaS/nLZoGOEvyxuUPNT87cpf/u80NE
rk3ZCChTJU18HGj81nJInkHDGqrTzagELclFSU3CA2lcn645SNJDf+lPn9HPYmOLMtAIYCjqYbFN
IwOOlUQt74y/LpsR6/WNDkRCUveexUeHJ7XMlNtcK3XyzA0Yt/xTaRlQf6/FjSS7kX5/HwOJ4fZd
korFDgtPHLYpbNDUWCGK1BO4mbW/TjvwHAVxWwJEc+NgIzTjMxDbkI/iFGXUcWE24TrpZMZV4Yw+
R6Pbc/ySrZYjZicG6veIVh4/N9aP3VP5WSdJoNgOw80FfbcflP71kT5GGHCoEii1X+IGHYjksoo5
VGxlzuHPrcqvX4pjNYoNea4DjW48tTgxCvzPW7KIvxjafsN3JMUcbkMC+zxiC75Nm94WKzQ49PDG
iJAmPouzTucqJVGp+bMkKn2sbmsZ9jMtThS18KEej1UnP8u947l6hY2F2SGCLwwo9yRZlCg1Bw9n
kgnooVVifGhXT/7IxExn+qf6O4AEHvhfa/Til6w6Jq+HTHJej77UbxpyRMn4OVMxUfz7WkSV+9eQ
wfv6QMhlU+Cy92cPtD65RHUB0bo1UPkhF+sMXZ9mxVWRUYX2emNMXGF/VonhFHQdz9e21DJyKIZ6
bbyE507kSj6NIkjkMZN492EsCz9KFLRjSTGu1h68XTLW8I6l4M5t8OrCXp6SJm+w1ZbKmIwdskic
hT62EZpRDPITXqmbOqwTgg0RbHPxG6eqMUVH9Bor8g55Gt8bT07AFLf2NKg32/0XVWTWaJLctwxr
/l0YnyIwnffJP6enWF3i9DD5b8fa1KYOi3ECo+BKRmV461vSUKaWvskVdtMhuYtVG98g9YX9Qts1
6TWa4e8/acfa7++/zVZ7TX681iCZPSrgHyOnDnr9TXuBTrH6RRyFyPlAvcArgmc74hr/AvXeTE/1
PMOKkofpMJ9hcBtfs4u37/5W2ykzh3KKNVzHwnGTUsVivfJkbeSWSlV3xLbbX2q6Koff9LRhZTjN
4HuwacdW8KXa9W5lifyEdwseXEM0jaM7VSIR4zP+P6hM1sOzbN/2RuJ1llxfNpGiLu6lov6OtdIf
8QUrrRDTofDSHeI8TrsgZ3gdTrSEfEzi5rYBsLIWqx53XTiHcli0kmcdkJQ/z8kbceRsgKWyHQDw
PUAn1Y3IdFQZTLsBmvv8zSG3rF5BCGPpd7EA95Y5FZuVrfMpLLG8mOhoAp8RqyIeWwanUNRb1TxI
bACLi6hXPcLr14YxD5WQoEVmZ82NnXx05aLZldBXU+plvDI1eCKrA5nvONObbD82S8Fyw2T6UNba
b+E9fJ+6ueDsGJCrTV61iJfsazwNT/+XqHoHAPrcTtqowMMpi1EqrVFLjESbECH3R5HFYMOVxOVC
jp2FAOPDUfMUbkAGIIqbW/rfphIZXy/n9dyFpHtG9Zzg2ZRljFLKJ1iub3nh9AGb2kGccS28UNkS
Kj2lKrDRmUq9+hq9yrdtJw3TMOwuWfs4GWd3oqggKScvk1D5Phc243llqyBHHfAH01R6KassYMDe
OAvrYw6itlK22mvpDtA+xjIgokPGgHyi+aVTvzVbAc43GN4cV0vYleTbFExRsZcMOcpCEf+lzL0y
wfp9RaM+WK0RHdmPuUkyX9huOrnaWeFh3dAQBmlDIUbG10DDAquQNeNWpc90MSOn8Z20XMGP3ws7
8LSjoa9qjfWH8sRM5ibhc4dYkSQtn0B8dRg4FxlbUn56HGIWAI9Lmpjlqo69voBl9YsaKDYGrpDT
WbzpyfQX77IbxyaknsJSUfJTGZicbOyZD1pMh+cVwK92ZkGMrUsowrACldN8M83BSpKenA2AYSnD
dPQSqKt3HlwQuRm9nO/q9/lte0Pi+VkxfirI+OtIj892XDmQQhErIb3/bb3yDm5LSH/7ws/VgQlZ
5Y47mGZleX9mfgPAk+kSPesslU79Rdf40hpgRA8esG2jqe4P8ku+SWnuyS7/jJPSA/892+EVVZhD
ynSGszCiN70/U4bBjwODLl61CVTXn/BJlzseRzpWB2RP4cxbSP+lfYtEzfu2ktnYjnDeqKZGO+w7
2fjzVbqhVBjYg/ktGrPClbDzaT2THlpKd/Kt5AgLime3JMDppW2U+6f8lavTvv4ccjrUvG6mE+1v
lcUipENHKU/7NHT99QrCbGKw/ahTwDY3/cbgGxZlxpO7PorRLAK6R/FUtMMtYt47XkNQKNsUK79u
yWpKyLq50JoYXoarj4NUn7vcSQECgVrixEPwLgRI+7RpiRHwPPhZpa6tew8Jpli77wVzqVrc/NhS
Wlt4hxrIudH/9y0GcTjNqmon1qmWXHGch5bNzoIN2bbxluOwwLRbhgQpnts+9Mgwj3lyJOHjH5+4
1nocDRc68yDo8hLnrZcepyUwx0K66ej2+IbuxK8rHa1Fna8tRPIwXHZ1tzDbvFOKoHMHXYtee+6X
+PiYQbSMqfcWssehQWcZyBwOOl1fGoiCFOu8Fiu8ChDvFGiq7pipHhxP9BnHVRYk0Wqjhvptz1zS
iTOmKfvNDSkbcbK5t4fo/JjdmhulVuHeyFOCjyBrmT+H/aT3MpfHmtqEeqnhN4SKuD9jwDRL7LCw
qLsgNUrOgbTrx5ZJKiqNQYpQpkThX29K0Yq6RM17rqp1eb99Ic0cKiMZns4+HeNGNGca7/RYolAi
eK82t1spsa58fBSKMNgW/hw+oQ1goV3q1msgEG45H9SOhSlXPy8Lu53OzS56/tw4hiXPcn1T6fW1
Oh/QMBTyLY3sDL4cWoRhhV7TJdgDAvyTHhZaoNnbeZ+pM+PvhDep9sqqsVOk035xJSvCsGvKKw8x
KxG/cxMXPzKLnynodgM+R1MW9p3GVGRuVsfuM11X5pGR9ET1fm2zzMTXfAa3kfGnaQEDS0Od/sxA
+p2+T+b1/5IIxHpD8BkF+76NLD7TUcRthR079sLPfpzyPCPdnhKGoZf/ESnem+myIOYI81hmZ92C
thuQdvQemn661BJYMzpEylnY5QJrL/ebHTFaNfpD/AqWtPkUAzuxucW201hwUQp7rFbmpwO0+GnR
MsFiXhF8CH6c2X+B3d/4ZMTCAZ8KnO+/F7YU6qMFyAd0CR8jdAh4Z8/CiNW/m7R9isNd3NlnS49M
Nk3Zfrb1tbET0AyG3WtZ7V4167k0b+kY0Vlcn0hoESOl18FSMBG8vPveM+iI4AEACj79ybPW5DK0
oTlBK54jOEOG6jb+a7aOg0eFxpJd+ivkSLG8f/DKlk2Qz2QKi87uyyezVzZ3tddhWXxjs0GOnQRA
zuq162Z691/mwG7STSJET6aUmsP+YiLDSUIEzOW/X6Le8jE7npyu4ZzaWSN3Xsmf+drJ0iVwxOif
u33W5ZXh8+yfqELDTVV03ak1jNSwzijrMr9auolyAhzw+Iz3asKBzD3KQvsWUYIY8IRAS1XG+zrH
V9haDczDb91f9FdWzPMbEP+u4hXG2pSj52BHHVHKAEBgTo48Vd+Max3kL0wMMsmVoiLMkzLMEATt
PcuP3uBSAnQiGwRc0CyBnNNEXpJ9hwpHs4uHkNAVFD3Jahr8bX2n0jrjBXwCinW85R3VKsPVfSVU
CnaW+6Jp4yEb/R919s55bbqfsaXjz94y5gQYoJIbo4VG1TUZ7P4Zlr5rm4mVOjkZG929O8HKXEcH
2we64nSD6T2yUzBn/1cB4WPNOVjnvl7yIitP/KDu27J7ynawTiFJUtJ3Fs+u1bbjC5et1yqH4nLj
RqV63vHM0hlnecp0NIgAtB4ns3HfzUnvX/a/LF4q5llUOKZZEdS2wzKY9oicuc/33rqt+7PgjGv6
7JRpXRu4GYOLh7313cSXN8fM/mpR9MS90BM1kSmzt7nyH67jCXeXPoQeeNBXjZPC717BoB9hy3dC
dHiwnyoWq/LuLBayXt3vF0/n1AwCwwToQnJKFRfcuMlS7pQRpwXtOGBdUUJR3OsdCCrah7crXytr
Fj+SAPOJEx6OmYDoRfopapR55eT4UcuV3+UiRzgu7c07V2rkbG9CwOhxHCL+dimWetzuTmC9S41+
Mv/wypq3qmuICGIinTNIQQAkSTg2hyrSqazmH+jVRHLNTTc93NuicCxfdyuLDvmaDLIBUfQRA1p1
fyxmGVJhoDYRrtf6Fl1iS6WiUZpTafkujSPpF4xrnlwMLVZq4UUE9sJfrSLPgOUto92M8aKRJE06
SvaMzPLd+wT/g8/XYpJBBDmCwrSztVexHiIAHoaXO6X1kW6Dn7TPCk2c9lDEwLwA8DZ6IMqprY27
mWGggXNWAVqoLgKayXYA+Lx7wgni4yZVTFuXFVamAvJmuLqZtRzHi8HaVPhPgo3st/NUNYDVbKIt
wNWzdshgFINTN7kUWnV229jh3ss7lyIx7ZLV3eV3+CzwADk24t4S1yYlsywAo++naR02jBhRKJsu
OGwLPf3ea2TATeGZ0Fj8dS9OXWZ7T4tZkz/jMr7torzvRQ9Gg6ilC3RNShyzfeDnu02LP+7O6cwf
iU8rS4ruV0xfKlHUM4BgDHJVkkICTDYqrk6du87VEo9P8+yHBQuktHDujDSaAAnFl5+iM8sWq/Xr
rtpTPob0wxkT9NwTbnL1nfs0AHgnmop5Spse4KXEeVBlgkaDQgixG6imE4G4nFwfyMHb6eMFlvGl
yZexhBVvPHudYzag0zHEccSsvN4FjNBgl7l0ucluoBYpjF4Ct/4/hz2YAyVe+GRK09/KBNm9uEhM
z2M6wzdMUvwwP+OWM/3MxUcW0Fw2OoEqJG9wpGAkGCnhNIwVRQ74nP7UXtGxMvDxrBuAWlIfllhT
Ppp7JEJVJXTNeJhPhFnGIMavvAishEXHTncp5MrG6fERWSBWekEXq6rl2KlBwuaoZFbVrLtVTrdB
8Tg7kNbsoICJPJFWEexKtiMC2WTrcON+8Z1RfYnmckE6oEqS6CTBnFDYPSInQoZrRf2A8nhS3KNo
slsUDNpewICIwvPxX28X4Fw8PDnZipxqYKGJT2ne1ePzzUGX12HlYsCPLmwxWDxgTCLRuniiXjCA
tUe6K+QsLAtm5NhLPX61XLdj21OLWI5e9GS+OTRJwpVq4GlFLmlXIksS71vtcZtS6Ibtpw41bzrV
OHACeCLEFo9iHeEYGdRLSpcTIPBe3LjEZ27dQ/SqmS64JuZW61QcHGHqzhU5s24vBA3vKQKtbZM6
nPD+OikUIvDUTwclOy2HVqhmLoCiV4vnZtE/lmSZr6B03ly6/eLZrGsiHGnyMJwerHJkQRkQouU6
hS3D1m2vA8tSO+PKMoUUL4QVGKRK7KU9+nAvlcq6mIdFYrwMsbDH15AX090Dzi8l//kRPsMW67Yp
XQ9G8Er3m9PM0yGbqaTFP/GL6qxU2/5MQi/fW+qEumKyBkXwbwszp4UjG98cWhbL0XzMj+FtBjzj
CZSsO1cSvYlGp4d4HIxNQ2a2kJXfQUQqop8y6aOiE0eV3/6mIlp4Xf6+JHLXs7zkUrHXfB9xU9VW
mC8vVhdv1QBeH6I4eDhlXO/1Inq/h7swQQzAQ4sj1EhWLhm9/zkP/0v0SMY62Lu8bON8D6O6KKdW
JT1Ixumo8aRe/Km1dEfSqx6f0WDGyY2KOMQTq9wR+eS0nRsyHRSyX2GSzNfGmYWjIP7bUYOi3hhR
maERQdZ7suf9ueihJZ+rJc0pmuYEoZC4YJfUmeWFWFUM270WsYIky2BbHPC9qRiu+vNqupglMLY3
OctGm6C8iPe1bVj5/6xknOg62vJ/i4vFIJ/S1kKiyA0l5O5vhM02PXT+DoP+5evF4v4TnEfvvK3/
cVztMYDDNocH8o4NnWPR8cvVAHx3I+PbGBv4YhPX3fPH59dMKVDDRGNRdPO8glwJks0IpnlHZKuw
T2yzCuc1LafTDAKe/ivm+s3tuAzzyCPnURGekEgq1+GAwq0BB8jpVTE4a+M0/I9TJ6+AxlUZ2vPI
lXj3KK0iqPDqPAN3/bO3jQtTm7WEFA+tyfHarAj606a00qnDJ7f2UfVcBd8dTWYRIXXXMyHCy16K
bNEKtIg7oYYLqV2ylDFQOzpNBYRNNff5kJiZ/NB+yJTHYm8juj7yRmtJEG6wauD5GUqmcdFy0gRs
0I5sk/i4UHfegMr6RN97YVswSnrNVvlh9JiWu4GbHFk3lOsqUhyjOLY4rMuj0nFCrMkhVInLIerA
acmHONNwUl2cvz6TFvFc9Rhc12DtYDTHLi8BFHWRDfbbJ58hhmVYZnlhzIDQnystDyDeuXC+GifW
Qw5lUkJo6eqTA1azl678krzERFr7Fz5LC02Xc/fplf2M0MPaBX7eWrPkyfCiHNl1qOWQKgQ6R0Ff
g1phDj/110dBvXhvanhOQoq+isOsahlJBwGicLCFRiWCIohDZ45Gy3UAEmbC9q9n0eiLUzOdDiqY
eRyFYS+HAhKNNzSjUSoCZLco/fhpn/KZwJBBPFCukRjrf7+OV5aTDJusmTAbveGRUmC3pYaNc07I
cXmmsQxRWqsS9jizjrog9bWrCrMucMpAkIwx2UFDtfLJTBSTKKGNimYhAHDpg1FgxWUeFwicgJBS
X5d0+Z4mH50Wo5AxAbfBvaVDI9GIHt74G4i4XnbzOHmN0cIdplUci3oJ6ZnLLU2J3QeOsBBE5KDd
V9+51xc5mPwXzwYFP/aIw6JhwzbX0YMj9mrUb56Dq0EuTfkWq3BwytJsgG1B170Jtooy0hDvOAiA
uuqXplTJoZcNXPlmdZrzkHPHeRjsXcfXD5NV2LrUuvx1dH8bpyrc4wkw+s9gFiAv/QjdNGmJ9VXQ
ZfaTinM2s6spePvj5xRhxd+fXDnkRapkMdQ/zyNsbYy/6m1u4hp2dscARr5EILm5ckLbx95yfyQr
dxcV86W+EInaKeZYS+aWkhP/wmfWPn/vNZa8ZR0UmDWcE6bUNGF25VNNLMKIpcJsAB0HnMx85qPX
Og04MXJ+DuxaJaKixy0W3Ud62VZQM2Foa1ZXlbW7hTbbSKqDl+h0eDjx6NRS2tTgz7NuvblOVQo6
IUKDwd9tctWWjc8y2CtctPkdryDVscmR8pG+m3I6J8KH8KUe3tCCj7ltxZDkoI+l3YcjNPuw4aif
6Ja9SdSNlHwtb7lmZi59/087piBgLX0bW+FT6tfdW5Eb6Qa2L9F8TR8D05DUVobsmLpM1pFyE+Ds
GBVDs0Ec4JtQWcOLMwRI4gwIJizYD9xYt603R7T7GhVxBnxlicK5NfZEPQQ1FCqJ/Qb/OTdHNL5s
e+/vRsZg2F8h2LwziIczDaCcHH3Rlj8ldvEvb7E8mgMCzDy3yOSPMkfYr6apqMxI9rbZIzzkIY9D
ovFwuyK45uLMdmPlr0Whpp3Q1Sypfy4Iv/m9klYpugVlQsowDXag9uncUl3gdNvfbb7jXRBDi9ri
lfxadLH/UPNuxUfe3Z8zrGYZWSnRWa8JfK88oOSVcO+VlkfBfad7Yqh/bQdro+7IvyqJ+TWARW70
nxSo3VQMFJITYb7vVllN5WVTSvY++xkHNgecaQTt/nImLz5zBmkn7mBV/VKVGpCcfkWNCms909Tl
4abWy5qbNeq51XL3dniVKIcHNRjDOp6gsERxWZDrmH6gOr3kzr+zvoc+l9pIlTHhFJSR3cQBRsrI
Ylgkjk6DAhtXsT+lKqJw3AaqgNl4B6OrucXdLljft+loZ6B77diyVKVihfMc1bSqiAVcuaDuG2Go
ZbTHQBqWmZobOUTkeVngsVvLtrr3PIqLkm9EkXVbTWSeQZbRhOc8PeNDpibby33AS10omcKEmuHu
7ZDdWK8rts+tHGVudVFOlFu1TUN+AIBTds4oOR+99pSrX7+JzhLzFnXH27SYJmG588OF/5PHJbF2
U88kOPUrJRFX7CBNaPcixTVYRcVUISnVzd321sTpjHw6isZTrlI0hQul8SwUbELIQm3mbPuccfqX
k7Km73zMvPmiyOGX3kwC1UpDz0R8oT0TtTUGjO5gcVpOsJ1iUpkTaSKEz/GkxTBENxXegGa40W+M
2b5tI809+HMw8Aj9QoDUbMlagC32uFaXyRm1qUY885TJD1vMMrF1BTJOOPOVgva8fp0mVZErrGeA
e3RD6RkVvKEHi8SZwQqq4R3UJFsml67+kRtEQyEjc823ux+Xqb0ijKmBD/z3cDQf2R6vylwO3dSY
8fjygth9gKZQRhn8REa1Mp+9j5seOElHXvdICDTwovtL/Tmmwd+XiQE0ujHQNS+B9HFVW1FxtpoS
JqlhDZjBSpZUCWgNco/OelMs582DmjevlILUCJf911V9g/USSclCqwUo3XG08gF/RkUx0UGmcSxe
6UUGleA7bj4qRdtfTeEu94Gsa6G4R9NBXTCpcsfa3tJVcS6Ip4Vl5MpOXc8MSBr+sOVjbh86NcZL
7N/1bsx13M+W4Top4+MTTOd/gEWQwcgJUA9BJ8HoeoWVtomGU0O9BLWr3/+Py9r0uKWl//8KVXc5
cMkon8w46F3SOeyPICcbPgtAUUyZ40zvaD5/94eFMknkzzF5H57H01hi+P8UJ0e8UejCE/6/H71M
GyE6V1ZEwVtHSbxuqgR1F1HnaRfxv8eXYuSG6/1kOPo5plqYyYXIXU+fevaPmCnzISBRN0v9bm7N
k+1po/cVpAv2tufFlZZ9JK6EA6Ss4HOcywrUi9UONFSuWgGHw+MhMGrLbxIRz45Df3m5xiCqRiFF
GUopq933rh4ZOvrgMsLgO3x32geSi2f7KJB0r/Kekskcki/m1VKyTEJ8rCI0NBdFUQRj+oVnP7Ee
blB/ajN4q8WVfK9Uv0Lb+Vnfty1JLyzQ47YdNwHLGNWBadWjZW78rb5DwrUAolIceB4Rv0w69roK
3htplUv5aTtPG/6Ak1y5adfOP36mZypAszKhInscLaZ0LhNX/NZoCHQU7XZH117y/0DoCwoGSfEl
ZrmE8s3LDH+Pzd5+vJaWWnxGqJMI5xasNR1IuiicBtE0Wr5YIgNdp3TEPg7iILxg4tPv5beyGTPT
ue26hhfIw9PmTTfqmrhHqFbJrUwQKz56c6QX5ULKk18hRUFB2Xsd6KQJFg9lacVMuhR1xIcWdZ6g
9pdpmgdVr5OYv+23kzcI5nMO/EtmPGOthkvvkcEtcCHxFPYihaNcZKnGs/zyjNfjdyZNBvawS1IS
7K2M+9sWFfFXF31koEi83xgOR6tJo3pyTPcIYyZpvRWFPLvjSvOhRXqN5plaOC7Bp/7d3//MCXf2
qwOescEppeaj1AkYvLH59SLBK7dJAzQgqkcVtR2FSqYzkJB8LDdRY3KWE9qtzdv0Xr+2A6iE4Nsp
4ODNMzNI63W8K0TlHTQaAiY9BNVZ+LkuHYlRKZaou2ut1sZdOnqm+mi+XD99p9LphizD3jOKmkvh
lH/NsdPEdRBc98h44DWfXOPZ6Uj7xJrECNW96gYk52XeYesTJ4xXZ8proWIQSNeMOKbpknQfsF+I
rLl6DEJ5RPcGUJoKVOxkqUrHfuJ3DQx/XtoSu4goJci+AobK4EGfY7anq7HMyCPZpf2kK71ZNoxQ
8qJ2EtV07Up4ZVxAvYJFqT+uTfD81V1O9YoUgw8+ux/1RzBaegtl+IDabbkc7bjyHOXS5wp1t/dE
QBBy26Rzw/eaRZEKCfnNutBS3Vqz6ifVgfvoCHuF3vJu60NFkmHq3DOoVbysRRDJo2LeOKn1Jbaz
y28YIU/pn6EPHvr5bUVfS+PXBg5jsh1RwHfnxi1815Bee+RQNgvrkTBhAs3lo1JDDaZ/jzz2n1K6
fLvYVk4wvDn/Q7lUvjQULJY7VzNN4B9XN/bdKsiJ80+VJ7/A4GWt21uJTdlZBySQCoGznIFDIkrA
dIgDObGrXMDzR0/3n+CrzyCTPbQjVVXhlO4AaKh7F1df4H5NKm1IVV1NYeQRC68/g5KjdZBx2BRO
0Z9idgo6nCPAgfevAvq9W6ql68sRAfV8pCpy8I5IpFTGCL+V09+yppBNLuWN1IIR9sGzkDlwyMOL
loNVnVyA/h91y+NI/idBLp6WzQxSh3I+fzgo2HZaSsyJkx+wKIG/NvTR9igQPQPf6afKG3S2iS3U
W2p/XZkj+PZXYz9sZb2NYfnCwPZGBe7eyM0vUuIGIJFDZnBdpcSTUu13f5Cxg8HqAMLxLyUhmgyE
uS2JQYIucPKyjsTtsZzcVGLJUUGOl6C/feZEVMgX0P/K5JZwuLZj+809m9NoYJvnY0AgtJAZsFvZ
KTsQd2lbRFVPBTo1xr7jEqhW0Bg481lDuq14A3TkHHKboNWWZrEh5z8uvh7NcUC+Uobpp6+4Zntd
rNe7+50UGmIMBVWoyP/7GW1msvdszn2aRYHve3nkGflehisdOclmW9BShJJSByf+IcCftvOrt7SU
nQh5QnvvWRNo5+I7Eo4GN6AjGAsJwmxt3LwrBrRnMr1J/YekQc/zvkv60mZ/kwr+kiTsrlKpRhVC
XKtneIIOBjGVF3LyIN0yvb45sZg+rU0D6jsUcvlEb5/baU4SK+wehPuSAINy+F+8aCrgAxRYbcRO
+cibWG4fKAFQwdamuSDK4hWvFznin1roLeAchFwGXJevy3Cbf1yxfH5AatQm2Boto6aSSZ/7v4wJ
dTQDTzOqeaC7xVF2HOFinxh9w/O9p07TswTyyVXO8Pi920kDHafkQwNN+fqbj8ZuTrVjKgqOXB0r
0VnmicM4yWuBVHkwOrsWKjdyeZq87UyHLoAKDh0n2HKJpi8Xn3moG9t4WgnhMnW0H6JrG8JuJI0p
CsJ9qAOcI5e34f8whUeoD5YZxOmO2/jRcefv9GumKRr1GU1wjvq+goztFPRDrQcaNnEpSAp3PRkf
EgT8ncX6MNnwviSN4vA4AMxiZ2qxota3DF+tC+Fnjzb9QR+DHxVyRE15J7MIPtuveisdvgf2KZlz
cnXP8NwyXJjeDSPmt2/M9JiuPmIUU05NplVIO+x7FzwsCSfTP9UqrhKAVpwIgTMOLws3XrDjI5et
zgmmZ2X6Q9b8ZC7E/aP1R3SssSmnk2nuGolhOQ9gV5XIQDLZuL9vKlKnP+z+9WIDy5lwa2vreOHg
epT++gwT02LQSamxWgSDq76FpMfr+lqhIY1pk1zXIRdPCl5DMrVfw560c+fB1q6B2zFpqhYO24pQ
avYDHPEGYjJpfRE3EgiKTNHBGuSYmpSXIGDrQYgCcRTHvErPIQ9jglqZeG4IbnnwiGn/PVqJT66n
vsUHNZMIA3GrskYnazgDdBG0rs/OYlHG86ICVzmWQUQdheEaBIhdB2KNsme1yQ4Tc73zWgr+j5du
dWfFq1jq8YT9XaQcp3pe3IrKvVvAylxeXEoy6Y+sPjVHMDi9hdyTCiuraWP8RnXggy2YVtJ3V6Zo
yztXBPmqzH3IU4g4X040rJrzyLyHUTAMZTImGPBKSx/P7VnUMQaFSSRUz87mhRhcbAoCccTsOI8v
EGBVP7NpDu+xUTKuqtDqio8fIdEdvx3909Q7tnpAxy5Qbv38fpPOa7jLU1w8lq87Zt/6CtYSCFTI
70hR0GujLpWb4U7ug6lxiejHC7aeRsjOYXxGhqGMxvw73oluqIgZVoMcY59jrAV6/X6HpBU6Yk5Q
9Ss5+WzeByB7V3PLCc1fqKhq0Ds1aZ82k5Yw+nYLONGyQzRP+BeOGTkDXq+GIMtdVef2zhLLvWhW
vefQ4+oeHn7ShVm8+eVSXLtvOL99hJHME74CJPMKURaucrOct7+DfSDN7Q6FJGwK0WB3tlqs8+Fx
tY09PxcMfQldaCJg65BVUHKo+PIIdQxUzGb6FDtWTMqe07BebV0hYKCY7xXLPWpZ4wdLdS3EuJ+9
8wkb8h5MIwJOiozPg2BHZNQt7lkllxohJZqphb8jsw52ObNgJUK0eYldTKAfceDvijWbNGWosWd6
AwHD6ACQcLlVQOr3xr6pbGGeVVvUXIwvjbui5w9n3KViaph9M3yagULEn+bd7vXbyU5MTrXu4c2a
MMEF4qxcme3+dNubDZyz1zhChc+BwYmMlij+LOLNFpDQwRulfXPPBnjEPRdPEKhu5cLW79YqBbW0
41thwmCeO926rnOmwiebJVNWKADeZ9T8Pp4t/mP//Dfoi4mP6HI/zlRoMDy8+mjzwGlQEPg1cCQv
rDG82rQDLpfV+1cOLTHDcaVvXK9CoyJPO4DbVfitSvWqdwq8dPnyP8KxzVKKlAoYxy8ZMj+V+uHN
Jrp7fULms6FiC2gglzl+tozRw1zJqjbLUdjbk9C5MdIMnzos88rI/HP6oSOenuYHrBZOksK11QkU
L+AiPDsKICspRlCarcREU3GDAgtViXNAxfvrTN5FmvDn4Fl7hWqlWxqhreACC6rHXH8IGNnoC6A2
+Cgj1otYeyi5N6xTetMj9eE3HdJ4KE5P0P7VrZew6ojnPSpfM8I/NrsAdI4K14IZ9Nz1C489NBV5
3GECOK0nFgNW/GrZLhoHgAuqn1bz++TsVFkm+/MiF0ObLdMpEoqWmc3hNGIsq1SZ9AiPYRkAN982
TgODX2cR3vXOiWdatOUMJpCLv4oNDV15s8whiHf2a2ea5UW64z2qVt1cHIAVZEpJW8a/7MV5bGSz
V4N3CGmPA+x49MhU5iP91p+MoQr9Umv7VJFaSkFdvovoprWjfnvFb8ORS5QWBg5m1mK2Z3FnQJn/
awVglg8rkTJdipCP0Bz+A5qUd0kWRf8fnd9DbUYfVLutkQqMwUEav/jRWKd3Hxbxbpb9YqcmUWC0
REJyReKbF470M0JTJ9X5oUbcWjXlXSJtp6ykzK9WHA/TugV3LwvirIR2SNNSzvZ/YM6wvmrGsESl
PKwksAPn4iv7ViSioyGJFxs0N27khvrrq50/lZ2xDOGuGA+B7vkRpJDG8ENIgwcyPsqAZ6dXnm/f
VsVPRDz9rP8VB+UowkY5nAWtB7Mhi6BklW2XTxwgoRGrV3HsWXoNWUJMsFAG9gkfjqRBjgCqRB3f
HmSdQff6TGOvIFXtct4zYmZsRSjOU4kN+GGoor6cTSWi7g26t5Cd8QbCp08rg2SjgtJKMRSiOC4G
rULyVBtNTXmR7x2yEH2WPUKQPw3JchSLkFEt4ZC9XQeNNRfLw5/Jv/MwQKfp5JEvE3LUh1ZYhsNF
ayy1G6tQim+ybJE3q6d2oXAg2VbYu6PFyqltq9xnAj5T7yjfdhyQ4Gsda055ZMn+afsm5Xo6yKBZ
P1nth4Nal3RV9i19cQ6cMN9BqofP0P9L4VTuR9qtJe4f+HSRo7f897it1Y+TxevE9rn37tXdtdN+
AiGkErEdHhfsbmDwwaZi89ZEW0LF4fLHfErSumuhNcYpwUkmJlckbxyP5LIY9IRdB2fnQyvg6GhT
z0ccAarksFaML90RqysI0gB7sT/asq5iTd7yPg6FXeQDC0RtRutpfZDGOstH6YER1vYI0r0XNSnS
LTl5EcTW1sHEFMk2LpoXBtiwLohO/n3mOJe1jrOq58kxAZYmbNAjEG6azts1XYw9j39BsD6Wdb7Q
tLVBts9SvtjIrMPXUbBGNKnmyCpWU03N9uei9JOzkibiOOF92r+/+UWj6L5hEaqtg1KxC1Gwp9m+
n5BMebSSmp2JkJFHjChTPgVAkYXABdNFP2SY4xm2UykaMPQS+foqrcLD4IiuSeDisUB11Oo5ZRKG
DIaGhvcxjsVIiU3h8Qs661HU0+q5PIPB30mJlaIO4nn/OEm0tbxspA1Wr+j7258X/O4wi0wa2EZw
eh24MCl8p8v1otFanFoUNP3e/8Br8jGUFj6T/WN6kbgUYa2MP40VhmOld+9HBTxMxc8uQcgdZF8n
4eaIdXrN5WL44G9RIwOAqWF/m7ttz0GL6iO3RKjArpeSvw61/+Z2TC1FylWPs5LQ9xEybvMSf2ye
iUeAl0Q0iUQYhVEjL7+0Zu02kGzCmEWKh19ttR8GBQyrJjU/ZFhq2eULgW1Bdik8sw9NQ94WXrm1
EVjhGsOuC8gLODoH8jzCEFsrlVnsiLcRcWm1E4hctTty1qZbNk+qMHJR7v6px649ikANFpP/tF/7
TTApgfo4gNqZik+nFfxZxYMyRmbh1qvcC5/Djj/FPN9mfPYxbbgXRUDEXYj9EDOop2X0H2DW7ahR
POm/5ni8f5D6G3zhvFBV5ostL+iJ3dBQtwB+yllfGipNg6kIujfIWQM6YW6PF87QzuRC9lYZRe6r
KiMb3VmDBtLucngYTbUndK0t+rPtXfVFRinvX/qkzIscRPyxIpiHtHIe2osn7ImwChyexeUl7cbC
+dsEr0UWWXrM/lquLsNV1MuYnQFJn/DTj93BKPxLfkxjWf+uZ547zoPj7nSi9Quu9bOGckzAHgGb
gHQMsACreC4FAZpz88z7n1oMlhH44w5/H5FeHtZEfUhEQElr1KW/5l8eC7IUS0CduOiG5fub5+WG
TdaF/C3Y+q/zLDbk/EBL7E3kR/Ii074dlV8AT3vgm8NIPcvTKQyTI9qZoTfhotI5S6RADgeZYOLL
OmZ9CrU8piBM/Jg0NQ3+pXpAtYeskvkWyTXvmq6fpPdWzjXY1O1hAGQ7YYyOAHAxSULGP26EtN0Y
bR3eRO3SbPsFkwBW8jCjaKCuEYRTASNhYap3764VwmRbT0/10hFIPjb9At3blkvBZILEbR/zS8rz
/rfz/xwbiXFs/PlsYn3x1C6fqbzFBuooa5odJC4wKSNtHadBP0M0I1z1ChMOK8RCOIZzbBwC0Ji0
TXJh1k072Nix9MjcQibzYpbRPvjwn4TYktXaPnIVdeUln0d2H2KxGLOefFNOZCndprqul4cWCwks
SKqfLpfYFYSIPavehaMZAt1DWF/jqMTaM/AgSAszkDW8xv3B/HzZQDtoaKsCkFU0ao0AKwE8Jirf
DC7NCjUNrfvHOQHQUIXsgFe6BReg3NCe8DWbpX4AfaBNwZHJ26h0we+oPvQZbU5TZgqlyqJAXoiD
GEMbNDzp/hNZgOi8mZyYb8WPxopgZDLtZt6CMBjQSKLmWNHFa6gt5H5ktuNIM70nGiiQY4JbcQS+
y3DspGhzq/HHPChR+/Ux6EGwJhWcQaOvlBHwolHXCOnyxNkMXarbeSY0R1SSXT21byhOdyKF4rQq
OQEkUDXiFLbP9jCtodtSFnFvnBAbs3/7vLNUePMn4wqbj9x7W8WAilmvOTUzYuxyJidDeKwNPXuc
BYXk89usNSqpThzOosAkOTpYSOXihahlITCy6dfEc2rIa8jVVIJXjnxwOHS/mTjtzT2Yq3Qwcap+
fdS89iuZf/yE8KCrAbB1bsq8uUpHFCm+kLKtr/HNnY5n5lT6207Pg/u6aJE1exYsRrpyj/xO2fLQ
2378i56JnY3jf6lBPSmKVG1AkfnzoIZkk/+tLv+RvAnzLKn2NpXzQGLAJpHxXycEVTBgcPKKQXNr
jKwlO0cuHwk5/yr5siQ6nLYcbBP1zYXZVFE2fyyDOa1D7jYqpIP/ZfDuiDlGq61QWmVkyS1/hVwZ
SMSgosB4eJMtjdmo3nb0Q70quycklvtjdfleIaQ4Abwys7D3dKHEFnIJ26wx1mY5iBdfUX4NISKs
TFK8cQ0QQoB1sM7C8+lhA1T3h7zeihB8+L1ZWHpP7pebY6yBqCpC2CJvSNcdKWlGYStERH/hTahs
Ggn1FLWCWcxgI9uywzEVAopqwRIFTLIPVdJzM68dpk5Banoogj3zflk6uf8kjLgRJrxj4cGBL3HV
MUU9OuTQnh9T7LqAxAfTtwxLs5EVPukReL2+F0+dVvOkhRUfGzwI3hVvMKWVGClll25p9Rjqv00O
sEqzpVZvHJzEzZuD0/G8f70bDivt186+1MttI+DVQSEq3s62YVOQimHjskaYvNWuEse1hqPUp8g/
BNQCfZkff1iHR2ZZj1v2Fs17hNxdJFPl4whcHS3c3wFRP2qlgbKakZgosGeF9p4W1Dt5ZnLUp6Dj
JiKKJFdLUFYxNBESGkM1ctZo1pBX1XYk/lrPj+dhLocVsH+I6tevAsq6+iRk0dCxXMQnHs9hssHa
nPKSXB0IaS3VipatCdrocLyA7AnZ4nUkzVH5PTdc01TIKHpoC56R3ZQTXe96qCNBR4nEbuUlQmG4
iToy8xqa99H/g/RKxe6GUpK3RgR/Sq61MIGT95elCieBlHgZqU6vX/JcrP+/xWsVmieyKfMOqzXH
DpRlC6WnW99tDTI6mNO2m+GKzxTmf2oMYzLmuBIFizCK56K0/34zUhxl18QRVqVpv20TmJZw9kA6
XlJs6BPRF0uAzM3ZWzVXSqvlmlaOhOhmc6j1iY7vo3hFYrorBftv+DdVsk2MFr9T0cubwV4mobi7
gpGoB91hz4682dE99U607XsnE+HRKuNilhpul9c3prA9NbovD1dl88SxH9lMI0aOpswvpn5bYKmD
eCkBZZYis144vqYqJdSDwlqpWG2P9xGwQhJ03ZqspWsdVZGdlNfzEZ/OEiOmTFgnPWOQUOKwgCkx
Vy2lMq+RktON2bnOTO1bl9p5Jz5j28apNyIx4QXQZKVsoh/lD0wVQAK5rsuId2oGorod3AvVPbGN
RKs33mg3+Xyb9Pqh7p2wkkNESVPGvKiO7HOzIZ8kAQQYq6+x/H83H5801GDh0U/mGs8LtU2vccqm
Ckk2bi5va5Ohqxbg8zjQAnbTijUftJAxV9bnWzvr0htELGql9hTe9KHvuXyh1p+vPN7dcusHNrIY
x5sAK2joqvkbFB73iUJdu+V63nUZIic+gl3bVwiunt85BCkZORa8qkfovta7eZNDQ4+JsIgUjwGa
O1pM7ki/m96pl7cRvIBGYet1HdBAsuj0N5RNnetvuyTINnJS4dT2mMSKaKXq/9Oci6w/KM32sZiY
y3XcMT5fL0NN+VWPXH6X5L/rezHYMS5aV4vY04puZcPjUzhZe6NZdECpTT0s5eZ6SP3khuGRjQL/
vVkwvfsWxuuUsNcJr7XrrEcJwLRMkotUaMADCQpiQVd3UH4eJrPaCEJyjfCwg016RCbXlmpc+pcS
5sCCJ3Y2vc4/DT/YhQxVirb20XCrhVHOrzGmhc7uV6cts/vzpw+vawfC2dp8ng2YaIk3S9mpWaUK
K4aOJsVGV2yn3x3u64gSOkkvi02EvyEideOUoVfzoJ9LIXJCApF9LgWw+e2dQkO+j2+Zx6QqamzO
r7BnadjlaHB7UY7zmFRcsx20xAaGUqPjdChUkEnLqhLq00yQJHnVqw/uONus6S0/gnvIvYz+O+ap
twYwpYh1Tuelmywv9JckAHqA8g1RYOAWbdVNgHYF9zpA1ThBT1ynhAUFVza/m3u3iowmrPsxuNIf
hUWhPk/3COPmG4jq331s4LymOv1C93E+294yNsVsOnEFYCRYe5zOCtko3OgPQ4U6DFBflqQGAa7G
0hAoGT2ZQNEJrUJOtElgZi62M2ERoNSVypbQ63gRiJb0KqQZxcl2tIMUvRC/V08VmnXF9z88Bq60
dyPWAfCSwGEOA63MMFQi/YCWIWf+RTr+Vm/Z9gPq0EzUvsQjB4n2Y7diAi+38ZTRsgyXNcPFVw8p
xctQj7eHVeHC/h/k8jwD+woBl1bgsLPVRmbyaEuGC9Cy7djKg6cxWym7qfrRn2N0AdggKUjGaXXz
oGvmFBJ5g+wjITqlRMRmNd141Y7fhOUy8BKfH15Rjy/mZ4cLY6zSr0kfVRJCdFWtxtN+/GXPGYz4
gUzIRL6ddMdGGbAyvYaKKu+mSzi2sa3240tpJcJUqo45xhA7yZWOhNKPp8i39glKqq1JgzWgOXAf
zgyVACkuq3l/fAWy9jWJxTND3j3Dqfnp4QQXp1aR/R+ZiP/AUX5sbspdO00YJpsopqfHhUBToE+4
7G6FJ37JoT+hvVEzrJf4NZeUxLmXMwzBIGWOaSodYlYV0XkX+74N7Hv39ikaFcn5iMYDuNnzhoTj
M5ZD1otPeKFJkak+28EyYkdInt+2nUMM6bsiMzHd1rwHeLc6fU7gkMCa+p6E/7uiprPD0rzyY2b8
P98E0k+BnHK2mSEFzls4mqaPAWhz9RPdm+GSXUSL+IZuLgy7xEkEGzcLAEFMjg5Cjy92p+YD2LcF
VDFBbRE8Yg57+zS15leXG1L8Zsl9nPgxsZKVbI9fMcvYA9TU2GkMsE2M93Upt/qMNDHxq/hbCBR2
IiIz6oo0j2+izPro/Yl6s+ftdgsWWTUh1hQxMmytbaKaAuGn0B/BG7n4jej00ZIdmZy9XdmJNWsZ
kxcNcHvbceKcPYy+OB+yQiPAtmYKChTmbRYWizdTAsVKVLJ1zrf5bp+1X6SmJ+xl+z0H4HJgijdc
09A8pyGBMZPxlQs56lgJKtxgSWWNwnrd9rSAxYxxWBdYpJUAzAaFnar8DGlKySQd+Dm68PNGedft
StiBiRLrE9VQB10prOVLmW5epwBAKoKZqybUwlTSFTv2Kpgn7yZfOVdjgPPZ2V/PGudjOBlSrb22
2BdEp9RtpMWe0F04J2RXjRI4eZSLRMt8EN2OIzmWA1Rsc8XXgzz42wFdpZHdb5UdJjUYUkU7eNxW
rXxH2t4D61e0NkkBEkrYn1kacykhHujAzHyMBrGYQfAW8wSWbpW4a+GtWyDLEQhx+gx92o1ZHGWN
tmdY5nlAfOjtGLiNc1sb0gJohsnkfX3V+T3T6+1GGLrfTWCB9KNq9sqPuPHVcSfzBXX/9Js8KnhW
vfNUp79RVK3A/Hph5eLODH8qq2+dy7CvGRu6/KmfWtGJR5J7c7J39+gmJDdnzY6jLlGtsB1BPR0f
3Fb6MlDqd/PcWu4+JmLwZmnpov2zeE3h6uPcREkjQzhtjY5H+1pcWpK7N6WLrcm40RACXlUCWQpd
NZyQ0rJ7vZmIoOLwGqCnTSSZJOsX45dSMT0oL8MVfzylq77C6xQt4DybuR1iWVPfYUEOxCqP6pXv
duLQHwjuiW4pvXY+KPgnjFdd0ceM18lMOxqF3htUa+bag1taY+iZNudOGiawIyUTCoLnZzEzGOWt
nzjWqX/2hSpqps8U0Hk7hNvekRJEda7DVCaH1YmUZeYU23LZT/Wz5Fvr4HEdxJu6uHoXu46x5KVY
25HfbFaib+GOqLrpLWimCNQ8hPlDHWDFlX1my9o7YaR3D1+eARpUN4MqIjCYgAcw4gl9OgYyTdip
BgZaR9qswTJ9DYKoRzXgZD+ZAQ+2N8IrV5yZZgbi3Xu4zCFocDXSPTWvd5+RqqBjb5kzkHlFryQr
rX8cZAJ7Ky5ewcPXZYZGroHN1AeDBpG+Go71LBqlZOtNFZhR/ru00mJqCw1vJnWGzC2zsP3kN1DO
KRkuU+d2K0cpqmtzbVmLOdXn87O1QqvdwiHXjtiYIIg3MhaPzh2pAn85EaWmuwkHo18zmlu1t3xk
h976MH6mc1IfKofgOVCIt4PIgZLyN9FNmegfdx6rsmTBAht/1+pFE2nuTq5q4gc8oR+CvwEZj8OF
erpE2YdQjA7p7axYeRWgUZFMbQQnltXINmeuUZ+tHdnmaOYbANgTaj9WWcPuhEEpIIc7mS1iLSXN
VxD5L3hB2i3mNJ0YJBuvMTB289dO2OO0vA3FxsN88TEV1B6JYfSeB27YrYeAwhHVy7sUGHBfGAUL
D/Pa6qmd5RvlTCpbadoLzQ1sNh1w64bKsr+1Zv9Wr3Fkr76XoWm0JglsRLi+0eLqOpS4Cb53okCU
J7C6qF+Ljy+gaiuh/6yJY3QRpj5NL0qALAjpi1F8NcGgrWSfeOUzrFR6LtqAEzC0CHQymujAMKoN
Flrk4+CRz8zzcTL7Jn4xCPU8AB/1yt20cViEVm6GO6LznLS0pGDkLIrb4qvp+AgN09I91z32Choe
q+bRpETkpLerV98RcXTAv4s8KO2binWcsxGES1C1GshUTCxuu5fr25C0T8unc5Vx0IYJtprXNDuN
1xpZl3pPjCzjADE6+5OWuwH9dwdMelnP6dPEDBnUz1FZgoNrxlwkB0HsWHSyFswwKqB2RN1r5UW9
PRN5VAVO5bVb3N+IQLbuS2ypcpuGyQo/dJ0GCDYg9SXc4hWRO6RJoRCCoKrucx4jJ289pvkqnXCA
92/d7A/xe0BzKmWd6znqmveUBV53bq8QtnrMih//Ru1wBsKJ9DHAXJ4ups2MLWYdhkg0ejCFamD+
81zsFAK74gNZtq5B3EqGndQ1AcEl/osIxHqLgKuDnv1wHcDLtVVlwucfk6HjF8HOeI2hhZzCuKTr
AfP3Y4NHMJZ8xqPl0sDl5d+C5J82eUugauuUieOk7XoySm3WGhPUTWcHZkzuoU20ZjxX92o/aX+2
kEOHUq17NmOP/5WU7qogIiTL9xZOzg77oSi/AsSXIhx8Jm5M3qKJv4JUmrp8uNqATjBansYX3Q/q
3gCrEHa9+TxcO+hM30k6e2x4/SekC+Ce0Ds2jVd79K+iTdC+vyTGhEzjAJW/0QDaOjxZ5Yd0YxIx
aJX/pA1ETLNDD5undGnV5oP9deIfS8OUhYcfVXaUlK8u58m2UmwtolFFdh5q+nxOy2u4sVTtI7v1
EQysr0POh/48lnpsLxRU9UBwqk+BeLHQEppi4U38gfm/ipC9g/Z2Vz+hr+N9ZEfls4vzxBKOm9ZO
njI2TCE4Av5SFzO0LQ4KUkpELCUGGdSoqSe9LsB/uTcb5h36zWkFgKR6o6H2J/y5qhTcor2LNNHD
T1RXvVWHXo5EIYUjwkOXDcL8QTmhwj3oCRs7hUYBwNGbOG/uaQiilbnFMb63sCVHx7r3ea7/V4b6
oobj5N0D1VYRolN1It+xmz7Li1oy6McFCYOHRDOXji9xMHmnX4724SxPq5wEE8pBJZKUxQVpIBKZ
6fdFlv0ICiB8mUz38t1pRx+sFTTNFsKJ+7MZ9WTMh8q7OZRPBc/NakZzT184veI4xMkjYNSgEWpI
tvATDKH1nwd+J0lHfTcLBDP6iSHrUwGj6yZ5Ft1QV21CE6i5GNZVFdEQGNVkXsabcBGkj/sn8jkS
C2zBHLOBi0A2L1sxFYlCM7EgM8gfU7q6jESIm0SNywIauy9OqWLNGitBBhkaV1KhMk5nRsO/iUAn
GpyAMsGgEQXZaYXdA15XHLqVRGZy/UVZKIrjJFTNroWed23T9VNBkG3ruWVuPxDkbtJE1Iae6Eyu
ocZJL11hxnqqO1yZEjGnhL2cBtAUM4+Ry7MpCRihwb7sH1GuYsHx74H7r7HrA/zCvnpvpQUwfvOh
YjhtNk+KXJvOl7w7uI4+4hgLyed2n0DfgXcIeJ+qzjlR/Z01klXXT5NjnCdOvmmMPGxGaXp37QM2
aTqQChOITZZWH1Ie458/nEJDdSVj/6qCQbpgj/kN9ulOCWbKa3irJvQe/RTOiIubMkUboYM6wxH8
y6Mq5uKgZXktM9HJP0l3MTtGAsDli4ylsWS5/hGrMXJRdMgiEAfv6rnbc3x3dzFmxYNY28cN/k5L
8KsKGvSCDgThgOd7A1eIl9mEosWDEo2tDNO/6+ZJUvDo/yykJWhDLxoZs6oDYLIJJYBykl+aosKg
DRxRWfkcikgqoMJSrsGgxBse07z+70ufGY6J2c8jvbNP58e0ieQgzaSr7BzRcaDCuW1S3IneNh+k
GJ2fi3M/N+jCpyjX4Ok9Siv7ajol1s/3cezN3WIYGyHSIjgpuFcp9NBBlsnn3H1X94xOy9rfAopD
5Y6Rr6DpeADZZrF9XfnGGQYBnAaKKiYux6lhdZ/1fKfKkMiyDu9upWNNhv6TT9FaH9btPrF8J0AK
LCkxig7UxOf6xyFpG7pj8xRdls9mtNs7NY2bTWzSkALD6NpSNKaZrkY9epq7jYcw99mrKVfDKcnc
wf1VLN4mCab2ASsagdWb04lQ0IKEDqXGTF1XzY9nuZZwzoH7ahqsRqHYKtmbRfzWuP6cgdB1Ejc5
xnzBDCMnVrW3I+CMCInJZuyESgUqxeoh+MUqqwlaKHuJm770DPZXd/79xnjC5Qi4WpQokrTwiM7Y
PmENw/a1iSlVgYOXp6Q1VPDZRFUr05SmhynlU6Yow1PtAwO7xum4A65sjjzTEzsZ1RskwMwKnRaj
uu4U5vFFIKAhcdDvbS8zGeN+1c4SxAhZ+akjvulQCWI4y3vTNcc7HXOiVaqc1hVzhGpnbLtSwi1/
pkUKHfAVgtHdKthh5TVTAokRaWDERNTYwV8QeG3Dp9YAHi1p4zrCA2f+AwPpirFU8kE5N/J9GDl0
aWEfmufvUr0vUzw6zJjWbV76TS+NLFr3oHuK1a38DEmxtIa4C3vgUchX/NlpyuPByqoPXffYtHCR
EpMxsbtYxrwRSILchMr6pHgv1FhKXOkB2duosxlEFdlh8CtHHMxv7iHL9IEC9C1LRORx79S+gyy4
+zdhEupV722tHycQqb7qHk6j+pHLsg1h5tEWcI3kVV31MkiZ8P6EBoWQQK40GWncB5rhO1wDDbZC
J00FVB4Ohw+XffLyqHs6NQlywD1A4L6oIO8H6zmzLxcjM8hDqKmB3z05D9oGxrgmhYObhnWbfqLa
745ja8L+AgBTvPaQX/I5d9h3o7RdgDwi6VxuXXA+iq44BoinxOvnKzLukfnHDInKHXyu6v4kxEly
o7BeNBfbjAXuvKGJlzq+SgtGGzvWirwMrgWpu5XKhI/GN3+vgkAHaCsmTghQSCrnduytwjCuhhga
TEYvy82lQQK3v9xs262uMRjvsNfQCXa5JDb/2hJuVBZAUgYFFS46oxwdqolvPBfi+lWczrwHzQub
R6GLSWtVWK7WtnKe3iUJ/dNSasMUtORa4crTtV+p5Bq8YWbhesZbd6OUZCY1t35phqskpmwUN8zD
8HTLpNFwC8QW1/dU0wRquZnuvHUEVG0fzQT+Zp6fcDjnuiXsnzedt9E3TMtUWsm6KjRheMiyfU4T
6UMQfNFik42io25LDC4mutieACXqjMjPwZcdcN37u1Q37XuW3MUpXeuhlF1+XBnYzl9T9nA3aNbz
4zsF7eqHa1ewgQzBGwfcpQeThmYX8bBBLr2qYiex/N1+HB6gf5jHFfjySg9AMVpSoFNd0IhlVuZv
xeof5JmmVbWoXoWZNPL3cexG6cEtX3UcfituSOVJ2HXHMivzZFiiCQ7KQWUTJDA4Jz766RGswjiM
WKHbINka5cUS6tK4mo1SC6YNYTGSM3Ni8GfoAqkb6v6+Rivfi6w+hLCEuQZHWYNLtezWvb2a20U8
TIzh1poNgLZT/F7RX+Ap2fg/m1WRuSpT3fwfbkPfpMnuls5RUujtZ/jPwyF+OMans7rdnbOx3+RJ
vESTJbAhjrXv4r/ZZ9e6wzF/YYHkNGreoeJv0eczKiMa3bjU/xPiwhrsVwpu0vhuJoEQMqkvdAix
nNLdRcVb1v5MZqSTQchs2WugJic4rB9b/82+Y3I5l/Ytgv7dAe6NXaWS4Qc7gFHqYcH20E51woHP
wVjv14uMF8+L1BoP0a8auYaRk74hkpKlJt/evEb5DAdL0/4xi6veRxNabfGFrUjQZzXK3ygrLYqv
Hzb1PlR4SC7/cm5YPPEgriUbhbATkYLgY+owCS/ppCtmzi5KEooLjJeCnqseeYGswHsKEfddaB9Q
Vj9fFsczycQgUPG0Nhk/tMiu3/6Sxm/W98vwJILg4GMoK3tJ7AILQk/go0WbB1Ff1BxracmO2a+E
SLbczRxPLm8pY9b/NHzOJ72ONKR+z/TfYvpYfw0bT2I2v9zO/jXTDnGItc21il5cqEw2SrL4hyCs
A4eLYQ0n6qU3kAgwnVwLBOaTC1Y8CUt1DVubz/LK39qB6ea97rRpR9Dq30AHwbFieKvgY97f7R3s
v6OQFMtr0uiI9cjzfscIrIzFsVbmJa6PFNaoYzfUWvxXzrIPQCiYouseyCOPbnl29bHtj5JTJkDG
tH32kZnMFe3t/lUkMhCjv6CBHFaam/Z5/vb+YMOWn+z7FpEFzXsqAumrMigeWs+RmYMu0ebv3YM8
QH2EtgWKTb6biAlMn/zOWyV3GNUCqkh9+ykRghNTAcBcLoSt2sxFB0GijmiPifAAI1f2ebmW4Up3
6LuPaAnz2GhoCVHjHI3l2Tgih/nb4j4/3zJ9UPCqperM8wrZUU7Jp6ggKtJAEZJKjNP/nUszcO7Q
USUX9kGnN6HsgnBIFiILNWQp9K4/miLjsbCSEvJs8wqd3UmSdhJSJ3YH2hz0wtnFdrN+6k3pfDTt
k50URbgigA1YAFztSLGRNRmiJ7Zm5PcqMCo/peNti9eSFtslGp7ZjteUlRiNlPPWVNudHx8dsyLK
oNJBRdBHmlyJEXbcFhT7iYEXWtDvHAQG+y092Z95Paf1ObHUzswfRBmcLvUaLM7iRfMstoMoAOpD
KrJIZD+9jDM3gIBoqZ6EI6oUzCaBITJmZhNR3FjzbBJ0UZm4uR4tvpzmsq6HJWemXTwXYiUN99RL
5I9kb2yiI6YRhgN1V5RayyIgklHQSug3ZkZoBNpAhB4+9yYz13xNmWXh6I368q2+mlgxC7cA2dY6
AUsmGQxyd/VBUynok/CaUuqVZI5C2mltxCF7ffT86k3cYoCDKogeRfQ1Am4teAY6ng3AtRdUMgE8
Y3mosYZcsshvomh724sitY0oPcCBXrsM9Bh+Wn2IrS9GqGY/jGU1HZ43O2ljty0IZNxgc/2dfV21
IOFBFLA9AR5AQmXgC/GWDLCr5E3HpiCZlfmRFuxk4OhAFxdPQpp97wNm1Z5n7JPhiLXV6Ov0HkF6
A+W/CYZx9D+TE3pg97E5acdI960u3zRf+lRsQxPNSZaidzygZTfrPDZA3m4f0MfaZNUnrnXAt/22
ZFJ6P133m68UG9v7jBtwCabEuNgQh0nl1u6VFyFgn4zqPhINALh7cF2z6pq7OzjoXejGBlCMmh1g
so5iToPfPz6+tkvPbSHBOctb5V7EGuOUBQWRrk7jubxAgIxPpeLRc/O8FvMIS3Pvy3jbyvLHXq8c
LpN4GyxW93WfWxgQkciE0fnGG6Zs6lbiKUF9IMf/TjvWORn8E/Go8Nk3LkHBNNu1K3ZQnvNveQtv
zyY206Uf8pxM1bFWJd/FcSSe4vkiK3wYF6au59/e7kBKOJ4MAZLUgJsxmYG2n0oyjAUvmiHHcgxJ
nibKiTSxMs3O7gj1OXWLvWJ/UfXzaDHZpWniIwia7ozujGx7VStLzBaZGxmsyv3cG9IVonHOXa8g
Fiy8TXlufWfEd1iXvxbwuEwzXirduHf/lHSD9N3hWPVwPhVHXPuMrwhFzs2TSnQAGc5thRW8w0Kk
BajzADClNJl+7/BhxbY3bLvNMqP6Lg8Segl40cPcm7yYZS+gyTzhi+fgAmeBRxnW+Bqt50qMB/6m
614X0MVR/1gwF8LMSs628NK+w0YPEu9WT8Gv86o4huYoOtznEeVuMSlGO+wb3eaOgMxUavtw9C2l
7UnQJP16bEqGm3qXbcqBzBtYvR80pFGYg+Da3QAAz2bjLkQ3SS0n3iuRRdgF91XgCI0kjQ5F+CHz
Ki/YpMikDGj96LrPMrhQLgSsoVBAQEKGEXDbAAxWKkgw2UiA8t1DioIwPTn5Wn7+0Q8Ht4NWLgun
c0UBqbNNHlVeVv5NO6e1/cYvD92ryjVFHL4d4CIjY/E3Rdv2R+6ua/zaqYIpZ4HeFzkFS/dmExKS
6sV1xzU0orZ18sv93t+H7Ty55W9/rGeQaWpdn3yEccxD50XhpzwpiyBGOKqODfpEFp9Ny8y1t7/M
r9ji0LJDLs+97a/ksHQ/LIa+mjeJBqWcByVCrwRgZo/J8nv6k022ZaVJZkVJCqpbX4tmweKsDf2o
nGJ0g5ZUq1NPdzBAU53yXvJSac5i/4RCoEVKqDHw+3Q8kiiv7A0xXy4vBrB9+/zYW8535Ja6u0FY
Jix5J7/32d/A6M5i1pj0/OJ/hpKgvt4owNJ9+3F5i+6uaPHfVM1j/wH7Mz7AdFoMHCNno2qMN4kU
dH4zplsEAPOwmi5UvOz4wsHTQF2KKoWmqTqdH8fJ43j4JtJ+9zwNjNxm9OPaaNmsAgcC2fA4EaCf
7fuCGJaEdOhLoj/h2alThn4q1p4vxeBtxVor+1lHT036BXrY6Qs3qubmNRyFr5+UJ2jbBoHSpXmm
7yDK3lW3oOJK6yAO7lxvE8YJiG282bExPVfV5c13Hjg7SCH5i0K2A7r/goMzUHLr1RGQYJeOuHhc
MH96ClvtFI6raE9AnlLH8ZqRmy28e6OJbpOXrtyeTSz2TnBDehk21lp/uVe0KvUmmolmtwHg9cI5
2RuwRh+0Gnuw/MbclV4HppvFas+39l6SCxjfZgqTwgG1VMkneT8Bhk2nERTKl3aPgcBFCpi0WChI
75zJIKYECTCGTCQb3K6jkuWcOuRrEYW5AtSkRgaujLMao8JnzhP65pYob66oST0d6Hu20YEw29SP
ciJ2TqF9kQ5G/yv4U4peJbdXabKRfrmJ3Vndq8mo28E6HMWGMcqNy/UXq0Lh1rVYGjFa7SBYO4bz
CtzmMrQ5qTgRJ1Bj2cQam8CIejQlVM1wK0Pcrt5w3FDKjJTKNSkKwoTa9V0GrunJFKHx8u4+Cind
UsHNWMDF1FHlKxOCFY+a4lL7mYL8OHDlj/TeXQS6bBl5kaUY87Nr9RcZhK7MIbwDlAXCVYuqRYVv
8oXB+RxlBbgQaB33olhWKZFl1lbEyE/urnOxJi0EJSClWQrHQOMuXjs8d5EHKKdw8q9d8Rf1rkEt
GnMZJmtajp/q0XxnVm5blnb6n2TJA6xcDPo4HBYsfhbsVX7WmxddF+0RJazyMu+Nlrw1ZqgeKzki
1h8newTG5cuZGN8p8tL8Uu2Z4yu5CJDDeJJe3rz0+d3fOL348t3XespdJEWiUpULbMQYZaf9kwcI
Zy+Jm1iklKl1TRSlSRKd5bRoV5pZA64R5ASoITDUB/pqgWKGa/tRbcBQJE8jXD/AeFSmTn6ZpL/Z
ZXU1F9uM6pIqgw8IhjSCMF12pzLCPiLMMAcl5HQMcrV+jqfwQ9gTfBWiNmJm2RdLp80KzK++Ye5n
7qw1IvnRzPCVvb5OcOydbj38qwReViQwV9QX0NMZH/t1r5YGGYnyByEGBlyIZ3ctcuW2jA3OjC5I
TwkBhV5q1mKJlsVd+4tP+Kvh27ET/a9L/Bg6skSuhKOx/XRwzMo5BagOv4ugfCfoKHoOR9jaL2gh
Invvje7KDfwjMr/8huSih0ZHm8o3RKqMaMszr8kaK65MZQScm9+2z40sSqULzNSBhNk2fbhgb2OD
OGzsZg1ca6CKPEgfExKiBoNLXZcGPW9QgdPYrS4k/U/RqMV5okF6vnCbkE15MnkzPdGoQKkx6HCv
booRlDREGlJi0nuSy91dZPD4fcj/LddzNBoyM0X3MHR8v/MAI6Tr8bnxg4qW9IaI3AvyyrhE4nj5
6NCerIOGR+V1/ye/ZAp10hGj6nLEGrPKzUt5Fnm86adrYcR5jxwAIRjQMHwwSgW3vFxfquC3gBuU
FdIxDJM1u888k4rgfpPr5+Pk5xFCXLxbhEi0fY83PaYPkD9csyj+pSxf6Ieb6Uy6YdDyZnVVaYVY
kuJPw9VSlzpt27f4/J0DEtWzf7HM+0Kz9OthsL0RKcPmrOugWhRYO9D5NASOrF55h189hayoDIqA
HMFzfm3R+PZ1LO4FIWjrDRPtAhcU2UWw2PKCg3AeL8iTvscOHlfaSw6IN+vz40eLdNnKmbfWPnA6
aGgqPw8N4jVramLeBx8jHNvARz/YSP6hg9ZADwWl+vAiJamDXXCH5JGiCJiXVJidYJz9AgBXFQbK
ShLEL0DAk5gweyQaKA1QdyIXgpRmbmAKv4zliUoPHnetK5bXiMrPlteeOSTjEzo006kaG4aIm7Bo
Xq15DBsIqK5ASnC5PnttB6Y6VJXXv3dzR9MNl0o2nqnKRN0giXNB6Qv9KXl8JJ9iVHQGOlRs6ErE
utjlMzbtkI5znPWh0sf33IiJlMIM7fYpJPWrKMTQzAXGZDwmh9SfJm2fEKw33Qz6oSak5l5ZDC5d
6gbi8P0OxBv9LyhY0d7fzv3GAxgt30CkhmT1EqevEOmQYGRiGWYqqSaEJcqLxabL3ejAyGb+5E5t
6gFrCS56PphI1tuU4OjLFhdom9ZatEM/dU02HeUsfI63ohCwUawOxRDK1ciLK4ziD+fM8Y5/9Y72
DSHCSLEs6nzTqIaUuB9IBQBaU2SLbakUGzQa4fF5dyNmpOI7yblYKOE5tapRps4ZjwR7fvqR+SLW
/BxO37V/CI0z0+usvoq/25o9E5eYxQThFqMWyA+8RoGDRf8iOzGWVWhyZegs8M6SpqnPPeFPW29r
O6BntkbSQvVgWhbGrOd3uhdDaU0BJHWl1bz8kUQv08OmlVDFaEgFS6jsStqKwOG3q8QwKHXY+Q1g
BzE3+pWIBsgL73Ipwii9PcSmjNxQjqH6vf4ETVfgskWtTAsoTXlDkpBqgZZ57dllhwmMyf9I3GsZ
6NOUadGSV7ff9Izx2JsM4RYWAO+mY+scwdysOpffaXsCEim4wdpPDxpYNdjad50DPCzW8sgDMf1v
RB4aavYx50mCl+rujbKMzo51x4OqT/R7+rZegUQR+GNVGf281HHwVH79fpChIdU7mV2STtQXf5Lr
ptelQGEfpfZL7WUJFjdmWSTMdfNzk7tobxoUbya/zVF4bW3sqNKxcx36fXGpbOfnbow8c42J7/dO
BkfmYUcqTBWsDHL/FQU2VKqH9FPMonSCoduAOzV/OquDbFCuqbe8DBp5iwKZDlwCeDQqEKplsEYF
JWPG25FhAal7S+PoyzeqiIoYmdOu9tVij/M5aN0suT/aC7N5Mdsjjha129q+ZHj7mYUOdjbTAM9o
ruXJnJYMzuUq7KDnqcTt6nhAgIs9muG8MG6NcpnMAMRrKXxI1804dGQ2o747pHAkfJoD8l6oidgV
JtukUXLPlIgMNAvBR+DDixtXr/9imtabTSWVcTJVtBxM0i5No/CGnsZHP4y7Ds141wyFWOds+npi
BMVX9c/qpACOzQ03uYhpeWPAP25C/wg8eJR07YjzuqeSsgG1fBpb9Gaimuz4Z/hn5zQHcJJGrC9T
pucVJHTxotglqOKygLUETAVSJoY4tK5vVhwQiAaE53lxAZDshtWx5iTIrKawm5uHm/znUPOocIcb
B4PNQb53YoNBpOSVxrPF6AaDFfAclyD3VEbFKZphIOVx1TPogBmIjDn/cyif3YRafE/Po7jpfwNe
zcpVdktzCAtCNF+jcBfc6kUiOKeJJZZZDGIIUK7zxo9mGGQC6Bc+DLeo1YbmPCWN18HCTUvcbTzi
QnUiMDCltK69tMLq4fIsTUZbyQz+GBY5D7jhQa0pOJSMnsFE5MOu1X0fuwZ08fybcmdyzRfD+XO8
qXm6HqZ+MRzmBAMK5R8P2quRk7kWMZe7WEObgN9hBTdDdHyZTheYuRoeI+oDQyiCJUN37PMgS8iz
/U9VZJccD3RWuRWAdYEZl8QxnTgWvHc628LCOey8tHr+GJzGswR05FiqQkQl4hIC84dP3WyndSAg
PcmZIyz5Nu3eOowD9NzeFbuJ3nWHWDMXVEwvJdoMzKuaS2ZE7ms0g83b2+BDt8zc5a0Naup9HyEW
YVpVRV+bgK3nv4HgfGK+8NcSGa23ra4Hljqg2WZHF755oE8MeJDbO1NS5uS9H5j/WUmDNO2edDSq
sDkQGJC9On4mdqauzP8YI63QCkZzL3EHl5mpB4bQR0YgRNdd5JuxsPTGoTpiQdmOF0oh4D8829Ri
XYDDRLeNGvXUm2MaTUlJsbi6NTBfySHHMJP/eahZgZF4kAfugF/dKtFOnNKI4tISNsEiFfVLx6LQ
PeclYGsP8OeTrelLgDx5llOXLpxBTybdlxQAHXbdiBH/XCD/M82AXxXEYwsGUxCEzIZDSEufQzKi
jkzLpcjcWH2RhVuSouMzc9R43VSASs7LWPvLbZf+UPKlK12kKj8dZRknGc2/zn/+vdIhi5hmHf4V
JrOqdw9BqS1IUZmABSyKEg3msrumADpaTpMstVBB8HuBjr6UXuC810hb1b73az2dcw5t8dz3FYRh
y8BA2z4esojdLK+kygUq3DzvtTs20HkFDP3d1o7SDle8bnA/QHQZYtlsb8BLSxL3bR6E50TVmoLj
H0mcyyjAFNsjwxM4nY2r2JKWdM2gZtkRQk+sel+4ybsLbjwdvOi85QmGxyqNuuzMn3JrJKmB3uOI
LGQHXmY59H8CV0yHX8wWSoIBm+0q+S4AENbWBftzvlRBBy0i78kHZpgfTZGccinyaqc9k7MGqCX/
UV2m2vq9K+K11YMNCmBrBSUH7gkS4RKrjGlWkXeQSPI2PdE4rPpcd/g/LJvXWHbkrxEwso+QklAn
nZSNcITDWdkLV28Bz1Utwzk5GbKYKXxibnPhq/EEIqCKm++FbVEz4qq4KQMjhGohy/cKSSd8m+EY
smjO8hVO66zpv4AWwjvM0qpY2gTP+bV0BdAcomBi7C5gcNRguCjO5DSx2WCNH8f7kWtf6R6O7ZEw
wFRWunE122ZC9YDQ9in0g7QnmvUu5q3aTFXjDwSjlUicNbEenGVvu/ISHsOyTTrqJIcqGrija/u5
wbzRalLiUiunqzsqe9FdgKp068JY3jN5wP8isCxrQ6LgTrUPiRScm6atNk2FVa7/5FjRrerpKhVV
3PNEylC7S3ojVs395WNlKTlrCC6z4NZuoS19YNebQysofYFZ/2b7g15YIl5KBe60XGkQqwX8TZc8
gN4wkBWlcHxWGv16O7PplrIHq6zRGsza9ZYsxkd0JoiyrNzJ11bZhgDWrMpMM69Uz0UB9qp123uX
A7tUfW8NvCjOX8fuco9Zx+IGFd7Uhm/KLjpIYqpThhXmUOvqZ+N1SMcm5Yz73QJCL+cVabGC3bhV
PJ/oVlO0BLWsAuVvfCssGEjxa+W59d4YyHDe8gf5CGZ1gJ0cCSYr9ZbyHod9BzeM1NAke6ArdJXg
TBj+6mhFtLyurShWvQO3ZZevTONcgtwaGaGQ1NhGXU+FYJzTpvqUvn4awMsxhIaG4iTLrq5EaYHd
7+0NVhzU05/UAlRrzvp1OxBWCf4V6oPEdEe99cxtBMLSUa2KqRae+xJFxQOlo0d8UiGvFcpR16J4
BDxby2LpGTbTSs5ugDC2tQ+tUHQlqMhGcj4HrAR8RIhSwNUUgebmqGEyw0xMikh0d/lpPx1uEEM3
R307/59d36Hj1rFqOOCAqCN35zskBh+CouVH9qm0EVlv5g5SqocD2q/uyReOkNfpQBZOyrDy7x6s
yvqxpQynPtRno9a+xALYuzNUyv5V1lyXHMeFfU4yaH5i83NyfPUyLQiWfBzm/YeD+PFJv1soDghz
1xvyhTe+enQyAW8Gl7Ykh0c42M9fdHhusHB9kTiZ72rLFY4FVwNF17W6eXFjGbk2FPzdMShxO/rE
jhyp+xGY0Fb4K6lrrjj0M7F1IfplvLIiZdcHkOHHK6czWuKCfkSXW+PYO6pTB0OzyWtFaiXo9vo6
M4gDuRewhKF9dq6fMbOck0wLKSBUuKPJyCkKtBtkgGt2XjyDKjjNtF8xGOKP2DtZwcYhOfDUn0OM
23Ig7ZRqE3IAu+uWpfHUDPbqhjtY33R9sV41SLhyjUVjwRNmPhEhgMmz3DI2lafGBRTz1Xx5wCbO
C+l8u/E6Yzhbl3i5zqN3NW1iuwDn4B4cwgcf1f0y0aaBa12gRFH2qdiOJpyvRmDNR4EgPLfnz/WQ
bbfc3P1NyQHzN+uneOeBKBDgtOhtL5ks6blSZSqPKdwMRAkYFZif0N1x2C60/aPy3Gere31GzdQt
fktL25iiF51pG1l2l/rCrS+P5Nc1YFueHeF+VDyw9lTEot7u0NLiU7aS6Wr+xbZfWqH9Dj73a0u3
VAbRN4lQBjNxPB2ZThEPaxTBN8JAhduRzBe/7OkWmuO5Sx7KMfidMxenNBhVMC6q4ZSu5NvKouyX
tnukbSnzileoVMFHFaMUfRhf7cm4pwZXUBSoNP3iemtMlPiu3LBHElxSevRDB4t1Nqo8+9NQd8LE
ORQGPPKSBZj52u8+CgXi75SbLGomRm0UU4y0Bo66y9iQk+sW2V/C/RgqQhzRIXxCqA0grCU6OLyv
ioBsisoravQqxIrlf+w71+tkKlsHv1Xb9BwumkmSeyzy98zYJIHSF+TExxZg8YIJpfTZvtIbFSe0
hE6V4F4NIwLAv3I5lI8E4gAJhT2T/KpdB2YfIGG1poDarh7TFLBVsd1WfAj83qhVD+WmASQHNPqb
eXV9sKMfsQKgrcg95yd52gdAWFrE6XejalKK8nEQTL31rh5NE4FMsu/hfaf5qDFiEmepEKDLMce4
bboOe8oVLaQIXPd6OrLzlxRfxDB6yREdfI912Xkg435/g2ZDnnUPFj05WMwebCMxbjcbyT6+5l/J
QT++cZkzX2kbpaHuHyuJ0DNWIyZD3An/1oZLZbhHSaZwlpCa1ZUb7PveIpNgQ429yWvTrKHG/HXl
+wGRlm45zs/65/uxhf4TLO2MNC6rGrtr9/uWxvT8OXTSJpLehXk2mW84OUJTgsREluSTGPVF1ZOs
dmFpygrSOcAj9lHkuBc0wxyDRnj+rwHv1n26ScbQ4KTM4Z5JSINTDLKZbK1dYAQAB/csXhWRaw0T
jPLJcuW7MbLXs1T56QvOYRvFrf4MlXlqoMOWAoQzdKhMcRgAHaVYvPdAzJ4zEuztMtjOpEyD4Wta
vOkUu2kiG51IrJDkIpgKC8oczpoYZeLjRDtJfSx1rP/JoISoBluON5wRcrrzI09IpTR/0VmcVGiZ
4U+k9FpyVVZKrsgpWvmW5kfhoCs0AKQq8hnXjh09k3pd0VZlUAdm5ENSo7pIqKdg5sBpf4113dkY
pcSuE+74OC+hmuVY0BFTe33ogh9ZBR7rzTrgGjBLmPOC5lL4/l/75eyfE1DEB1Ceg65EPoKfCwB5
AknGMKplo2aZkTP0PxjAGEkNyzRb/Yw4i8McKx7MdyOYw+zOB7gtF2q+diy6MdlzBYyEC1XM0oOK
kuKsRg5GVqkWuBI461R5fI4vm8F+01jjupbJHxv2FdfHdZHylZrsFm6UGb1Og/Vru4wW2UWgW++b
yMjBBvR8HhAyLe5qNN44W5jl18ijuA9joiRKechGWi0WrffqxFjRTw/iIJWWLYpKcUQ1joeYQFFj
ORjBveM4EGBRY20uVDQjSY572GWNcARrtgWpX2suVcXAAypadx2qG94frR/WgQ1/7v/Kl8PWuvM8
m89/82x65uu+Emdhoj7CZaWaePbatlBqs1aUSszChVIDl6E3EW4yKYvAE8YrH16kZyK/bS/9+7qE
Lsu4GTx3q3RhfMGaaBUiJgkx2DnT0ihSEy541prBjq62DUJ8g62zvIvufTpbZLTKJZRdCgAuMDOj
NI1dWu2myUQtnO8u5WqnCzcoB0AGEnv13mIXWTZFx11Ih6Fpod/2+HjPBDxLpx9Ui1qQZv0ihlPu
4lpjGyvmjrwXb6QJziOIycqU4znaVrnOh7cqi6s63FN9SI5pW4Ik7/S+THuznuYa+ouzJ6BmY885
ibrLtVe/RyoJ11cx6tDcEy5HQK6H85iKgXnEMM44py6WUfE2xpEB7mVsh5Nmfj/qPzXPvegZbVGT
jvGeI/kn4int1rvS5Uuoei0UIuTq+FC3Tsh3WUlSnKRJbp42HBPChb57lRAOaalgqn7le5eAy6yg
8o2GMcS2/ghCcxZexw3xXeEop4g6uUGZrln+pRtCXP6xRZiPpPdMHZ/cZDj9gCaZOX2RexTrj6Y3
196Fv2a5uKSzog5/hMl2Tt2sLO84e1roQ6TACWShJd5lVQOzVdoWyCA4/Uz3BCBC2AkB7PF/wRV/
6IGP8WYzZMSZGaCZpF4qK0GXFix4b7f4wLLx9o62oPg1rPEj1WPgx/SqTAPfCX57HviTjrwvZVoq
BTFj+Qcln9jOifID2VuRgOA/FKIKsRiDWYrb0YKzLmFhdGhKy0AFman4j7TWNFonf6RIf+pJTA5f
YL6PfbHxCZdGhcUuNBGDnMPmEfdDuNjoTIkTh1hywyY5l+tLj4VVtcFJzxEZC9x9FbX0Fia36oVL
4NeieLoRAq1/iIQ5h7zvbVvIfxcz05YVPioNCng1iGlLNotTI2F0EElXe6RlvobY9+s/eybTW5H5
Z5jotdmlTl2jNqnwmKix/+8+GjwWQqq9wXYkwc2Jla5yNneQTdDtYucWBx0rCzp3hNAd24UJ222E
HmmWqHV5jvJrrnsdX2jB/lZgGXn+QqVzLJOY73S40qHuET708dGUHouSBag2PD3Jk6hgS2vEgx1y
Luh+T5Ved1sCBoSeKhJnBx+uWxkDnj1cCBiJ+nOE3OUQvXOSmXivYUZ4OIBdd1g3A1gFqn4rQfEG
jFaAysOqPKofi4ZhRxPymCdr3xh1F2UELaHWjwJE6+An29cC5qId/zCX51L+gGEVATrH3SAHJvhJ
izcLygKE+op1qKD3ebVn4JqevJdDGi8ce0xjAZGdGZkt7St38XTJgRlfNfZh45Dc4j+2rJFatKj/
Bybbzq1dlT55uPpsLuJSJxkGIAGafxhqP6GVwV7PaSZmL/yXwatHDsZ8oO+frCpAp/fH0VebIRE0
D2ob3Nl3bIuY1IhD+iKZ5Eu2fLwx7AWjmFH9ZYbCmfV6JBGJVFHcKZkDO8z3be3lDX3DN7kkji+G
t3sumWzMmnb1UR+v8OTZCFyfHdEnknbS5utroFsYPbukdG4Ctl+h0VlI4O3dOSq3/BZH2xhLRul7
514h226zEPZsMRBuwbPwb3yRiO2a395qyuhjIumU5YraaLXudyKcJAxvW9ASxMFD/wvsPavH2gHK
h3YuNtrtccsvsoyNqXQ//p3EysWBJX4DaXHuhyNaSJFq3i2fsciPnzDjNe2yJj0IK+OurLq8Kjyz
+hwZCpSodVNA2TqwN6eQ7Ts5PlKE8nefjfYKqhSikObIHv8LSqfalZNKTcMX2dOs9UHbe4q6afeA
lEw4vF0LZJtUB50xD7lM9+fmvJR22Tu/vDGZ6MYB00cWp6gDDG5vOPeVTdp7Qdqf54KcGio8ONNL
iasjpTN+HTTkUFlztDZZhyn1NU1wbEU9kjC8WKSqJ+THZh5IBm48XO+pi9uI/dn1OciymuNss0jV
NkQmm1hf9TQqASVG/c180ZANUPvw9FrgZDlucPfoB/im0JqLS/jpb/jdj2yt2HOVfnRi22Kq3Nm1
3C5LJG14/iK6a8T5/aJE9rc55Az2TTYGgSBcT0c264NWM3ct28Wwd6MOTBQiFTc4ZdTSFf59gIaU
aI0pYa3ijUeWhTu5JGMdeWrP2tsnqvBAvDfhHJpIC2D2DeLTmIxsSWLAkf6VibVe2DofJnse26ck
XFGHBRd1VmDfNyIOL9uM2q+1x7RbD+zFJFTRiKRI4PQFy2K6Bz37sNewq3QyVIs3J8auNUpLNZ8F
n3V3Q8iJwAyhGqKZKR6bFktwZV1mC+V/lAyR4BxEkSPjs3dYUrfMd75k3F/0ulcXLwNwIN3Hz7hJ
BjqK0WUGW6O0H2/mB8HLP9qZaRim2lPdCi8E2WG94uZrC2YQPk2FF5O8E8J65G+09UaUvEBrvtey
PM/DqLjXgMSmJLd8Hd+s56NJgC5Rm/546f2pUiNDb6B8OOsq/VIfPS0oIqXnczvpybFc8CfzZt3A
XhS/6Bhxwhtc8hxFHRuwwkNT8eJxvlYLnI+XCTIToqfhjdarivexM5dzZIvbc54LErYOtArFVje+
9y2Ga1vjnQdMvYlYZA4pMImGZ/eC6wQjHH0+uM1mgvlLfyddWiQ/1U6R2SqZQmVQdivTiqIVCTIe
uZ/Dm9ae+gv160+2Olm7YlQTvfVW37yHzjV6/uTdSMF3T0kAxzBHmwRPDWIRrBqcdMYHVX+IM5oG
z/AX49r38W89HFHbDl4x2SlZTbIiYzkSsjPkuSjv+KRbDsAb3V7ycuoGNA/lNEKynlrMJ02I9ReM
rr1EOKjn8ZDdui1QsfHt1V4a7T9bAAcbdXEjR6vEYWdDY4CnvHgd5h51Y7LH8z7RnWhiTAEHTMob
L3rU2hzWYt1tDGtoCyQkaOY9nKEyGkpsGwJvs1K7tvv7Cc9hf6WCAYKYnPCE7IwwUi4VHCmYLRIV
J9R6oPW4yLfCyzKi8LLjuLjFa1UtcXV6/MBAFeUyQ6zr939cZO1FLIFfZbTY483RBhWNjiatMxGN
NN35IaEc4CFsvThDCaB7JFFVo+rMLnURWyHNy2UqpT39UqzQ7UOvKoI/qlnhnr8X0SOAGzCF6l7Q
wnStE6KO++/RquKDq01WYSpRa8VAP+P3ZHKSjCUD7yQowQJ8vuvoXZy3sbcs2qlMs/79AGIK3Fyh
EmKAmqK/lYiB/5ouSwi1AvnArfRza4apVBNQVbkQQ5ZlH6lbgpQ07aFq0ER6MzNn9H5euzXMbFh/
NDNp+JIjVBA1wBYxRsYscpGRmCHTRT7SFraAYJRPERUWwukdzPa+DZ7cTc/7rkzduK11zpkYll6A
SWIZFQne0lloiRNuhrRfWDgRAzUZCQR1b3X0LIuWPj4JgxxB7s8BEIvOkyQqjIBVsXvh6YnNhDkn
0f8saQ7STEebOz4jGgneBtxFAxH+vQuaqsaAVVqyHdFgzzBkVFkeeC8c2KGr+arLrxme7w/Gvi/e
1e9ku5e4b1Rg4zdij3Ya+L9LBVimQdYWJ7lXabM8tPO51ypqfXaTRyE5INIcRwVw5D32Qk0wZQ+H
oAplsFe2q3ediSt4QRTe4hV00jibsl+3Pr4dIPf1d1E5MoiIYyMXeTP3WPenUfdjtOYhjWvRIVZ9
PodTTKPrQur9kp2LEW8NNxB3oDxmR7pYSnJzav8sMIhKFUfH5F5MTOWiNhv/G8hfuuLHL4n66tdd
5PCgcRKMQwK8mGu/eGrNCnPoQH7QSC+LDFqNg5203pm+1DtuWJjM+tZB/HQtYxw1Nfp0z10JOUeL
b4li3nVS5rFNg6GlBK3UkR8l0eauUJNwZ+qZTP9Yu6Jq5Y3sGT2/cFBHDUwkfJiRm8tx94eORB+H
+qXrXJknr18l/MHMWFqC7vdj/dggFDXQtdEjevtiE6XhfDaZ/o+W4iHUTYFF3nundoPPwCN9y0YT
xIGZGXJvsmLjCEYJoqXUGnUiIk6lwAEUzmhBQcQ9XCN5f/5QDBReM+elqQiB2m7sNc3wDpApdkj1
mHFv4i1g3WAkShkK315F9ySzY25cvWGzB3UcFV1kbwFDWz1cp8Vf447ONIgf7Yi8WQiuR++mOCDw
al1ZYlp+ex34glL6kuWGLOLpt2amybbi/KaPHeDBqP7LNbayp0uvV4T3NYdeH82tU07AM3EDqWOL
Mbmjn1E5UdY4iOF9VsBM90LnClEEYynI0iyt/0OYqxr/U67JRsVuQ+WBfz6Mv4ovhYoloHcDXZB3
GrxRGrsSB0Fk4Y3Z6hRNAK96DPSQXspea/1yHTuleiqbZYPoKalpYFAk1JEdAuCuCMR2pqBrsFq1
48xu5eCyVDJnZ6KX7xh4q+Jn4j/wew33chFQWvYRUJ9mADfPRoggUZj7e0Mb77Z0wouTShkKsPh8
K16heAk9LEsMrqJlYlMBBKZS/87t2Ca4KekOxc9jf2gA+vBajnVV/UEuOAEfKEOwNJw53SBsMWHX
nZSFTCd4X0c6RpWmsrOeA2DsC9irKrzET/fZZE0Dy4mqfUurR4N62mthl9byZwl1TjtWdSPW/E07
N+Pvyfg0kT5o8KsVQor/h8cLRtMIkAlSGdzhFVKoRG+ght3AL1j4IPhTOFY2BtjupuAF9tVFRCYU
cv8oCzn8dtDa40LJoPY5X4QNtV1TYnK8f1c0jvcky7C75A5J514N//FXvZmCxIlCIWtuHI/q/eoC
6rYXUQSUnZoSr3j/nKg/zwa+Y/aJrj0KTgsvE0L+fm7k/T3dPdF3vDud6f2QImvFbFJe3QYmSU34
SGfbRoV3EzWpNNmqMWEGlBAdfjkC274PnwTZCmjFKsRyaiTxCccnoOL0GeliAibx5Fe3thfD/9KG
Wmw+tSecUblZl9hda5Gx/+j5fMfCGST4x3ppp/iU5K3PqpwCwVrljXZjLe6mYOqEDyJr/pp6mqRo
I2g+hbPRPMGhUyBjXCz9ULkfllsXoV6+pP85ofq6Vy/hx4qwyk9AtWaob+0hokTZmUuRfMii1ucV
mD9dXqtL7C5DUMLxBcTrYfADxzHKqEEsdNuyWukBACLoAxSjIH201Lahm6D3gqKs1zWOfCMNWRRV
43fJXJo8M8S2+hgRbHNUjKX6fQP7oFrkSIjsiIEZ2E0YAMOm56FqTwdTxk+QYt1n2/K9U3CSTpBS
P/uMJxFgX1rXZGT2FDqKZYvKDI01ENz8kMbSf+2gzagv3gjKB4QmcILzY815LJajR4e81coNpDNc
7OdUQxQC6o8YCla3C7gzX0PTizx6ajGlWEbzFdIKQvWgsHgqSSALBYI0+1CXT0gmNPOfJJz61DBx
A2z3tI9ueMHUmNCibQSD83Ilj73NN4TkLBT6UxzcaLfnvug9iifq4L2cveyLwYXynshTGmBg+xRV
bnR4b3gyHD+pSuP0qYub2+Z26gXgHL2+61VV/xPFEfP8Gvy2VFOY/4KCsmuWMvwmh7A9G/LELuJi
NTBl+3PDn29vdnrko9y+XLB8TeYjqKkuc2Ja74kc0xguqVLLunhITzpbywYabebaxjf4d+O/E4VY
KKA9cGRt5valHM+31Eheu2hq/jPktMl2imRMWXipRlhbnFcw5ON0KjhFMdzJs6luAYb44bbKkGoe
YxoCGyy/PRajHG/f3xoiG+DI32XiWt7o5E3rZEjYr4fXsqjfpLHGFUzQKOeI4VNy+URXWMbNbv8d
FpQfr31+rTWdsK8OtMfD5GsxdCGoSMpTx9KxJBnywKow0RL0kWfcnsCT51omDCHP5t//IWD3Yfub
xvTBvNEHc7ACu7KpPcBNhggGSUTOZgZwpA6tzvAXoXu+p5JBW0tPEtMYZkCogil5gOTX1f46SwTs
xr9QxEvCm4NvfEyh0vAaNBL/IPfYE4htqFKdOmSC2CGQWT82FMvuKGCefi0jreljxwfkwlxGdeLb
sdnPfmP12fV+f9pJxBKAIHPNztNm54CQzXlgyahU6mrmDnO6QcYe68QnHGzATvYSRNCp7kQovNEb
Xmx1g8K2pasUJ8cj5Op5yZaPT5cv8r/Vt70GbcfsiecPSLYO/nie6tXRNNGQDnGTV0i5qwQZ+Yh3
15a+xivVmmZRxG4MHQglyW0As5PshJ54WOhXjxtic+DSJ9a8cN2sO9KZ8d3EWZkNJZA4pOh3LMj6
ZgueZEktcCaW07P67GDFxIxsEBJSivPREgoijT3ROfalsvKvJo3+5XZ+dX5DtnARl74X1R8F5Vav
OEOY62BLGHjkGGGAP5RV0ZUHMMgk4xx0Pu86rfzwImrTIILSdLMKjhQnVjkWewyflo+6g3NK0e0l
Kc2JkACbtwmFFwJXXT0oqm+NxBCOCklYOWUAgy07xtGeYJmSB5xaEPZ2fynnI++DEbYaCVMM7DQn
Wr7JOT7/bTGPwHN8g0uS07CgRwU61RXZnZLOn7GpZ2s15QERmShFj9FYYFMWydc7Iaqda/qQ40bu
KoZnrxwTz4ZEu9Wc4rjCxmW6H4kS34nZyx68ntIykWT+yEcRoBeGxa1mR8z1xXCJKtWYCQBGph8Y
iq6e891YHAj22ScrcKo4dLlFUyVEpW3O5fXOvhF9aN3F4UIYs2lLdq+w0Icllml0/xb4l0krgISG
3GsxJk9Tddhjsw2Heqzpyrw70HNmb12lxzlyzf629T7lqnBq3z1pLP8IsnybtuUoS20m3k+JTCLb
iJG9Jg+B1bA4WPIgZfCDXz2e6ujCoqee9jcqm9s9jfooCadH85rYDZgBlL+6O+29xp6Y3TM6NCTD
rMwcWebzbGoAygzCjkAGmusW1HHxbY5zNm+mtsGeH4T/hgrsc8WX/TTEmzApDuVVecF6Pp0abLLT
JoGAfe/1l/n0+lckPYBSBKlE5tmlj+WpU8dfzcfQWi50DT8Z3Ke+jZHN2UkTa46diIqTpcSQgXRQ
Z6Cf/YVUsdm6TxOrqiumqw90QOa96IT2WVZz31uqcyW/xKfMq5r5e6W3nYxfqlt8puN9OMh71/2w
4nZ+mSfTmWwJ32h0jNZDV+w4eFyb+xjUx5JQ5q9wZUY0zKrL8vB0vdONaZ5JpXl9IiOkgfszs9ba
cRnulCaP+yrwQ1BG1hacbt2EJD/aRNbul7SESkWX0IVgU9VCFnKRccMzVt6Ze+q6TX/R27cEB5il
iuwyn/l1XoY6LxjS7DKo87ZdOYBcVzHfjc8FoZtNhyGqzOgB2iuVqiLfmD8O73qr0m6sUj0RM50R
mdInPJ+NlmqufKEhfySiV/4PnjO1imQzHzeP5StMYHIXkKxJyfRek3jDIUckZHUHazCEJ0OhtSs4
ZmjSjSWSC2e8CxMuSIPxcbinGi3245Y6CQzJv3n9l4VbRWxJK6q4kiEYRjuh/s6l1DTyVMPyXjhr
4/S1M6pezsiEnSr1w4LMI2vx+ZQpwuKCqG+L2PY2nCRUq08Dq5Qq3Hj20pHWwg4M+Ost2E4qyEFC
Fd+NEqA89p8/AFXZLI/IISGmqYH81bViE9mRKTOKYhOOEFzr/pYx+toGRwn5MQ6HrS2bgc/t7Ikm
3oD4QCorFIlT2z3aLiQyV/yZZHAW8DLl8CEEhh1RVbftviSYk7gyyfE3tI8uB5VhflYOvIccKQTE
EOwlnVxf/DSktt6wdTr3ArxwEkEgsP2Dggj8F7CbEynmXkTJ170wfGnCgMIQv9w/r0RS4O5rGMC6
UzjQ2AN6lDnR5ydBbTsBdCzXHnH3j5HXMB6EcA5C5TIusC57TyA+pXihpGL5+ULQfHUDAG/WAJYY
ctzFgUWGKcJFOb1eNtu4vf1KuoOE8zL86G5IUyUyIaACp5/v72Y5nSRnVv9Jo292aVhNgIQDPmp7
Y3aEpzFY5ya4twC0BLM5m3MUSldvvZvsGwMMhRQCMaBBoZxcz9210WTSVBP+MCP/oVXRxjB/6y/x
9rM2pVajnZT+ALp9NIiti8TUocd6k+vuGfnIDrrRKjdGUWYAkqPBMLB0BOpMgUYUsifK5TL1Gg31
eT1VU423QDJ3vAz9FpVEDbkw9ud04if5dvMNnW+rcP/H5+8NRJRaut2GW8gF1ZusjKqhFFihnylJ
7+H/Kjf66mCkxZJW3Vb6skH7mVGS71hkg/pqLxQJNgLxS4uWL3mRtuXDtVk0dPgo5mE69gFcjzZ8
E4SbnxzOqUpfPg/NOyHn7RdGP2+gu9sIWC0LvOwPZYEpPQeZM4e01vQsqmAf09TCl1S9GisdnG2y
VNbtoJ2GlwuAAB9El4JMrGT7xvdt9iB1yEyjlNeUlnSwsN5kwT9D+XgyGg7za3XVdnMmcGKceD0X
IZi31LgqHCh+7h1/KgakmLaAhaw2vxmhIS542f5JDaKPvePV4NkdVenCi+fbQ7+IX2RT96FdUiGS
1Di55ohadzZtQjHgBrunheZNKGwly1NXbROK9S+kdGz25HUQAH/uVnc/QUq+QBjVHpqA9ZohbD6W
uCe5eBxgdG6A/1nc3zb91Vpe7dZHeyFOBH9VX8pNijrO0G2miJIV+h/cjSRQ48Nk4QFMHkuMZqWF
EztrRyjOeQ9+TDEoBXpheaYo75sfyGMzLBmvVG/nnOyJObp3+GVgeYhEqED4PJT7Ii9nU9YdnL8Y
uRgF+WarNV/1N0kNmMJdANU5ETaiqlRXumzXs2sILU1Une0xE1gQhDJMgvXO8EASUkt1E+Crp/xL
ZDVqiyMtSVAmDf0pNTb9vPvKZlL0gU8fpW7z+71+AZeZ9Ajd5oYr5rfuR5K7TTreCFKgy2CGhn2L
I4DUE88vPQRSr6SDUW7dOrUMjV2EbedMp3o4DJly3y1BYwCwIE/SlFhKhrs61Fb7aMAyrQ0sd6Oj
5tRyPkShHoy1XPPXhtdzNcxjDVB8xgsHyLbwGRPdjIQk8oqpoLYTVZD1T1oaFTvy13VxmDCmEvYT
E4D/8U7zvmLb3E6bvjqyJsBfT+bVS9GSkKgNkIwjRP3AFnafTdzw3rJoWmdAzHVYzAEOHSQ5iEyB
WNVvW3oINLdgx4vYWouTIDmnaqTfM8vFWG/4JTdw76QNcAzVQp8sT10cEfbO0NQXiS/9sihNeKgK
e5v+hMj/gWkVxXUMdd2hFhexmo1xAdTOcVQmQlqd0xkA2NGqXpK6FCrwDQvxBRkBWJCOdPwzFUV1
XiW36bChEERmuVTN5ibSh0o0sd3U70EI4LpoS07E2vyTCSjbFcl3wn55ZRpmT4HW9Q6NXCI+2l3p
16uOcM5lnWA25gxWycJBP40q6rlVQ9K0jaXk0OsQR28J8o4Zocv8R8yfRNhcTSwk1xsoCtqND7BD
YJdxeUxKu+HzkL2Ur2t/f1e3UjUoSK68PUczFicBtK7K9B6HdGGJLZrhJ5D+QxVtwuK5IYj1ziSz
Vi8l0r0LKfwbPgI1CvA3p1IA8GNAX8eQPNzmmszxef60vVrfuSxh7lR/TkWC2aOcK55H6dt0oDk7
7xeLkVjQ/iRIb6taCPwrpbeOCP4+W2CMImsY0uw/aspN4vR34FZ8SHJ3Wb2ts1JtW9Gv6ORlSyZL
v0aPVuh6QeXfnivu7n/HLf3fhK/Gw36rMtEfs/giox0ulmStEZqgr2Ind0ZBuZAK09kLpZI2gyAX
9QBzMT83SMNSnBT/A88Qz3h5HlHoRkqTafZPGk0ISriR13DQtYCCwnR/19/h16FAlP+mVP7rD7sl
W/RVh8n4/U5Dt+hZ+EiwcYOjCJG3mJyaphPYywiH3N17p83ArV117rxfMJCZDJv51IT/Xge5abAo
TkS8ctv9l1QYIsluI/DLblfaeTjC3Zi2vkKrXQg9vJ+bEViO4YMVr1gDFrSFWZznP9n722NmOiHR
85cUtUJx92c96t7r9rOCgv1SSUoxprx307NnnTQgYvi20h0Y0qYAS8iUVO2ZPESdbLpSx7X1HgIV
CeDt+dcFRxyPJLBl4PZk+LmpfMhjJ+W0ewfcF7ppR+AkEXupDYF0KmeP0Xic2QX28eKkgL5vqqaH
TeW4fZXnXmlznrue9HOyKg/3hP7hwPUS925VN1ru/7IRSZpGnyiHW+roCbDjuNzlmhGFBnlXnKqE
zH2WSg8DeeBL5y1G4zmebS7kexzdu7GOu0NkOSC8X9xswPGCOBhWTG7xKWRIdTK7JysyK+QAaAof
TVMSPJqOm1Ya4l3zssQFHfOqxVWjWOL5CqlQa4VS3rWoBcVyxeHXjSbb6eF5/NcY/MljCpNBgva5
lpqnXPPQdXpI+53Ad7W0mgY0FFRq58d8ekln9RLaX608y5C65fIJd2GERFJLgr2bUh7lrsydl0xH
sZvtoJBQwAnQD6ZsHoOJ9l5HB+LjiMH5Fk5joVQ6mzyA6O2m9GUurp9UtLi91pp6kY50ChN1BDl9
9iDZWfegQf7phKFEkcHJ/7aF2OEEnL3VRDRfrDSTjTH3CbrSycTBenGL58dT+v+oB4R08fWlbAHc
KlvcBYoBIsjOU1ALyfB5jektPfj6zf/WIewAUuETQPv8LUMWfDQtsPEpdBeYiAJNi4vmCfNPgXuN
iwwRKTek3aN4B9Ig+xpEdpurf5BJOpfIJ1CAN5T3E3lNvhnEKvIAJBPuRuHlC4IEgxxFY4ZpF0xT
/adDOFi0dMS1JbQmYNoo/CNDj5YtdzxvbG4umvZx6zwQqiiv06XfZ2rubShpWmekjwYIlFWkCIy3
DLONzTAPoSqCsHWEVYid264Utabbz4GffeZl3yMx4p/pF+mkVichO4jCUlaQ9msZ57zmh4LKiEv0
HKpv31tG+NhVw7qzMI4EGoviPZ5G/3YkCFps/8qsO3QGnZV/QhuzrZ4yHrD0O+oX/1zAK3UxhFxA
VCAblDDO+/wOuIJgg/BfWz3qk+LW8/lZUAIVHzbGEUCLqtDPaSvvhCaZPuoaxkljue0OlGhLQ9hv
A26xT2YHCuHkzU5PLNpw13ZaK1Y6nuhdFi01g5cQeOVB2I2pjpWPI4CIKTJzpH27GFNKvCS0SrM9
2wFbCSDBpPLp0LtpnPinVzz8m068HwUAwVqLBKrGwD+HHa0FntaC3iyfOb+ixvwP1GTKM4x/T17U
HqbVywSraLlXu6T96x6IzgR44YC/zg7PLL6j2tzYTL9bbOOHw6xKDo8mtnWcXO9osK0Eoqa8O1sN
mF9hYWb1/yW+eT3W4hPxPep4sL00fDswq2wuYzPvcAp0zds5RCWwyH2+ajDOorc1h8LAn/1eRgnB
7tInfuLV/8M7wM0eefHXduAagpQ86EG/yEaZmyAr7Ci0NDyfH48hrA9zHOV4aGZGEU5oUL9Nx9x8
SbYNFN1njhjtG9azisVINXDpVJv8CkA9LeOWZvqALzxhqtdcCteQO55tTr1vzvRS4Smo8tvO9s7W
jT/3Tf6GAU5uLi0le5Srb3l/pzcSePQow5SyYYb47SPedXR3ecAxejacdFokeOx0XZIzEpj9Bbnp
lvSLVHjSm5imYl+t513kLblRCu3cn+DaJ0a+AUgKvJad0ED/KIR+TISgrazSOZmIZdxOSRd+YxyE
UrbnKMfFvAShTTwwh0V2RiCF9jv76SI8QYsQKJgRY4ipVwOtPF5DqIX07Ibo079uas4mdeAqZyZo
Ckz93uwhw3nh1Hf/BLnMHDg0G2Nt0cM/hG2kTED40LNpMP+fpQml3BOHVZFlMpSOY0RCtM9bBPEj
NsLQveEJKvF6xoj/Xz+mFIFPymZxr0WzX6KxT3tZ8dCxFxHzTXmkaogAVe9AbawRSaXH+5+Z71zs
95HruLxvsGS0LvOh3azlYF9nP65bYiQEoAa9xvDWlTbGfatWdCOAyzZEZW/cf7xLFhZj4KLd6wzM
UOdbS3owPXYmHUNlv2GUnFKZN7HxsBvjb7VvSBIftYx3bdNw+K/7WJf4+FTTnWMC4dr87JPvW2+p
YXTfEaonnUf61t3G2KZGoXcFj1cHDuMhlFaEE57cx5v2YQJPMUFS8Rb4Veoz1ckQFuiCQyx7J1X2
/ou1Yi2j/KXzEO6XvPt5OiGrCZMAr4HMG/XZsaDdgn+fQj0Icqrb4lU8yRYMJpC7CXHuS3A1oqGE
rUfgqE4Ni40ZcohJsWT9uElotEatCTFdY5pGtlkYx/i27HO4KyIE3qJAWbln8WtGpW5qnVSpHWgy
3ONDS5g5QLtuSqob3E8WRTur3pqMdx5FSbtRi3Odm5gHQwtkNLRwBxuW09rfZ13R5JuD7KbuIpOe
c/3SLLnDGIvE9Xy40YmIaK3N0EIUFjnY8rBIgjWYahQ8rSkpQ8N584viO3ymJ+KTbPsBputb6scr
RPxdtBAGb5AD2FiO1p5Wox/IpCO+fLUVPJhcD4L6vTCtXWjnartYP9M4YWnpL+wHhwrtO48Yn6/w
b4fqc04BVZZ/xErolJvEiLq6naa4+0Q1wT/s71MLRfBAwld7rJJDeUbHV9Nay/+eqgwXg03KY9I5
bVwyTiitiNZXLHk7JAPrc/EbDna/J1biC+iMG0j1lxM1Nx0SupSgHA4VPSzicIgzYBUX2c3kIApF
4kB8GIcQEuzrCUAqAc3DcH2XjfROmdMY5/uvrVER2gbx1mzJYc8OTfgJAlLyKkZWjQNVramnZ89Q
Gpexkkr5iyB0Te6kM8ZDLy1qmf1FvsknWWoY/SyN7pWchM7dld8jrofVd8eeH+uB425qiPnEC91/
W8DbemuzssDXfAXvVuzL4uVame9CTx1iAPZpvyc52Edskqs7SMBWdDei92GAyVvVidsDe03+7yp/
7T4Jm88btECvazOT79ecmDNfqE/qS8ditNFyCyOaS4kfMU3ZQwuc3CE8Cc51ixAuXYwuXjazq/9J
8jb63h9vL8E9IRJnjSJg2/Z4LXfNnlvylyvNmSv0Qo5HbfHIjUaidTgYntBNp98sQArj4rKb5YAZ
O+hZ/CgDDSv9kUuZ87/rrteEaHd5NagWD++1ohOUYe459e4NgjJloK4QHJ65hf07sDoOg3vTMOrp
0vhxsvQ2TRApKcTSbyXuVOkAYRwCkL+fjtr0jXt+AQtBLh1+3rPJymXaCHRVgJoavaxIvYeMf+M4
IBV7BMQtGPzyn8mAdmvCTS0faQDdAq5dIbDUbV8OMhNpIczdqbEjJhkQBkS/LwhQsoDKAo+oZHdD
gKv50JEMJyW/GYtUQWTNBY9uMYBlhe377ruJZwEFZv3B/E7dutqCAiwU2T+K+gW63W/ctq+hbsos
yPA2OHcgqgUtAlpkNypTkna8WS/nBRmv4k5afkibeFNtbHSEZ/aXV1U8W1srvIkLubJeMFRcZNDM
64Yd+pgXWlmIsLARR/ApLxFv9NtTvLdwPcZ1Vymsg1zZcg8X2NOuI1pmjJOXQ2kVhzP7Ys8og5zI
I1r2Bqu8XEk7xT4iN8oOqaDFm2wWCxuYaofW6NKM3mSkkAqETfw8YQY+aTRXQD8l1Sh+mmlcNuGz
RV2CK9ntWSqXsTFCoXvTSMvaTtmJMaWZWtCZ48xgl6WDSlh1tAhtdTgIh9wOonv37pwagKfe7ZIM
7rh1jZb31BeE2BQYpGh1hyjMpEAhEVeXSYENLZLG2kOB5PRXuHCJpnsC7i+50BUkzGWDsiZmApIU
tVO8Z038zv+n73ie0p5IHmGxMduSj7RUvihHl7+veuDwxPD6VUbigCVsYSlYdSeSjn2GgDeq96aJ
ad/lWie3Kgi2jTJWwn7r5MIxd3sw5r2VB5uCORVi4DNxslGciZja/hUCa7aUe/iuw1ClmG/Qc4hM
0OmkLWYkB2fBUkpLfdMoLjHvyXdes1mzBQ6QA2RhgUqokZEuMweW/zmtXQHZp9U0EjKeNxNGOgbV
JbXNXKsRscVOePabEneGAUx72vGYuJWOCGcblwJOexQ0arKerr+ZlPMJTPtVsUURvAVDtQkUuBeT
WHRflKe0cer8bm7k16cw2AR9BBzBU2wx2BCxHd/h+e2WV1XrsjmXBdMdEQerTUfeSM4b5tcZ0MgY
uGoxrTj3aS5wB49/P6KJ3jdrdIt63t7ZEUQ7b8+BeZB/8Gu3DljpokIgsApzaIX05+iXOEmumVjT
mlIBrH5PU1tVr34ttuF1acVlbW5fyDzf9U/PiVc64k9CQRvezozd3Io9l611fE3lRdhG+2JJGhpM
hUqjLzFSdC0wQnR14JMs4lIERFETF0KDI30A9JeVIAf85Jk/zWEZT6oZKyVEPfUAHfg9iXlOTRA6
lIdu+lsyrX29nMbdTCH6DwzCZjcMVsce1GCjd5TnLHRVLBJHihkYEvx3zefLKyuZb+nThLjdS1RG
CaiMNmC+tUWacBJfwJ2eWAszVPnmxYMudeHMwehgCFGgeXMqCFcdTxTb0coLZEOLE/f5lL5k+iN4
w3sWvxZlONcrfNdWaVT1L+hb3S8d66DaacWRJl47hziMgxGbJNPzlzLUDXGb1811LmvTamG/mVl2
HPEWmcI3uB5BD4QvTr7GtfBZm5zuKOhFlN7c3HxmrYMkDVI/eC1NSAN6PXwnDi1Lh8p+ugoN5xf1
7lw9EMhWOozs201poRVzsDQOQ8ENuYlTcSDqnipdecEZW6eeXK1lQ7UMkahFMjxcU7KORP87XD8S
vIkYRRyGGNkEMfUt6q6yoz2q3Mxe6vIN8DlYHE//I/gaJwZytDkzsRRrprgLkPnsYu1XXYRbQeW3
spriQlD9Y09OuWOXgJDhfEyTaE9vxRzaX/st8XUvO8V9USgjV4lQLsswvVXUabtlAJFYYw6uzGaF
4Lg3RkeFtVqJbA8wWtKGQgiKVCq3zQAfZ3doWSKMXuKIbA7RZevEdOTG92Ynn8M5dx4r9Xpvxd5Z
357knxeQUWAA/oXyZYePHxb1IaIAD/UI98oLNFNyvOUcvd3wFPV4Iw2dVlcqp46SNMn/K8oeKcxL
1hxqyiDrm3oU+460LFl3baYNngM/04lIxD4wo1R5+RojrZoWvzDkZTF3GvZlNMbepAhnVNYKMLh9
uNBrB0scEcAaWVhEFdKQJSByyfYnVttwuWhQ7mVfJ9rZxbIXrEKn5/gOfRyuenbaMZDjFRJWpILX
gqVAc1D7AwTfDA1+rrVA37eMAF9HmSIwDTfvjFSsqBel0AZfP5Dz4jS7KRVHh+xYjm7KCwy9CX/M
MN4ZiykruETQS9zr8iv8HNM4H62AqKl9Jt0UW3bhWocNOZxb3kcbRbRIoayGaSbVESyiRH938Kfa
5+Jao74HidTO1Ruhht3xBXv4MNVIt1+TU5kjzgOwidobgoQep7jD4LubsvOamH9p3wyL69fPuTKT
3gFZrZ6yyC7B19mS+1slsbkRmJ3ZXrELnQo1CpirzbDi3HX3sFNmtrpC83Dcu7C06AScdZV+ZO0R
7YUmCtbKpdpkj+ZjMtWVgww9jHdL2zG56WxlfnWw06MkAvgsjoi5f4nM4MdXvW/zKQuG7ig6zITr
4MudPgmEd/uF92h11jaI3aABItmHmhf2QAddYkBDKDlE6dnSlkqE35m1dOKvkUpw1hSrlL3JliEl
IcXjq6kbInWGIEo7J1o8N6TzBCjI2hDNzYDCfRwX8xRBDPv5tUN5Q82Ri4uFU8o+foojBpXowdSt
bw1ThuJni36M0y2+GU3ps32X98YCF97OBIQuC7qTi+SHG9J8XGTtcQhBJKMb3WiopYDP5bUcUCG2
A2GEq6zUpTt9WQQR7NTSdX5hO5RqExBfk9dcijELMtqndEQVzZmyP3gHpDznmc9Kgnf0b7u0QNTV
z3gf/VEMu/8wsuVIG6lMQG1sgTcNH9hmzAqXfbKVOsf2HGJYncbwsTNICphiuz6FQk69rkoTjbaM
ejDzn5XyVnSzc1WxHhfY3+AEPNl+e0KtciKWH71piTFfV+AiHVE/pa4MIw27ORzPK9zB7RGbuRhq
03M/LJPPG0mdBKr11hiVUwZVBiLdVgIYZdNDFvj6sGAcZwxGsWSiw7LtW0CM7r5apz5PCDk6H6Cb
Y2NAvvJ/B4KuTYWnQjqHMKAd1yWKSgaxVFmYmqVF0i4l32erX8tCoWCEqSzTCHn+/wSS5c6HuC/u
LRv7HBF4Mbp/NlP/ixEjRCLIrkNFLMjiEEmNZ1P3tTdPqZGkC2MT8qqV5jjtfc/lZU8qnu8H/4Lu
/yYCQuNoqo/O65QxAXjNHiAa6rpxPRq8Dpb9Gsm27KUmV/PZP4SA0q6nyUAW9mBuRBWSMcI7hqtf
ZBydYC7ubeb6Wj4/STNyF5+6QPRHuNXHAkh1CICDmO6/a4ekxjWvZrZDQO+PKeTfoSxII7pbOxpB
L7lfLkqwcr/5Yi3rvOuoCbHPzKLSpFhzK/WwF3hOr5E9a79yaw8HPuJafC/gDRfH67mJ+1vQ3RFo
q2ciSog2sTEZnS0eWgo0Hye7dqgyrWgvUKy9m+uQzG5INxEGlmLG2DlZE0jMKfJKefg89Y0Gjcsq
oYJbXMjHtgBDxL4A4xVp0cUNHfQuC0vDA6sxY2qBVebWLUv+oKSVWmRUbSbbiUzkr3kUduq04tdL
BeSmbdtfaK7MIQp6Z5+IZfc6WH5nPKpiJxXUcg4ExyEFF+Ee3yVIsZkVOjq5FJRgPtrKSVsjmTQR
E8elluN2lQmLjrIHyAvmibXHH3mzgGzREA8h1+0bptBHynVELyfabs/Jg8D7nZ0TYnvY3UP/PfPs
K6D4TF5RVpTtTpwnaUlOXVumt8U2iWUCdLAJKo3A/ldsJFLAYlrGmFpZZ4O6eHbnxcIBFqTiWNdz
Cxs9MnsVHn2qjyaQExm1EBGwFu3FXh5/NJTqVNYuNsczfVpC/flW/Mo+hVLz4vqFxkhw5EHtSqZS
4Gsa1gkpYaficc2YjHB4wBu5WWCAkv/ZZ748xAnvMzsliQinigEsICxFhlN5NBOqyaKpHImid/5+
Ca1PFAKYVaWwQ47Gi5dARK3YSDhaAJauJs/oExA1tZWMlkq3xHgoEO+mRyrGk4JFcWMOONhNfLzh
syzw1MIunzlnP2DtIs2x+5HJ9LjkW8tOZ/xT8dn70eFm624t4F/oCPBLwGnuxmQmo+f2y2EJCXk0
ngPpIl/D2ay7TOEvb/az8xqyvwW9dbEO0VaECRk20kIzPuLJ3yp5fzFJDaMEm1OdL0owi9n0l7ye
NfvR6c4zN8SDfXrjPgKcviZZpmSiUfGLoUaSKHsvjZs+cCuEV6NFeMTuGfK+AuWkVNUe0Cj0/bSh
AEiBW9j9MNQ3F4ulgV44ynz5rl40NCltfe9Er8lQXspSRtLFKkU9dtx0rRxDyBFwk6nIyUhjCDWd
ov1BH3GE5gVEUxujp/0lB8T7oYTm86LJv81ySGa/OZbDe81O/lvaCGVW1DZA5zgvVCYiGYRCpyKs
Kfq7mcAOieydofttlU/Oxh2467+rMFzPWvxctz3Andm1JzQu0LhOMXD+yH3X0Gq4NMpGYhg9ul4/
x+fWZmnFIhWPT/xMbcvT9VtnEitwy0tKwUDBWvW7KwTmqUf0pbzony/0m0rCX8kVMBaFU2kl0cFI
7/VVUzXC/pyrn0qjW+8d5b2HReCAFB05RQ/GYVCT3oFhI3cSrvqeOQsnTGR3by1armyv8TPpV+Ow
3lPbIa+yCZKEn7eNo5bh5mo6pL/b01e8+mh2I55V5WdmbEOLg1lJO/7scHoQClOSvULxg7yvTZ6S
D7BC1sNccZrPpzHt7E/TLUmjv1Lx1HjncNO76cyvUeT+03EvgGT8pJLdbwzfDMURm6RGikqskiz4
gTkDAEKg2WV39dRAQEThjlma5qk9iwUxNbr92Ry7AoMrQTGHDN0201S2D0fWDby0qN5FPEMVm+yK
axihZaXp01+wtnC68sfQ5u0KjzxB/3un3bajdYG7psmXLczQYEZnYgqyUBHXlb5s4oPFAAq7Ph0f
+Gk9YSr9HUOYhVHGmoTNEoU+7jmK7gx1VeqJ19pqgYO37cvnl9LiTuqQMBzSo6rBaCkXB0gsv62t
zm5siKp2EhbAC4dYNnhEuq3wnhQKNQGBLRp/ghj2g9UAELPITD+RGBXwjqV/qj6rA/gIq8Dt4OZk
B3h9fVOrQTVZVbO91KgzTXAzk29zatkYNJfsxmsTutyv/fInGAw1WbY07lF9qB6wZ8tsUX/BS0wN
z0goUPljGT0w9Rl8P7rIEbpus+rhMci6vH5pXclPv/gNYSe12dCp/BNXlrrX0y8ScDlyny2K67FR
6hPA/DUcufuHnU390m3gLolgt5IKiVSAHJ+698HP58SwvVvHz35CMTSxmVxtbtKkY6CfZl4x8WpM
/rZQwwx/V6C0amtfDv4M4J0+p8K+C1GE/9vJRHNBlKAop7kn5/2kEyluqEKU7zOazcxyITnPt0ad
GOpM3WbJEyBGZlHhsPjoSu7FHRbdFauR9FBWTxSoBinKvAAgXRyR9qvzuZ7s33dncPC83F/aph2w
gqT+is6YYNCWwJ97QlBplvMFp4d0YfwvISOJXcSToGOGqK2pvTLWuaTVkwIUpS2rljzM6EtUUw2M
Ga6xjFPxGyqet2lXO8yeVBIh+PFmiYHt8xKf1uKYM/DKDAkx6vdm0Pru6JnMEOmJER9j1nuQ4Bte
CL6PoyBd5wTd0n7VH0FwH2Cq1pkc/IIj3tVzY1/hIoGEZK5JdRYEXjUL/KNX5PrX/Y0RAI2EGn0Z
gBv3n5mf76E+ViYMNImriLBhR7EKF3I3R2iDBIlChRP3ZuHYefUTKRY5EA+M98qX89Has1Jwv0xy
CRiDDwVXqqyc9HTGv4nN58uj8VWHuIIkYsrK5wKMPbshab/itogp5Plr8cWIor5d0cwuph4BvfQd
vCKLR32VJqO3bDhfFn5RzIwREsqPKSsjRwmbylPYEvfJStebVs/hMkffbHC89Kkd42a2c9bxRq5g
iD7K9unyV8M+94hSQQ+BCoEMsN3xQudCctnWG6iVkbqxj6MNsR6nvxCaJ9yHdODSdDMpVo9nbquu
GlH7xCM8Ucznbm8S0Zl1szHJ0hd3js1M97GdxpDRpiNaQz4QaDUQX/1qN6iVkQf6EgN44HfjCwEQ
wQcK97iHdP4GEGa8gFtT4cyJaAIRzvgdpwH6HtK73tPsw0XaUim2tduj717tTm0aJvQb1J8FFtxY
DgZbBsZAf9aGUn0acOKdQLHwuob9xPnt6Aiv9KvnquglQ9mehpF9ZjGTJrJEjASCpKIqSxVhGDBL
QwjXmYfgTwi9HiFpLAPM5bM45uZ1wb/ZsAner0f9znO0rLHnoHK0ChExLXhmujYd1OMs13lZRdHf
TEj+rh7SZ8MZkyRpXYjieL5A7fgvkKxLhRpDLGvsMUN8pozuVKSC1Pl50jcrw1vNEot7lSPjxKlh
AJFzKWLJxcHBHKFv94inOipZGaUIf877ZBnglrYehBWDyo/MM6qP26P6k2JcGG5gHqUx6fywDLOp
h6GuIe9zrS1QtK9kvTDGZorOIOoh/n2+37OOD2VlnYnkzGQNZ0Ub5ouadongUlJc2OfBDeuKAjHC
DgnqLD8wgGYCQElR9CXkO07LT/E1uHNFEVvN/7TgLAhPlbq9ti2u9qhXmUvjmh+8GzRycQRNGv87
inJXawPrcqsTudxbkM29t4DRO88os3jLTDRGUuiODnOqW7HqcMFAWiOYL5CutxL5XZSb0V/exYSj
6XUhajco0zowXaUPCg+9U/LWyxUSrNvrILXRzRyVDt1hPELcKkjsXw/n2IcOfsJGSE97C/mvL/Sd
zDWX7Q2MPStPlbhldXHpaTCa7gmE2S6RNjTWOL8uBdarSUJicpfUYPs61Dji42WSFqjG0Sl7XAkT
V9hWxsXvAJ9Og04EonrRlpYh2+8qjtpLqy67/GR4UiVsTLb6mfRJOFCuExv9Og9GpAH0q9YGQodZ
6j297rTNtO7Q1ji4MSYxc+S+Q7Vv2l0vRzzD7ONaZyKclGXpYzQ/2KFjXF1D5npRuWhCQZSJFaSM
lRaJVSduKsqWX6GW5/gM/Ek+p9ueVECyWw2FTiZT2VrwcOxyTlMO7490h62aLIOE63YroFvO7YfB
r051qLW/hPlLeW43j+ISRenEgVRMw319cA9CVvSIBEmz1KCmIyi1qtNFxibXy5iFLtW8/ClM5peH
WkPuJjQUXk9fnKOrF3nCColP7Y5JWFtRWgf25tHvBjJEHEkU+0sOhUH4VkieGx3RT3+kXli2B3UR
LroqN4odjxa8RcGXTaVhtHYjxj0+okWRsl/7lI2kBY40U9jBDSfIj+2+WKlPVP9eKOcHNs31n2tZ
ljPt0gQzbsxoMMNQkbzX+sYVJao74gnwFKsFgZGDUtSJn44BgDLrPQoz/zVJqCTWgYRN3cWHpX/5
TVSlXD2AXTzD6C3MTpbLqr+80FnqjxoEJW2zmApRD3QNqxbJlNq7li0twxbGb1vLIhwFbpziFf5u
CatiG3OBd+Ve1kwAiLmjP6Zj9oPWFyKECMstn5kF3eOlxClXhDLy3xjtlul4SmKXmXmxfNIgLkMV
c1QM++X31Vlwema5cw0myj9z3h2Tixa7d/W0eQqyx/uM1L1ZajI5cOyKLn04QfiXrradEgubvrbb
llKdDI/n742UbBZKT4hT3JQyFymZcyC1Vf0bqMKjGGjMBkDxmg92/AQbaB+61yWQxJPBVRuML+fU
uGdM9ByfnTRp8TFQ3/R9q9rtpi5JrOqujPTqkh4+6yV748l2BZI7+3J/woPVAFKO+3ddxgUpw8sX
x8B1Dv8DrOmYkJyd07lRZZyHrVJX6b2oQL0Dz/xyXEaSvbLQbzT3dqu2rKqPb0/OCvOnApuGxuml
IINXKwFDkvN9iJtfTGY2E+fi5gXfHojvC6Uz82R9KcXTUZ4efk/cxbI6X1spa8I/fL/7KoYF0wg/
eZERW/cSkvVUqG8Ph7m7FA5uZLeuj8/glPKybx38I0+AOBJRPVAUCNjUIc3aaFjuHixFndDakFUa
ZpAfsdIAESyZzob1FESUs3gofvgI2YEZdaBuAUhQ3yVbbYfdX1uYncN+pgv3CWG5lqaPleutw9VE
d553H7HnOrff6YI9pTApr6dMk6ungBC85C3nQh0A+GIU6RM5rpdMpCda5gccKSZiBx0tatQ6x6sJ
j3N0AEALE6arbUWmyoZz0mRRJPgMA4cPrRYrrnbmVQYOpi5BLw2vpwjIiv9fNC4OyudDJNoMxZOZ
sEubSIBO6FyqxHB7gpFKheGhxtOTBgtPnib+Lh90b3k2rrfGlod3xSmnhfT7xc6UU0kjqAY8NOjt
/F77vJda6Tww2Txr8AY6VdFOm3UAGSnk+c9xIfQCiyCI8kyNRr75dLb9jWWrngpleu1nWnnZXpFu
dVRAkLuB2MAsrdK2se70vQgVejhJkKjyGcbW3pb3ZautavvTgshfFVFPLMyrnPUFUwAFGlhaqu45
TDowXvAH18/s2s5qImgamS2u4WmWAAtu/ETktwbnGj5pirkqovTXiOtFN3e91HXgTgO936CyB8bt
mR1HRY6cLctQ+CaSNN+UGxplcfH8nhabP9iNtcKM1IJw8rbR3545XHslvQPUy36ZoP3GSszO4z9p
WDi4JwV5pP48T35cUaYZIqNKQCSBLGKUzA06ZUXfcvRb+zp80yiqPdImOLZikGxxb0Yd8JV3jtmP
+nWokXukNGLMUOt9aa6YEVwD0xmeLa2fF46u8PNMiyNXfbAImP1n7ihoVQfv179qtbj++Qr0i6zr
HaHmuUFHk7pCsDpNZ0VyU7ZPHWkOrRDmgY84KF6QORgrAeOKAR+68PtE5/yTAU7P74X9FhXE0At+
yYcPREyn/nUg06vdGDJ9dfWw3UyP+/yJybuEdCgeneOQw/0fGF4/bzSFvNb5UhtTfKt9Wd1FdEcW
bBbgrqgDDWRajiUeYyDXr6WvpJC3f/oOQY/nT5TqYy1nraTh0jAu4YPlhnPsZFA4BURHqiAotKgb
jRqIjXCZgrqGlup1jhmMM3KQalYE/EASHb4mz+vosFbvKuJNIc8jQlE4Z60ZJDMoIL4mDnLHrAjD
1jY5x8DPELA783puGdJfCBvqISQvC8yIYsuzNEXc+CvU7cH+aOZY73+HDNv37oDVipfvd1Y5ErAa
I4i71eNwKicz1UqPqbCzTcNPH0kj49Cn/ZJqs3SM55w7QPzSlhzUWvwM5PWkJPVK0Fm4/VhxgPBI
atupyGWILK07FQDyZoRowZXFVkvo/e8+79QUEmR5cZRexBom18ijCPajSrAcUhwGUmumuBirXGlm
Cj3kteq1s8N6dsLn1vINzUFJGvGpQPOwrA2PsjnWyrqcRkiC5R9t/AAy+vOAYEHWp7C4SBZwHzfY
1ue/fVxHOplq6odMt8Hl5oj5TkCW+IAdqla8DB4Zoq6Vvx9Dgpu6QuFJqeXVOoXLS2ricj8C+Af7
j7VhQgZ5Uqhe/1iX2LC3SBY85cFcgqXN8JuE+sepKiXTI0Q8PmSLIc70zKVfZuKESLWkwjM4vifQ
LFhS/JIJ5ijjs/NIrOhcBMUE1FXuFD7tNCNYd90tonbF88599Ge9oa8yD02W1/Cv2O3GQfyWbFj/
AMybgfxO0MZh0pd7PZE5uH9IEM0oZq7RXDOH49LVd6P3AXhooHrN047rqsCxAd5noZ8tVlHO/uKo
uo2h3kCYvlIEDp3RqBffCi2UTn7YR19K6duG6ouqqMMNrxaBAG9lvUo7AGeyX1HzF5d1k2LAnEox
q4IrEXP4Kb/nOGMKjHX3yN3bewiVr9mt9Bp4b359tVYFQhphTHCu3ZQZoTXM6By/C3QLXZHb8a+A
Nw2BYQJ4UO/g8oXLIhBrJT6BCN5o7BhPNA6VDjkXXs0vkd0e5RPr6/YO90RU1nBKUGuiESDvaFpt
4Kz+gDNuegnPPXml38qNmHXCHnEfPLr3EzzQ3PZ5uFPWRuqyGTN21wYOljmsqdxJoGmC04Mz+Rp8
Awyl0Zcl+atKmXcxYZBh8jY9iaCzFYIpPze8IkYY6e1qEUadrrdKOieCNbQJCZ2kuxSaB9XEwahT
goP1r/5v86mDKt6bgSc4DEiynNCHTl/3waocjczo0FOtkGhZ8DIjK4gWRgS7mO853HZPMcTavzn9
IIjCmTr4ENZlMDz3R6n+c+ikEx8mHdLVWCBRn2i+j4JnMsisv40RgBaEUJUDWWe98uQYOgwJnd8b
x27lkyU3FLkKCKTCaSU+8V60bqQJbYl7uDpgcd0mOE+aL6ZUqX+bqwaaxNKj1hF+ASneOU4cscNG
vS1zmtX/XXDsGsQOvHUp/wtQuXbGzGSId/1zF/61hOIVlkWOjxNH7NuYPss31N7e3Wuh5yS+hMLE
DLGPJ7fkC1Wct9k834hkA7OAJObQas/9B2A7xGQw7ed4+epXe7HzzjL62wo71AJ4LW7DQAB9i0+9
/P7yI66cxWzzPLZB5raekGAJPoiIQBL0NaU8iJomnscUgUVZ0JMQ5a3r3/YvDfOiiLr1/nK+bxwQ
8dcIUXUn40Le6vbOk0wliBq20AN0mKAiJclhDKVKpPYNj5qEPhkpU7HAeBLqKM4FftAySqPfTTdN
4bx1VWk3bpxe0zcIK4TjdVmEV8fCIrhFeGm/MtcaauuL7/5741I+3LgglXN7nQTYtqL/eRgEVTV6
TiXqgKm4S2wm0cFG+CmEtVNdKSGKAvXvMmCVVn+pvHwdZXLm69DLsjeyC/cLHrv7obhXuCgMNlFW
ziaov1/4m7vWZxGPT5oEoO7wzvSn/Ub1vQRkCh+kphSHDgHL9FHapV1NZEeNJCg7hSLTKtnxyAAS
J2eJwUKdlKIZOPGFoYxeXJBcHxtRPlrNZ5Aj5oMokQ445liJ3z3EHI/Yx/KxnxuAukv3hbG27WQ1
yQWZKylHCCMjNROtf1pLhrDbCSmOMq/e041RcnrLXC+tXO92BOLQuOW56iah7z8jiBquzai/DxaC
p/Z+8oVjga7B25VbS+0gX/ZNsZNlvSgEpQkunM2rpszi7vgDxiQ7V1rdrsdgbeIlTgjXDJbp4XSP
TgLQsdYDcUkDUE5KAGkm0Puz3vl0Pu/ijRda4Vk5h+AEXLvq4iCBDRxVbY/cgL8fNwcozpZgGtX9
6YaktfJl8kBqUuMM97NvbMbqSSwvCTVaudcVfUKS25+Dq08OwTgXzbokZ0qC0eGueLvfUId01Qs2
WzuzKpNLbAJUOAKxZsW+sAlXCxnLwbNNHBB2pdNvKXcfx2BwPuIhcSeoavY3jvIcb2dw2ngC4Q+Q
vx8awD/e5rSxB0p2z3uxUHFm+fZt9r+3gLjah8NwCuJ75Esrw1pQ9JUwmqhDRZWFMbu9j4Wm4Doj
2+MXBV4GLZ3+urzPTw3zXJLnai+eaAMcgFfZDEMPhVBhJjFg+SvtyXouQ7veuUSgIQxnH2s9vmhw
UkXbBPFih/93mdMsFq90WuJ4vS2YmBXSNulDvvryPouE9plD4FMwUxdWjTXp03K0JeeU8Hz6J4wS
YTFidi0ZQ0YmuXu57Prdagtr0vH7eanQSO08JGRDw0Y2BQ8uzCe6JLoBtd0kojnJbHXURxZzMD+M
yUEyB3t0Osdo928AHAshZUJrltd+3Z2+C5Fdj9PyrHO7XLOjrAPg4WQOrvdBtTFDqMoAjHj7kwbG
pEAx9F7c4CkLXjUYXpICvVUJMSlJTqP3H/PZtMrrCBG0uXdC5nh8sLfUoh9JBJTv7JWmob3F4aEx
ZeUimA3aa/wNtZbg+8mzMexoFaGxJQA2NuHocrczw6ciY34YMf23n357c+JoBzJGZ84A+JLkVIs8
iNVwxdqiRb1Iv3BZJNUWyu9Q6uc5Ls3ZhUUgFmu//1ijDYoGyD+MU67egr+0oHbr4z9iSU+IlxII
bUjSyBOYlpu/KN7oXBDBxYxu/hNeJC/2HcTfxlR1OtWlhkuKcEwBQolbg0309f8J2uS7ruN7JwHT
kkXiM+81G8CwpaLDukqnEFEOBGHSdfld9QkwpjeAuw7nC1qrO3WYLpU7lsPlEQGlJafKlDACE/jy
kxPPtWJc3gNsDF5XZDaMTDJONQKw9qTs+QXr8VierbTKQYDC6DySlIxB2VoMUDQI1OEru4njypl3
FwuuCq66zy5siwPx/UfZBvBZ2OiM3BdOGqhmwh3CAh6zwnynIBrsLZFgK6rRza2pnKB+tfrbpcr6
nTZreor/P7EW7aBuBFEpkV7rMJS/Dk8t1DUjFiozkmckWLqKVwl9Cpo3vVNuHO4qVObt7mK+LNBT
qcT+CMoeABHX6pl+pOJr9+ljf0dOcMov6i9/2ChW/4hSMMpAFLza8Gf273s2PCV0g2lffyhCqqI3
rOuKMEgIPP4zVUbhOLEOvt6BjE6JWfKlACnxogbXuDwh9BhhyDpzkkbKZJfBlTfluf6w5Pco12ox
wZS5KgnClDzau1dZrUxezH3XaM8Sn5PZoVOj/T0XMXp9TrkpOJkEqVK6cPyhVAYkquvTXFkt7kmt
hJSqg6abMVoilgoFp7FzlfOkKGIo7hZBrrGXr2l6FzeEq9ZD7ACQa5gGKoPJAWxPO6zU8eXk9MAk
eJWmk4yxYDEdrZfsmrCDgq2jr84yfNLcii+0zJR5UVGvmDuj+AV914yh4qs6ieuRHlqtzO2/P8cS
Yt3peNyQw9aD5B/aOBsMuV0erKxUlLOFODdbMy0surDfz68BjIKBwiXWwWBPNlkrb/rY914pgIV8
vkagXo1FT/SBBWwWEe//zs3yfU6CY2V6VbbtD0XOL46OVcESk6ZtczqH1Yu5xS115yoO/+QYpJT2
4YK4Oq6NuPTu4ADxd+b7vw1ff+gxPCPeRo41ZGShqx6UdTrzxQq6qYNya1gut31FpNTq83ySu4XV
4MCbUH9A1Qzo42SftObs37Sga+IofpbNWAWRLQ2eCkTAN3bwrxTLOisTKVlK2vGpEUBZt5HrAoL3
tuCrey9iE9ZCHSmHTzRvsKEu1kvw0NazAsIMBTdksoPax/GAFTHMzL7fIxh75kWP5HTpx7d+0Ep6
2SovP2S5rjcl6qHQ20egDRDktCtfwcL00o8TeVvXizGEei72MBfbnXUmj19PP87s9FbJYs9JFE3D
dzBUTwdt0Wpgn0ki+3MSrM3+TFyTGJVJ2MKAtdZbcForrbsWSSzez+C7GQzuPTTNcyfhCbFd1cIu
RyHHGd6LljlkfeJ8OPSNlorGM5HG4V//VXm+XHijIrUocyz0t46nNYYrJnhLBwkhsJzlJp0KpPAo
Rf0MsneNLesVIZVERdmVZpp8+0sh2D/zdpJ4XsSxug2jJEyOQpZKXlWjnjAA51VfFXPKCnFi/eD8
iocYPWMJCsTJBM4nJVjEjbi6vpgaTh5LapNX/VgCqvelynBJ23IcKhIE1uAe/fwqMebU+Ps4jaC8
mDNuVqGVGuRGpJOE2MVE+ervPAk5RiOqHtxh6rlzvY6pyDabJFl0YYWd1lH63GRPwCqx6yOks7D7
RxEUQM4p+5wjlLBKwScoq3w4hJXXhcMLnaOc3iU0jyl2TueT5TIOlUP6N5IukAdnlT8PjBMKXQtB
jAPl24pgUikla1YEqMJQJkxhP2f3h5c8yocBtJ6TVC4LMFrBi/ti5Nnwzlokhv0hc7QEGP9nkQ83
WNZieW+F8MPALDvjeSyutHv3hpjS1FhQySijqiNCVXgv15QP3afl+o+ZpN9dU3msnWkb1zdzdKhh
EPbRXMu0za/wD2WtXsiyDSrnXGXiuHBimFd+Aqet4q5Y0Ty9Y1wbE+cnkhKamePClLPE5K68ZViT
Uwz8/eiBie6asc4bZSk9TI5BpzlIbPU3vuVoTRjs7G6d8HV0czBuPtOX03eVBOIaYs9Ksc8CVRLW
HQQb2meGyCGYGkSI/IYYl5zz/x96uJGNgh6SFd7KYyUWJzRvpZmaZvu224epwZvFEoWZSyMxhO7v
rdoNGs7peMFFOQvalTIEJ380dXlaXAghvWQNX9dAuKf+yQ7BCaJvcg/TGDgPFcWbrcS5DFGS3pPI
Ow1hYirGou9FSQZBNNkw1s/HktjJG9aE912cbLPIttlhYBLBaqfP/G4Le4PzHxXQJh8lZ10PNXxV
QIYUnGaM6q4t4VwgtoC2I3GmYwEaPxPHJPyCqAY1uSettAGfNED4wUEuFEum2e7xAnVKlWDczM2G
sSh+stNY6bl705XbDnWIMNHNrhAc3v7+8XaYUQMKrQkM9VXvu/mqajY/90s5H3Nn9lWkAJqeQFbq
elFICgHqW9rOz3or2kdTCqnSQP49zOj2oNPfUSjZebRKGulIGQdLzEcf1I8Qo3Y0uclVOSejMoM/
I75Xz8lvqY952l3xl++RZTUC6kgCkRccaGz7TyEQdHCiv/i/HPoMPZWytXytnZJyBKORp+B/staP
6kJR846jcJ4LpCbsgzC3Mb7qXiepmo++Oj/40VYzHyr3SUlPHzCsw73ej2vKX5u5TvbUWmgAr/JS
bDuBCUCABhShd/KUncUVpVjBANfPNtdgAnl0RbaBXDCcbtUPGdb2sy2FnEMmTY61kSVWrAQ6G8D1
wHH4lsNSQKFuDmreUuKJ10Tsw1XK8J8QSYdAK1+AP9daUdEWJkeh4MXoO3eZbHSvSUgfgz1xkhC0
ujG0obDUf3mcqota8oZPrzhFTT39Na+aeXdU8ZyjH+6JXVobEdmSca/SxHpA2hEpSFMlal4Im2d6
q2+2G/pXK77BmKktjsMc0k9cp4nFXtbGDDFe+nKh4iXvJvgsPd1/aKkCMeAp6ztXYk1UlFEsBtnu
vTgwyR5GTyJ8XbUV7f4gt888YF01fGZ18AWPqrpF5O0HaYurVCPseQupwEar2U7DVER+PYklSxIb
2oPe6V8t9rQf24Pl1r9z1lw/QUHmLzUEmjmEWqBwfTUaM8agfQXLMXMiRYQIrmADO0uq1KVRdpus
QgePeuf+lZ2JXDtjOtmI1vILV5FC8r5ea32YJpZIcc9FVoFt1trLrNFORL25uEJdacMq3IC/CCJs
HcyRmk2Sp7kf+Q2pDK3WX/l9zGyGeCQfuh6v+s4ZKXX/XDR0AgaYvlQoLA/8nM9f/4eZHAo9Ez6P
Xu7ZDzvFxTei2rx721OFsGKEgGUa3yUmAec8w8EQNDthEiY/+UeJ4Cr0FzwgwjfvM61wqEM2pegt
1B4yybwX7rmZPzu67FluNorHqG+bOZ8Ce4oLW6lXpIytHML4dzfa7oRgpfZgf0g07Wmxn+Fg9WrX
itIwl8gYw5ziCDYLg5lz5wgYmKkx95suSHtQ52diPrIzetlt8wqQfQ47aXFvHxudY5QoEkiLT50U
b1bQSyCRB7XHTNhhlFzpbfyPomg08owbwxkWgVcEZPut5gCLWGwIWKZdWU89pH4I8DrGTCbvtzTi
dHVMqJDrXfYFZzAExgBOINJUd0yKGNG275VSOVfnbNOeGrUv9SNOkZvfP34ivOwPGsAejBp8OCOK
+5i08ue9BB4FBXb3RPdhUm59yep7dOcocIOpPFqYMZbJCkI7ApR6mT3fDB0OgY9EfGZXfuLu/I3K
Ju1RyVzVoxbEzpl3gcjHDlrp/pK5iZMhrRir0gVcJ4uVq0YApfyzPfP+Kj0VZCW9W05gl8JUQ0IR
KMODaraYlckj1n0sqnNUavOnwrHi1+/MSPRZdtEhHmT5BHqVhMzdRgnn+e9ESx+TOJqYXJdR4s7B
Ommlg+1RkMOFQZ2hR7KOLbe9Tf+lC3LaEabBHq0i/rC8vO7ZPc/zT6uEuh9P5vTkot57L2pnDe1+
PSWhlPQpGNWeEFVxfPl74HmRYsTv4lpdeV4u7SfXFeQhKgUyLSEcbJiiffJ574IwZ+bt+G4R0qAG
Yk4tDNCp4q92kg8II86TMl3x7EpO55AeFIH0G2YOkDgaXSRtt+Mz9M3Qd0hMam1jbIj9x/Fl9Mf6
N0jyFmR19WpXD9/OHGfvZJdzaEqlbVCXWTvwRftnomaQXBLBGWyhoBhfcoPoRHGKp/RwleI8HkyM
GBU7CYqOR4Uhd2/2VmLuh8befLuqQH9u+79PW/ougFaJvuvNfEEVwlfKIp2ha4Z9OV6+gkIfEFDq
NVj7qDdEKXJeiBFQlv4JMJq/sd+TJzw9FXSTP5rrXGuCmelxAllR5nI1gNXtstSfpae6w8XNXSgg
dNQoDFVsYba/y17hKvTGfCRsdlnETgp+YQjM8M51QBmfJlfU8JYcUqv1zNXZBt4N/CiJkxPI94y7
ADSYa0MaSrPpw2udzXJjjSmkeNMV4T+CBoZfK5aNcIfy+xllTK/tRoLBKuI2pLkL4BwQf0YflZQq
E5JtsRAzm179OJmoollFGX7vxh8RYH7TaLOqrL/cltLImRmtJnUsPdJDj273XtMUhT/q/yJPIPfT
TlajdK9Dn+Zn94ihW/F6Q0aWHlnGRpyhOOQWBIeHjuvXhyQV8PdpNCH9DGm4A1F5bm1MxnL5N0qr
ob757n1NSDda96+efVCvWcFbUTdjqhfs4EstX6A5VG6nC8u6dDjH8wlwy/3eYT/1tP+qN+7nWOqA
GNGLOV94EI7OMK6ylS8umZbwx+z0KWAe8OR9+Wg2yRBiasGMIUqRBZyq/khvzenfaYDxYL2/OLkt
JSthPKH8Li0NGgWiNfUAjimIzJbrb4zSNy68KtzSdJl0lYK2YZlrZ8KD3bQuOo9ywCDaiTYQ4+2u
zAFatCXdpRpwJEAN0wxuzJgvWJq1Fhj2Ne5qgSQHE9WRcblz8xWpbuR+2GJGF9RxwYZqHYe4UDNo
ukmEva1mSqt8uTzhWCTT3ph++1E0wjn2X3YDEV4jf0tpn2l3rDf4bPa0ZikGM/SR/shFy+WSTMdR
lV1N8lVQ4VP8b6g2fhpmWeV0mGivL++DIDdvnrbwQpaLNCfT1T6p4cqczg4IrPba4N4TisfBIhPQ
Y4owgyYj5rUvsrJgODri2bsdiGnw0QmZGHSR6NeMOPFEwTiSdLCNa3gbbk2BV4mejAB/+lnPhhQc
tKQHsdGMnx2fDRplUboIrTCi0mjoXN0/fzW0Z4eiBNSMKqqwY/16pHw9Lusu/zVz+Z3DtqtiN9R9
PUEFPlycaXzlYcGxbPZZs63NMve0ITJ1RRg+4Iv9et88o+2u3DdbfgavXr3qPj/jrJuFmXSkJjn+
u5LwUWbYjwJiWMTumlo3Mx2nllY+6KGMh08g86jmSrwAUsvbvYqvtfJ2GCDEdgVYeUkowXDb4J0O
JW0fdb74zLmeb1rSeVIr/k1Nsphzq1UUdOXmXlW9HXiCM/5tOmeFmhbktp2WxtOyy3Co6h7KeH11
OrUqDN3yEbMJa1umI8FJnjB3RtKiKy5JNXj0pQHGy8oq8dtcoTKzd8ERkyNC2bujVxiQazbg2cZw
4LQuVa2OlKR2XLv/8kywGzl0B46lyUhfoxlzoJaICH4Mx6EMYTQYpUd6ffSS3xc1ImrejQkhjxmU
ksVQ9RkXaHUINm44Cf3dsWag9e+yDZBu0p68yx4L9cmEPx6CDywGQlvVfS1oSCRj19CTp9+jOCsp
XCFu0LD7f3u91+mPOqf8e524xjMl6SVEl44AtYartpU63CDUaMXo30meqs6AwZSWQI7olzKkxqGT
8/f81gOsNCac6hISaSWEi5O1y58mxo6XNLOGDY9s59JdsatjZOD1Uy8vkF2Gn034esO00K+930C2
ScdNjXZepzFFwhLF8uK+GanbJ4N8zWmvDKOOhjL5aUDrwP/PXZ7om6eCCX9XVA/AVyfTdf6XAItJ
6TE5phrJRj7JFyzCg3zMcuMoZxu/QVyG5+WFMigaXQOjOXGbmXYjOJ51r1S6DCtlbnbXXXV8kAgP
p0IKMAeXT+axz8IjvOsHyD2WQk2EF6I2n8fympbAazcbX80JibpL7aSsM5nT0wXAI4l1O5eiFCmH
9jZ43ARgh2WUKTdlpLP+FTMjjxshlhKbpJd/vzPHfLIkO7IICBzqeG/TaxjcXKyV+owZURuCwOL8
dJeJP2G5+YR2fSPNNLBAfjoDXky46qPZJvV81jAV94hFSp2u2VvdptJlNQn6doAkIBo59bsECFvv
F5zTjnyl0QqGMyKnVN7Km2616o2XzXsqF1U+j0i1xL12o88X/+bpyY4uLPK2EktQFCflTTQJbJW4
2aYdp4fBqHqESYNWVka3bVcDcocoWShB2Hr6rvs1NDdvZmEDzUr5ZbFzhETACK9IP8hoJ2gqIC5n
8m5kVWuQ7TAUDc6nmla8UVYh0KXT+QX/M3T/eaBRsL21Hzzq6nYpRY9tNGMZnHnYSx4wNXgTqCzE
Ace4LgCz3S6SwJGkgoyqBSovsqyFJztG8hudI3Nnd0aTgZ8/RRMhPNAEyybYu8tmmbqAghh+HU6h
NS3PYhhDqX3BOlW7jmLcTgDJ58HRvdaLPuA8947d61Noaqw1CR1UV7YyjgyDGlSYfdMy0Z+oGoM8
KU/QBmThZbmIe6t8VCTQyiAtj1nW5u7W5WjuTVy3yXOlE4Qp1giEhc71728cCrgNk5VF40X9oyZ1
OuuS/AA0KtSIQsCopxPZ3s8/kXsjR/PnEOtffk3650bh3XEOBCFfpxZEjEeRHZZz4R+EVDPFY4XF
Emtl1uRtE19HxsYrEmG2cLcaJs8RjhQ8Z30IVwR8M3+BBYYg0XyJzUOBhkpcnjTnWzDJFDtzM8Yd
StTVqCSZcIdHhqnQqYIpVhcP0sOwvsghpbn9aRACspU8gOhE2hm0gRTZw7ZAZSkz6xDdwAED8FBi
V0KdLmJYNr+ctQRYzzZJs8Cx3jNPi9jOVijjqfMiTprxeU7WnqCUyfMknFT7NevLvIZ/VfbGM9S1
GudCP5j7I2mEcauOWyEY5DkxtjvS/LtvVPVyHZvVHizkn8WRyHdZv9MC8FXWv4ogucygXMXYQtmW
/K9y6YetVyXlIAmHQE2wT14ZjW1TJDMdVutqFSMHclOT7oHzTBok1jBxtVMmNBIhjy1/doUYPbZU
M2HHPrVKeSnttxsdHn1/9/ltKTTD9PjJsf+wErpt2X14dNkIUCkMrwJsxLAH0aMnSZeS51LqNJ/F
KmbGPHbE67OD23H0sq8v3cSmqzXzjrNhPsY8ytM4ijRnc6YKLNAyURWVwt/BvORqv0pRWxdl5Yie
xxtHhgB8bAmzR0cYt9V+dT5SjgLjQ1gmsF5XvjwT13mA1gHtdsICDHBg317yp8cxhBn4E0q8D1qF
zDhfze9NtHtsXvpptoeTzjnbZAeXsEnd6EuhTbABeWLgmYoVIXBXjVpKFdPLdH63kMyyAZRq6wlo
zDoTcKgUmIWbuJHApCzrR/sEk/0gpqZSZf5uyhW+yq1Sz8gzZatAuW9wJZXt/pFHce8FKpNbgzua
m8qcT9A+xqDrQRHvbOIpeAaz1w6FZg3GGn6dvdjRy0MxVXsTKhRG/cChO7GJIQjueNvP2A/2iW88
B2lthugAtrIs6zshjK8eIk8mJJnp1HbszjY/VMwZxvy/vgkoqNObBfRmhliNAFUEtYxj4mDrV+in
YO++wjWIOHoz6hQD/EaMiOlaHylioez8/R+W00iG3OfbyMJcy1jw9s9fjBEy1SSu90IzVBOnZUh8
88ZMKDStMTbJAeOl/+JhOP7mp6AGYrZO+C4Naes3BnpOpfe6gEdT+H29sT2FJrjGL8n8EhwHkFlu
U/6/e6uCWI11rAdtEQH+WIsNCWMsUnm0SE4/JRVHOZUOT+PFmFiF6wNp8zOKtKkF4oF2lyf6hgvM
nOzHVYt94p19Oa3CRKmdINhqdHXi/jNjupj3YRs0XEOpq/nGyA3cVVIk9cj2K0DFrpUBt5KzJUPa
2hD7SvxRo7G7s4mvPls81S2sqXTdGursehYX/MnjspneQDjaayBw3P6aTsTAKZcu1l8tyODTB+9z
gqcQeP8/hlbBJMM+im57Aa3K4KhyRhZpnwn3a9K9le6kW52LOtyQpIUmBjRPZtF3ELdwvZp0N56r
cCogc26Lha6JbWX50btYotDwD5uPKtyZl3gxpw2zwuZqiMYhS4onCqLGD8vbl8XOP9ZRkLBtEMD4
lQWQULg09DBXsqIzfL75x2/jg7BqQaCEgLmjukWVyYOq2ZOzNXy8z2pjoJ/8jNwaMSSKLO3lOlgb
WGrFFfDwrb+F9V3LeptgVgRtNG3bL9RNGtSUFEDsa0lf7vRA4xdK6zFs3WtOe092paSJXHAQvKLu
5EyrALsKCEooI+4QHxVXGXmd0g7k6B3voKkL2qeC+WHqRGhAp+XIkJ+pgYZ90VX8KFHPaNUHpxB4
EHpQqmAIH5zl2HMFkKli/sfNBDtlJHUdZd6Vc6sIapxmO0+VmcSnn4tRT7xr+AD/iZpRDyXZRuyE
ZYZxZMmXs0pcjRNMQf83/aQAqcJShfr0+CLIU3b4C29tl5nVGk615yxIv7TPqHcWdDbsw0utN8eI
WK56DeSjwtXnuYSWyMcjU5bdL1ovvV4SS+4tRFZY8dZPFE51qj/lFZuyoX6XcpEEV4A9m0c/vjtY
kZWxWvhb7J6F+VnEyW7kGZzFnlQmdhVziGVd513En/AlNa1mAW+O01/DN5sgR9whHWo64N4doCYA
dAUOGKLOwJklheHpc62ULkt3zrBNYnADuIzqF6k6xBNlviB+JiBB0CTTSIQv/JMw8BrKSGjszsfk
DzI8uEAGunr5KMgvMZxf4IHjC0fj0afizCJB4YDFkzRBeN1ZxR+h1xwlHzCgUxv7aFO1AwvXIp+c
8M/CANVa75G4TNLysYecmzFqWleEpB9PJ5UBb5m7pLTKqfx5zd3jSfiZEY2XGsPOr1rxL57mAxfz
Uc3p08gj7EMwO1PaqRSAYnxUkvTlcTHSYmx1dKwFqgmPkjjCTo7Ru+F6zmn+cBktA0w684uaQrEJ
B1Rq9QzZ8h2LhetWAIostd1nEsQWcGvqvAuktpyB97uacvVrnwskxU3z7qFGcTEBmvIrSAfHQPkw
C+3Vp7mSAnZrGl9h9X4kdi49GOa0IZwZOea39i1Sa3PK/xmrnndZLTGUsFvTADbEqZQT0sCOlbz5
mkaOjN8uEztqlKS3hJLomHXW2hDBJcuLw2Edbk4IJ6MFss/iBJC6C92gbayo6VZ6eIw3nWWCps1q
qDiSb3F84QNnZO9hDgJBMyoRG2qq5UrBrF+99tDbYpzLTg5Spg8lof6aKNjeegmDxwlbYTXBPKgD
a1nRB/Jqu1oy9VwNd4cAVLcGkIVyIHHnNNxVnAAVFKJjqk6MAjfk3iN/ftFucQzB6/sjFCuXFKEz
IhrVFSSxhxOuLTyFRVUzaJBgmnCmd7bilB4/nbbcSJ8fDJW+2OL88icuJRxBBdAqIsdp5mMVya1K
DudbLzRykZVyE2E8M2rMh4o8Mz/ogWXUb8icRIrUR6+PMZ+igzz9edfUFMLnjSk3Fp2f4/IC0frc
AAYU0rO39NsmwOX3FLx7oyNppvP8/PVEurUqErejWFh9+dfsr9kOiReq9WiPGVc2WGHRw+B0rBAY
RUqwuIZykIpCyr/da1SJRSH87GX/p120X47p0x0w4IVCDbR11gt3RJaRXSanRzf3yK0eO1HgzNnY
t0ar9BDDMQK4Nv4zyzOa2c/634R/BrBlJE46Mhni9W+EZkfk3Zbu/shrQuMzTf17pKHmyeMEQOQy
Qn1Ymp6K4kOrzl3YKpCDLqzk2PU40IH+plvbXJptoOgAWlGeL5dAfLNRG1FM779HGbC1PPSVw/sK
leV6xWr0FaASbZK/Yoi4bplkvr7zRSfrtJArEb4UOBfzau0NQVdvun/tIdrUoznwo5q3g1qmJ5a1
Lx32swtblFzM9aruSIfzqXdrNLHX8/lOqd4fYov47mFNSddoS2ZKfA/hiT/65GQtpw8bBhFP7Rzf
sUTzncB1J6kZ1TATb10jUpWT2S+B4MWd0hpTQNdBCOnwNl/kHFRD9pBmcqJjTXqYhP170ktrvmg6
4dtDiWJKOZSxW9X38HPx3iCDpjbj5hwHCqwpX0TzPbmzn0EzHW53sbslf9BXlJg0FoRch9KBV7GH
DW81L6mk1au2iA+3TAAdy+ixAxpyI4uP0cKM0G3FwE/P0NYdayZ+3fC/yW9nlusovp8lYxTV66a8
ulR/jqoP711qgcd971NCzS0URSPCz6XC5Np+P7cyrIWGELHBUmx1k5c2PX201ntUxyuTXXhcgS1Y
SCWI+2HjewblerLlbqXPDPO+bvznehRLPcwLP9QNK0V88RaruYLI0Jh5kYIMRKpXgmyUjU4rOEHt
OokmxANa7MQvriduFG4We0PCzuY/GfwxsOfxRVvumtu6ujpaGeRWCrCG/Gt98T8RECN7LeH570ll
H9HeiNfPO+FvS8S1dtB3TA2GCYYUrsYIrLmxQb1rps2vDYQoDNW3iDggdqORer32OAyu6awD4jTS
TyUYN+LoDQskHBhU6N4pG4gYbSTQgUqK2VmRz1Ffn4Y9JbFXnYmqF+hsZdPFbMoMRvJHeueNJUks
hEB1+wDdHm+vw76jlfOcmiDaUv91YyichkYGdfcMefAQmCbFJl8gKHv28fGeV4vAdIJXzgmjUdxZ
Oxb80pHhJN1UBRxYcIa8ExAr/Ml+7IntSqf012GW7TiMsQSP4XSzViKKnnPJodFuJEVoKeLRhF4g
D02abXN4N+OSbw83YbhsZGD1GRLpKTPzYkw+mbQJQOxkNF4kHh1WpTImbtbIjKVaE0GDut81phlN
9Oth8GUlCIU7r+m7mbSDhlrQkcsZYnTzMfaaNXiOg1MNiypm7DQRTu4gdzp9uUDFckAULldYDF08
nYJyA3EQ3UMaQDqH4lwhCITE0Ek/zq+6Suy9GjlScI4B0XX7mVqHfb4cRnZKVXttSPKcHwI1w536
oMRSm3zkeCIa5c4aJdgaOwL8Ki3IooqOC/oN+Z/Glgwe9vQH+kF91ic1g80wIDfvMYqv3r3TX6cM
kj2Gz1HXgCX9IQi9RvctiFiCKDlwri1xMBBMbPUx/4cObKL8WzQY+ZqEEgwvRDrGWLqbvpTcRoiR
jnay8bafspaFElTzobdyVdenzvelGYouOGmPwLSPxayn0VU8IvT9aRJdWqWR/UKy4JYjTuC3rukZ
+fY+QplASz5oKop4XACbjVUyS3qIfFI0d+RjF7hsSy18Shc0WjP9VPATGs+dMa/73yxdSJJPckL5
3MRamihUcQu9yQhcAUUAzIf5SEk6qW3WnCVmTVRKJvrz06TDyEU61KRt/e6NB7mqNYsnW0B1JR56
XanBUqFERqRVAXd/FibDXy/oD9iPm6pYXY1yicjgcxSoKTLltEX+/ZSU3OHJgczRN9+6nFGdIe89
mVDnnNT/RKSeWl4iQCv6sPz9vm9ejbTCmctwP9eXakOHX4q6HMDi3bahicEx+HSlHidYlhm8gSq3
88G9Mi8v4oV4AvranrpSItYXFOW5NyL4V+K8LRn/q6I4hw1lGn4B7wFMXtVqW13eNOTVjuxQ+LPn
9V8tc+/1r0d2oZId8meND0oDMCingK//n3oQ8Gl0sQ/AVe/7soxso3XG27thpqaZTihnV0vh0wJl
0QVx4kFR7vnXDpJ3BunXe6Qkk0kSW0uCv7/MfQCMIzj823sO2pehwVgZsbU0bNAsX1MPUPvHMZEs
e+EXs5XgzH1/7yKiRwPslQ1nAm+NWrQEUrIOnIk3aF8hZnvD/+nBwalQ5oCaCTn7Qxr7IKJpsu/W
llAx2ck7iYVcu/mEji3G5+1Ciz76APAV3wuXoWSS3OhaXB6aj/BHae8iO/OCMRBENC/Q9tm2WeBX
u7MUTyUGZeWKYVPwhxPJRdycCjKdWCR6yU6ox/2Qb9Wxti15HAwONP2A8gv6VgTa4aE2/U722mCy
COaSleP5ECAiIndqB6DuO7Z9jDo1E09vpWMAvZMTooI1gQObI0LkVdHFkUYIKb+N4EJQo89g39x/
r1wWw2I969uatihGFVKVsh8zy89gQj/nkVGo6WRBT6krsbBqvfSjnSbOKG1plaiU957/G8bdN2P2
VRI4YToOlEuiywlQgegrqM6UrEtqcEv6qh/fK6Rz/AwVQYuGJtRD4q8YdfRRNwgH2dhkyuzEyv+1
z8aMG8hYR8vKBmOe1mAgvmwStUAAp4gtr/01WNWAm4j549u4Xf5ihFNU6HasrR4AbvkuzBgW0C3y
MBZmb4y9In3GelfbvDpz4lGCCQ2cKA5l4Cn9lgnLaeFJjWPPQFEVGxI7BlV3rToZu49XMdaLM8L1
n7Tl65sVwyEyQkHEptHiuaSdkUCJ+3/4dUDOOG7C/79tLXffI3BTiNYw7nIkoHv4vY7RF11lhrFq
m34uWZGdco+6yxIxk9MQOQHWNtK5GKIm63LZ/yJaeKfSbKvItkdrM8OYCYHqGnEVlrzDfYVumHTP
wKPq6DPzi7D4JBil7RDjWUEug4qc2JZSto65u4GjyjN8E7IS3z+M2npsengrzfFHmQ/dwwbZ5LbM
20MAln0AMbjmat/vldsT6VZXHAaZkx2i7ZoOSgJQS8+JM4edvnkz1srzOUNQMxlaZz+7rzKAegc2
WEU2HHEtOA4HF78MDXSs5m+Cz7Coqbshl3UDJZXaoZlQe5t0RqRPm/NdHhEyI1ElsDHUcalvJYCx
Y6H0/Sf6ldehrrIDLPHMmDtcXJHqJi5OlOSJRyAi8UWoLy1sVkXhPt3o/Ci0CYxB6IFjqGVaTlL3
QtZDqa9K/KRLyBi1Kt+f+knOmkIKYQNCtFyNc7OkwN765F41dByzwlKmUJ1gnTqQ1uf5oYFLv2Bp
ZE0Hnb+2WA2p3szvTK/WP0bRH3JIh2eEsjJ+q7k/MT2wOoE1NiPIHUbun9m9XqpJUoEArlWsG6Pl
sG4Ui75Mc2vK48K6ne5s/b8+mwMKZZxDgDe7Kvc0zdLtnubQR8IrybZ4bclpkL2XuiA3Ndnjf0JU
hGFqq+8IBN+n/mAfvTSdyg5V2n68rW4gqBxJZw49AL4VxzJaodDPNDA/w+UYhnMuWbnZofWabtee
/IH7SltqrB5IshcZ/87a3NqMEIKj1cXO+WuOl+0bxnu/U9MEk/I4WiHgGcvD2YNZHcBXGlxALktF
cPoUoemOcYIHpZTXfqDIu8VP9JhkzxFLHfIz4ywbgCcQLtVVjLQmEWnZ4C2Mpv7ljEyvGgNh9YcZ
ChdGVo/NuPrIOXsjN25C5cAKv7zUezrxipoGt3MGUz+T1M0BDPW9V/edVhC3eopjn9i9qduYRyXF
AIziZk+3jMk54dK9YcJGETA5m+VnQODvM71aDGrImDk2NrBkT7ez1O1Olioaunux/CpXgTM3Bn5b
Vvegvp/uOsgssoTU6awmbfRVb2j7CyaJRwV60O5J04QV/EVnvnnmmzg20EUOYgFrtISFeAkKw94M
GK+UXipfIfsAZW/iNj0JNNdYEH8nv7p4n6/UutZiEAnWA9trjCGTyNbL00tubztTgw17NIAkj4tH
8+JPQSHBQs7WjmxHfWMHC3fzlVYDURmOg0U59Ym/rF1/vijcipPn8N2ufRJpx/GWzQnB5YC4sr2y
XjJtA776cCLs4+6xqjctJz3Q9r/9Qz8g16wTO/+cw+Ymy/lmczUzDlCqUs7Jj4pnB+0AqAjlHIWy
AD3mv21vw2IwBPYbTKHbsm3vRM4bGnfOPY4l0V2IyL081KKsbtojndgcOG2JoaWsFFPdtolMvf7X
MyGr9/oWi9y8TgiQY3umG5rzEqANdsPMbrEBpn5e5O6nDOBP6VavFBor6syfWuBSydcZwFteghtU
ZqW/m3zsLJRCCPsOdhUKcudRyEI1PD2BsBshNuPEWlEOAn5OOhy8P3kfZPMLx2yXKcLlXXFTRUtB
FwMe1hIYSUUo0AZzxcNFg9O+LT62R7DmAXcjQIKl15xoNuwi0glmX7AfirTNA1fcMV+F9A3yXEE4
lrNdQkeEIGlMYlX0bDNQ/OIpo5kRGl1SYNaobLWQwnVcDdh7RnzYsGt4SAFuZNCWLmoZL3wrXszU
+5IJvn6zHm/MjBmqyOtvt8ng0Vs+oDkUahHRhRZ84NXCSY/3albKCEeS97A3Qdk71PQQOXXBdrHh
gJGhV8EDLb1IGy/6AEjH85NYF6ipGHplBXbosU+IOPiRYJX71dPV9o1Q7fZui0xoVQ+IFHqhEX3U
lX9PLFNz4jqWZaWKCOCJNHTXRBS2YseM5pOYaZ16gLpvS8SFfVAy+OjPBPhAKnmMxFqz3KS7k0ES
mttpceU3GzwJf2UM2F5o/S333J3/zUjbiBaB4/S3n1IvGkApu1ScvpbjYmSsWmhMBEzKpnO0fPpP
Ykw31yhuArOidmR1HtOsmPSLM/t6uvqnIn6qcrhnJtnwufjEfdA9VxZJYrSqUN5hj1gjv+GQqKqs
ilmtvJr6axn40U+cObHlfBlS5vQBwSNR4B3DnLLbAhf+KLEOLIwXVbSXaFTeDvDH6CZWKsPor8OO
fn/k/FujzBLQDqo7KViVnfcXWfp6gP/5N5+D9cWZEkB/+BUT5JnQlSFQeip2a1u+sQ8mll5o8nAX
OUlBke6O3+Sdad4sRcaHLabBSta9oYpj5fafL30qIQwLrU4S9QwCU9cuqok3nQaXvVdJjfmr1itH
5/vzo7mY+kX53j8Q9oTBSwr0Di+dEpO+h4Pf3uAOlk7mhb6HAqb7bHmeW8Pv0TH0UozrYUgvPzHv
tNQwmX5s5QsKOs9oSn/sHZBLX/yrf6MxPGv087nOqfVz17y0Bb6buJ5E+kpPBFQFbBatBrWXdlYu
HVg/+nDCmCDsXy2KJeIiW9aYBjF19G0zBF1R0qy6IUYkqGO0uUy3kgkXx1lqNchUq3o239lF3xhL
vKRWSO/O7p6OyGyg5wv7/7nsgnYq9wsr6GhhrZQbrLKsWY8/DKlDa01wTyYULWvyWNoWEICpbHlL
Vb1zlihk62sjLwATcl4mWfjRvMVVl9tiVajtAkfhnryXUcncq2urkMWtZ2ntp33Hx9DQwa5lDsGx
i/OMb+sF2JMJRtDNLD3/W+Guedwv4tpQZ2K5k/mWJ3Q511X1VI3K8rtBARez0I8cjhUxWA8S5zVK
vl22QIP2F+i5kBuwF1h3+0sU2A/gBpkB/OD/7vl9dY6cPsEXUxlXGZFXfNaELJhziHLNIa9K5VeU
slSQCCBlSfEwLPJ1ZyJa/amEZuTlbcHw3pdT7qj6DPioMiG8f2BEsSbu6GuQCFsqWMdTn5w3YMVf
9Rh5Sep0vLZSJi8ilDXwyXi6xA/tHQpd9o0/h38pNyXqHypgJJ0jKHW71qDvjALRq4hfmjD3nwKJ
KR0PxMGTdfQHNsd1yil1guqJeeXjTcewHIE87QYYDLa9+gZQUjmoquYvyX3x6YSqNQs7a77KHSpb
fudWACpsQnPA1L6Jjh1YuADs8zj72GTcIqBU/RwMxK178n01qYlNlm08/cTJw2EarRwHygllQpJD
yh71kxb0jL0XFTm9/YQp+HajwDvLttAt78eVBggKAdB5gpheJetEB16PhiL9CvA/Di9lHwmqHzaq
O3SVCpN2n75flqARUAhAvxbv9PqOH9xb/zwBhoqPj2XRvb+dNzWCKyX6wtZ5X1/e+XbLOshNZ/iQ
A0nLPJtjkv1tHQ1ZhQWNiPjL4uOGHnwqVL4Cc75g/0LDEnqFTJh4W/3mC/BOxHf6FqQAr+irVi6D
Az0nukoFYoT/ZvTMdN5wlG7L9WDH97MoFViBr22Hv5by50vylISwIM/ewCShDV9lwUdxL8QeEsVV
Gd/aXMLc6cbfJ1R1u4j4SmqXvYSi6zfSLo5MlLcRI/4nZoIL5RGc/E/EU+KGrzJpQoCF1GYsqqGP
9VLp1+b3VUlWlr9wmcCgXYwy2fgkLOnkF/ADgs3Yr8u/nxgXGXYHPb8tCQrcRHmqUzaG2KR60+De
h+k8HpYpStnAEx6VItdsa2jtHhLjWYQTsEAL8r5gabZOclLf3SR5O90qwpaeivFXR5PLxj+imZl9
81FoAtvWrMdOcF2FBT7sYdkggmJUmAWMWf/5PrR01U0WCp41lQiL6Gn8J6EMO9a0PK+wXTwS8VnL
pOFji1RcKeIAsTezDb+f+3rXmXJUG5+UipyqqA6sgJVaDSkhpmDKSFAM3uKWfWyT6xpZAJ/7h0HY
M/R3Xa8JWIcXRjVKaiGSvH9L22fkHlHY9n9UfpcGVt8dNn8be8roc+vYRJRvrP6zSw1nuRbkeAXx
izVoiPjfZ2UomPZ6wWmBr9l1iEh8it9Czlta4nTlSbplfhdbIjSrsXzmayxpAoEW2As26RRxXrKt
05/o6HFZuCnpVAvJ/bJpF1z4nWK19nx3zxz53kgfhuCa4ReSAOMpMjrn6FwtSZKSm/sfcg35Tz6o
CQPLv8noLuyI/sHckIRWsKtbBWZaIVARFNxU3ZVRh7Dvp+rXgBZJ9Fk0uU0ihPQVy5TL503QRxBt
PNIyi7mGE/26TGcgF8VaR56NbM8bMbFB4xKPnL5AVwZYmEKHeyubUUYMctHPe9y5pqMHE2DSwovI
QdIO9/+Q+lWo8xFzE1MDL7Fen2jjszyyuFbASYYSPG6cXZKsibp1cewGTW7odjCpCeQpU1l+vHlb
OKMNvhdULCjEi/iYc2LSYogxEfNwVhBGGoZM7JQjsFAGsP5GYN5dj4fLnnFMWFkv78ovO15OIqvm
ugvlXnDeLcEfuhvuookwbwz6ysuVNxeRGS/MLtAfZAtxh3q6Buhp3heoreuqoEsW9SBrdUfI2QFh
DnE+CHcdaM2rlqFIgw66RbUqD5jKPOkEgciERnKD01/38eZMkXqhj8GaQLdMtlg3ncynePuK6edq
d56m8oSlmOyTfHH2SjCXMWDDmCZq3b023gZ/B2JxnjCBV2bexXiUoZx8q9JFC/42vfaIV0SMzLPq
jaU26oQWzj8MIdpM8GALR/BMc6FE4cGMw4FoqsCWgkjcreKBnVod2WzZkrCxLDFcIyoVMJkFtff1
zSrV0boGcHVpc+3rqqwHHBfdFu3H4J6civUFZQzEoWu8tKP0JtXrmeYR8a8+tU+OkzOxqJOtq3ss
mlLejnAr2XUY0VoEjuicIyEBDLOWl96U2UN0/aVI54e++fwvOY/HWSwNeQ4HbZkCFax/BplYY8I6
m88+XgFVNFeXjkgXahsxV0LXbhyV8hHWqpn5wfDra+o5bATyaNyatsOgPH6UXDI8VanToMpb9PDE
3AWmTOyQoKHuU88s5yYtctXCFFkOM9QanFJyQwDwu6g/Oyom2a3ecjDKT3H2ODRFGxOapJU3KRNK
k/EfTV8IKA57t8ZcRJEpeJacYLctS6/hDIlcTnkY80M8mw4p5QPc7IgwzLiA67A+Kc2+clQ6HFBu
XKK0XJ8qBi0ueRfAaJ2jDxeCZLO1kcRdALjUbKDiNcwEYELF9iz/VY2mCWvke67H+TxSoz3/WvOM
iDJ7qVSdjP6aSynLLQGPmRym7AUjgjPTDc9u/CrskRvX9A87e2fomVFkzNStenLjXKYRnkRFXoqv
EaqIr2iU0z3+/d/X5FdDNsSLLIAc/zzXAu6GuswKrjdcFRuvqbvFq2bD4lAfkNvXj4fk0V41Xum/
mxXw1YV1m95bbZRuhOZhNM/uYIARl+41IgvpCmroYT/4A5HWzzQG80/gKJnW2uBlV1FLx+UfYnY2
5s3zCrfjrOwqDIMiH+oj5K8c3EsyAEfZ9FyWexCgGpjHYu95/1uQf/7XLkWZdly8LHKLp1H+8cFu
XIjiffY4i1BSBSIcmIqc1v0uLTRPX+ufn5naEbn74shaJzqPeelcYA5DJDdKQzTGov0/YDW1DAlN
P+mLcQpTbe9SSNL7shhrSo8puTrGegVkGWifp2R8zEr2APBdut97gOQ/rrym9D75ttuy7Zeka1O6
nDAoWJ1hmOb1fNq07Ad1+2C0OoOlhYYYOlaNB7kMW1xmJwjJ/yg0yn+pHUwA1orjrrZ3WfCpTB6n
2nyRZpGXqMSyjmYzQMTJiLohsRL0BH6XrtS6O8XhRbUJScfcWinZrWpHKnK+8+5vDiUzILbbLSX2
HUgf7Wxnb0zC98bzVhdQdSjRU4gKzfPKcHyml37SwfQ2ykXS/uL3hrZOCEk0PLHhV0O2qAochTaM
MwUFa3IkpudfWp65Nerf7JHT9wNL/L+ysBhhVRcLjAl2GFx96ss6kHVtWpJS+ibpVRKjteLWpSI/
qP2qfv+RYFbDwfyaYUUc7hhT/Qi4ohQOCCz7NRtgO6ZyRSUhaZ9UKNltGCOZjwEohQy8Mf5f2msA
1hJDITVPLnILHxwlBjWyuAV5VAdvJy6YkfBGfhmzb1CENucx3aHcckc3m8qol/wzv578DRCkp47T
bE8nALwqP38Lq6FLT06UlqhZXHIYQmYxAK99D4eulkHBEr7Xyltddf/tjRwZ4VvWA/SA45NSo5QP
ZQVbU2FBdu9awbt1aCQPhpoLeV5pBUB87SAxY0UD4d3T1EciS5IOTBAVbqu1uZ8rwlI06LcoMCMM
p73EOsIazConacW5pr78eqUXuAJe/KVyGPA/TJT8V1p9rCaf3vEqn2poLecXp0/LPKpzQniBhhuE
hhHUqX4GxfHVuCoNJAHqMIqCLdYCVv9NDh13SoFKmIe95M1UesRolfY29SfhhhkRTKdTQ2bsnVAN
vmJ6RsE4ADdO/3ae4oLNoyCAN2MZT3uXbZxLSARGCCWCEtVyvBO4WurfBwxJHIJ7FQQXvi4P3vH2
Pi2tuQmAQppIYk9J8e4oRvqWsPAxnZVPhZ8sCDVoKomLXMo5kjAL3QJdhSWO5BLKX0PwDlfpjM07
wiuyjTvsFj2cEMHKWaVBbvuBj/d06oZKF3chq8wY1QBJIIOxEojAbXN9M+7JRn/kSWinjI98FJnu
r51ekGwyZzZDI49U8AA08jSYHFAUpT3JUj1iBg1qI32tphOQYs4URBfw1f7wycul2yz4Z9b6wH/B
vbQB+sM1R8bTNIt7po4gSWHB9y7yGLirppSNHzgVwRw2otWTRr2u5xNVH8bTMT3A87XNxPUEn56E
0M2DQiNDayxsfJLc/twfTpmtee7G/0DSce/knukU3pYZngGOn0Of933XRUO4ZejNy4YDwwqixd/x
EOGE/Ql7SHQp/q68p66mBjn/nB6mCBn+Q250UkilfYOWuhWUhHckq8dQR/Z770ORm3sfBsHAj7Of
pZFNCMmTi+Zsncc/AZJuZ1c5oPYXB97SP2dUeFJgkAreNRI+5lO9VPDg6ieHUctHZnVOqfJki/9t
LEtMLxQnxzluh8TcE0L5CIT9uB0apuIvzpTj+fp8DIgxQtbHGlBgHKnlGiI8/x9MI8PeyAAAYQzR
dMdQr11uofcmnDS0l11PRYjJgpBip0gywdrn7bAaAaXX/i/tcDrx9k1DA8fB1WvYIEvpAOJN+ofN
ASCAnLF1QGvEVugszvMXCBcPoLoJHhZYs6d1vJwElGatxXi0GunukWNTkffZTMki/K0Ad5rZUN4p
Bby/78j6QJ4bOInXN8wlr1M/6w7eV2G6cQHhS93GutlkxskfpAmiw4+vxUjTVAWDX1ZJsHe1KnIw
t3XqdM35dl6QYECKRa0mGH2/uTwkie2JsMz/BEhoSxHclZ6Jlin4MAMexCnlyqLOwfUSIo4P0p3T
ozEmvsQANOQMHm8QhEeP76y+RHfnxXqYSoM44JXd/aXJCn5pc0ZW++ddjNeMA9TsFC6RYVcktho3
kn8Oek7nbrImBnt6l4YupRF+gXQo6B2Vds8mCUfndvTheJBOt09bby0U7uqvt2//weYnKU0HPxiF
eHJG+8fnO0asrbhHuU+bUZsvdSXhd1S0TuYPRgSSOX/wkTzU6LMqB+ZqfYWTUcsjAYghkSlz3+TE
IictIQNE0+aX9l8RgG97OqikEwedBn8IfeFZ0j+kfBD6dczdHtd+RMCo/xz9zRAU/5dfa/zlGT68
yYkBEzXErM9OWryFwYha8wE8tULauKpuC31DTl3roObtjOiqmHuve472h0SouIpP4LeT+BVpMRJ9
Vid49lu3boJof2Prp0PL/JJLmqGuzF9OBFt16ld3/NTzYvM0160C9oy2rBoWC1K2Pwh9J927IhY3
Z/xWvk3SJ+WfTO/GDRL5bWRLLY+xkxj8qhIDHhxPJXrNcqjqVxYbz0TQgXagHbZ0fgjwwOMUa8Nx
abhRuG6y5SvLSvMoiKxvn0HpfVAkmuqRZgI3xKkhyxipJFmGhrxapzsKK9I4rybzI5uxXVcyWsv5
jrpJvki5sB2YtCTnaW+LTpQzKi36dVBsp6f9TxJDcyBBCZ3RkV6RY/qGxiKnEik9vlcqiJ1BQQ+a
G0whdSSdC75qOg3DjFVepYHRU+gi4p50Rxcv8MTkOPs/CJOLBX8TRXkYJ1eQ8qNGSwQL8FbwD6ZH
ZqHlJk695tumiEsPIbrbrDhL+70+foodDH6TdcZFnMyzMiBaGWEHEnI3fyIny7PfBkjzlkpnngif
2F2hwWEzVL9HpXnZD/1VlPYzkNa+Uwv20oH2Lm8QYxvwuCewcmPLIzzi3TPINdrP28bqX8u4IXCo
Mu58DzNY6ZhtgVjrzTZ0AXkYi8tGFZSZZ/EnGEUvcxjNw9DrZtumqaTsur1I6eDlNQeYrdEZLQAz
siHWSbF16BCQ7pFcDdskN/AOKyDgeBi1ElRdgHFQT/k9X6zK80FBnOjiugKn60fhUjSy6eYHdjkR
+wFJZ6vmCRoLCMQpaooiAiJXkgP/udwrhnWP5PiEFL/spWJ56eYIe5VgGobim1up9SCOXOLBhp1q
ov3ZqEnEn/Elkb0w574/oe4OQ9J0aN9umi8bA42SlsvJCq3LwpkwzgXpEEFS69/lWr7q/4sKwPLI
DZJZ8S76iPiiQJZ8FNBpsV71UuQjMgSpYCyuvgHhQjvlDP1PFcP3pKC4yJzQCtS+ajzNUprNPrQa
n6o3VV0ao5KbJpkYg71w3xfwinO4zx/FLQRc4iBKczCzAsvkzIGNYCjjraR9YWzh5IdGpdS0Jfwj
dK65U1LGmC6guohTA9sIkJWoI6uyVDwbLvgc2F755DcUm/EbmwLtvLIZzx4o9nLOeCeHMHhLo2sn
xmL7j+TypY58VwzA8W3pHkoU8Xnp84jhJtncosgHDqULBzB7KLsKBRCL3jVx5EGg4Jb3lT15nfiM
W2T3CA7nt/PNtIYm74B1TsJr+E0d4o8HN72mqkHkZDMFlv/P4iB7M+2Jc8bCUuc5ehmCnTnjcSR9
6w9XUNtb6BKE5RjGmYzOa9yf+8mHzAmXxJ+4i2HNSRrN0kB6unwzrQ0yCY+fJL+eNdN8XDiWnwnI
WrJV6C5v/S4Aslu7Gm2h3oRIxBKw2ddtldaA5lnlUH8GHYvF4+SrVL9AgZONcuR1pEr2tvKdml9D
m6FqAsCc9gxfi8E0zUvyy7W8K7e0sQ+K0jGP1sltj9qmuYPCM+T8tdZ4+IjuUUMls594f5uj0l6h
Ra/9lH+CEfIFtGilBW5mifrbDrYqWVYmQR+aHsJT10gHoDEUeLTfwylvDyPZaarLNuO7oL9+6bT7
GHSSaEsDrjsldDngqLdjgYXCqfabGAtCaZcISHXbmtv9bZtedQ1RWdCHudNBA9VhSoel+ic2C9RH
oAB/bGbMZrkmjnorg8aZaDTLExpL8UMplGt0OClgjQWpnOWu2uLIg40MiLnHEpSj8OzRSjKr2mQW
uo+IVL+9kL7bfwNw91AaQdx5cRWPUyt7vDnKwtCm+FLb00GbEJM1f6mjAmfD2l5jMvA5vEHBWtV+
EXkDdfxyYjq1kP1psqQng5TUGpz9Xd6lzVjN6qcS0H16LfHNlbZYh26XR0R2RMZr5fZXNXTVAnl4
7zclSibnJRGnj7j/THzO9gxoWxjrVsFyipAy4dlv/YIgXObl2RaZninIm/zSstC74EX2R4ZGPiyG
f+tjbYTzIffWW3hEbHxCNLbOMhbJ7oxz5BEHrHtNQK+toFVNUrW6XFzyF7LLsBSpUWLKioTHBbvk
q1OBYAQuLvU34tNHcPup5FE6uKPSkVG9kSqIFUfmfm+QWl/mT5snjjIOtGXxqdnEagW37jh3Osfz
T0gh4W+N5car0BRi2eVR+LkvSXuiINAPD5zcdGE7LMPKnu0JaBqAXKcn0fbJ5uz7g+TJg/IUXQba
AHKW+MREkLswC07kG8jZEZSMJCf62BW6xxonKhR8z3PYZ+sUCqeEFUvp1TABZx/GAaEjd4GOEqbg
SqJjk/Ks1jdzNJq/QFDGVq2mYnL1CtIg1fuoBt2w6Q2TrfMRvEvEFZse0Fj2P6zfcH/hsqCeNZce
hliwAVc1gDm1HhSWWKRNYxeFG8qwjuhxJpZEC1bTp9q9ehMLn1wcMOgxQW+avvCmqjbHcQRMiFdM
xowbWBAQvOtssJdx1ir665BBeHKNJG7PBG+R2AT65C6JCmHPHMEQRghnDolFCCa6jDhTtBkN0eW5
7CTY9hd4zl2rID22yeSOpvSqHvT4oSuJ9EWbYG8YQxumhT6Om7kfC4oeWH6QSOyhbVoscWjbzGO8
oYdJn9HWaOtkrfvaBrJoJoy/ImIPYh1rVFChxiphINfaTp+tTGCdGHtPPapo6qiMwPnZvK7jUSbz
eRVqGSkov5z9GdOwAlH/8bktlEVY+v9c1Sijf/heLLqMHgofEpnpsJONoFT2v6jGy2SWAFbN5NTf
Rdkq8sv3tz9/9ExaMKBqD7PQisM3YdyJ7g+ldyUE5kywBX0exmGVsPwZoO7IR0HrV1ioY/hZdadH
rHeGmGwCzmyJmHw6guN8yoieHRERg4uGV5gPC46JWHbsB17SCJlROWGmupCf133+ZsW9VnDR800H
+vDxmavu3xBpc9/ss9bB+A/cW9zMHVDtciKZzZznS/ur5FKw9hhhnOvl9L/4JrIW9kIcrTbOGw9s
OZUXqe/5gQ+3G465bT6d5cK0cw7x6bwLlgPbYZJNXgI4JtDZOI6M1IrQaXpxdW+mkoeVkeFGaVb9
MGmYGoW7ueR+xGOESx74UQTWCpFAfFI06o94TlICQnw1zTqpAII+dLvMH2mKVS3Ixl+rpfugczyd
hisJG/CNesPR1vDZ0ZkxJO55hjkPcso1vAeTnwmEmXQ6xRBxu+lqVKFWSQGw3AvWWujXi6mA51CJ
JMbzN+JRa/PIrT/H7UEtUpRcXZpXIcxHPbaZmJb0Yan5uqNaBVd9ecAhRv+iZhRcaKrJa4+hpDWS
4q6btTSO622kf0SHFdFd8VFHff9qPvy57a4xa6o1BQNjIxnUrID8T+WK3cGWp3//+dScJ6CIr8l5
imrrzaqITHEOgchdXSgFMmT9XZH+U7IvrkTmp3nVv8nu7cNBytqtHZGBVQYUwCA220+M8WDRaDGb
tlSAE+GeJ/k03gHdAmFgV4OP8uUS65ACRIUkRTW7dDiB/rfsoeyEwPXXSwo+s8gnckJVvuXlne3g
ui1W/FDI+omXWjySJD/OKds78+oditLxZN4YIkbsXgcRpfLYy8scmw7yzbgZhD7kk8ozvtk7S2zE
1GZKuUfkQvscNgFK5kar/+Oj0zW1+2MoDvE+cvY204tyzjIWBm34hODkt/CWWfxhfrxgidtquhrF
OCa2N+PFeOqdzW0qP5hv5O5xQKhNTR/NqH+rvAEhrylfRJcW1HdtZ2sKAcLkXhqIaLrfV/PUzrA/
/FDNhpbYzV863DchB8WbB9/PzB5jdEjuYL1addPFd8ugK/AJTDy+Z5jePtrJpQXh4PKK06EZlBxx
Oi3CORI5b+YXxe8NG+FsmAe/o4zMu1Wl803CVRkRiLS1itOfC6tnBDfmXW/FjvUDgIkjAq+qNTbA
kvvTFFV4x/lAeEmad8e4gmrUou8k8j5nyaNUrBCWl0Ceq56d2wUTQ9reVZWn1AQyLcOjg7RBbeXl
7m7Hz92hhDg1Zueqd6bRHk4uMDtTZfiNnYg/KCfftVLnoi213T98BN5U1kbHUYfdr6lNrIAGs2LS
+TKghuZ0pnqnQjo2WX/g8yVlZYaVJHwTqcLaZSmTp/ngg9dcACBxTIblpZ3jByG4NEs5z51qkwie
temsQE7zswJnSwp4lQxOlZf19WqRgUrQia46u6NxPbZ/YDyiIeC215h01DVmBhPwZQrz42fmYYuo
elIpOfRQ9apYrSJxhIfvNkRYG0Ba4KXRBoA+RCJackczo79/PIiffUIrR+tR9OST+lPXHV/7/lx9
Cfz6vhGAxnOCJvGpd9lVVZyCN1xtoDhut6PRO+djLDEjmZ3O6aAANoaQYh0C2/+PzQn2R/5r/ANz
A8FRwuIOntDF5F4SFdKL4SMmC1NrfAY2lhNDVD+Rr4PZQPou+4ashgvSzQqR4PO4ZqZjIpJrMSXf
ZxcARlMLU+JtzgJsrIBtc79xpDcsQx2FHxPkhf0ZK62FDo5MM/lFAgGtIt4pL0VaRSdbAOtytnRK
X42HQmMrNkKFPcpQM/vUw4AbhpnQ1jHO3vMUJmTVYXZ9Yx7iwJn4qnBA/TCdAEzzhurE7AXOC0Vq
PSmVtmPKYOGxkMDGPwCt3BZaRVmb8Epd9zLyGV5lfBFEVCSXnt25aA4mUyWAcE6DwkzVGGclF4YH
muyKp9ShLRzd5YhonMfYipxrr9RX8pGD69PJZ0YexYubphRdsmIpr+Ng0ZL5/kCmqYQJq95PUtep
WzTxTuXPOjgjnSdWv2m6zSBLz42eRomIxyskmjpQ8nYwzFw1AI8EF0zNKXnnaCL+cpkyZUaaFwUI
sAR+KIOKOQmX7vs8qU5ZFHKp5iAkU1WuASlf2BoiDVKWCflOOlmobyVS+zbiTN+32oui46d8CNhj
GzjtbKMZoaopN5HuhAZlgB17dxY+qoFuRMcGFeKd7I1cKRZDRUHS2tAv8Uz5rtwS2jiYQVXxYzEr
HGvgLcPK9g18yDdxi4LJE0mcG5Rvw0O6IPnYOOXP9UG5JPlfm8G1Vhyn2JmW8XcHMhxzgPyIDPQO
no7S5p7ZFCw3wNM1zTMB6mI+GHjngdYTGIAwRynzfwkXMsQBvtIoYrj1Nfy2Xnm4wPksXo8JekOn
65Tq05iidk7Knzj//ePFuVCnH249j63aasnG1pXTW3Y1yghyMOGhVyATYjyH2+5ZziyzmMzz2k0x
9wg+YBFLP6xfIEqaDmYmAQAVQVFTzTvfdAZzq3cr6UGDhWvVueIZu94sH8p+UBxxGAQQcqjtP+PJ
aXVNsx9JLGMTVNDGYgHzQbWCzuZk+YAtqxl1zn6QeUGjza9Z2bLxxhvMaHtd9w15+GN+3+gO19Go
1k/EapxYbweHPJ6AtL4yMqv4vLXRckedrcQOQBKDc8kXzrXDs6o1cq+9vqzxqq7hhMLlKe4xds7o
2zsbhw1rVx/YG6wnYzXYt42Hsg53YBOz2YVUmspVirLMMFTYS369lUXSsOI/x6PjdfWIxEPt47ot
nPSFcot/cBBRI0P1LjS+Ih0IqiPftx7fxuH31WWxkY1aZemDt9W5JCFu+Kkcuh04OQfoDZHJlVbA
4sScNgM8lJfdvNiWKeKvOFJMP9R6eERhHoKJl+Bc8XHyJ8urGC2IzxRznqFHGXMXEn/h8RNmfdD3
AdphzjhGweCnLI/lJtpOheRGbzTvKXLFIFdSkaQZpYJL4jA6NPhgrP516wUa2RykbhP1+oycc8Th
Ey0ubwS4NgxteEs8Cr9KllmV+3NXmUJnvFZIj568izNDkgVfFo/iRYDHtvkLUrgrjLS6FaPLwfmI
K2F75uBYwoZUiGwzmU6ojghb8Pu0Jue/By2rep+I4e0mT3PShEud2Ff+qfECczsnZ/zLWp5B0dV0
ULURqQRheqHKRsIN3XcNegozYV9CcqdIIbvTMeQPMb5rBg0Pq+n6LgveqUepqwGTqWo96pKwWGc8
VQs1Dv8FPc+/fBBWMgbdO43tPmPxmdKH4SeMDBiDO5HMU7ksvCfMB+Wa2Opm/Bdbq2+fBAhk9IX8
aGKnir0uRk24dXHG+7AlR6Pj2eYXG+Dsps/Az7B9m3hpNWuih+Ozwr7XLebNFpF3drLeqspH0T3N
iNA3N2L4+9UGUhfaBmZZEHd1dhz/+5WUivT8u0fcZg7sO4z9LWd3FbB7/opKoTVhqhthModnSmUL
ecXeeQI21ll2515ThsWZOSkk9/iDr1X+e0fFYf2RJ7r3jAB/ftnPHltQA1uDFNcGRdqNskJSCSz7
5wbVgE+YSdTuvLy22pyvazp4vtmaMxOC7KEL5IxtxIoIL9EKWyh01hTnCoKaeBQaPKejUDAQ94mO
dmHl2l0QyFaOc2/RPtN18L8HJKbV40WO7otgDDdtePGAo8FIpJFoygf6mFX7YxELeBjS4jRYWuj+
wHaa5kmvr3rMflPWqv1nc3XjYOgBzpgGG/bpfNzujDwkOVhCQsyuw0fv9MhUlCw5yQnzonTIgFC+
kFWfVxqR2r0CZYXxp+xXiyqQ5UINemkL6zGQMWbQtCS6g2J0YGa0Bl4vvUbkWzM68m5Wc4B2HDL8
kQi56md7TbflcyUQBRj4gJkB+176qI6TkEHhhkn34svgQezQxP/UoxlElij3ZXyfUslOL1oHfu6M
pHC2v8dPHMBTn1+Ku4wAzYnuwJ9JsU4ZuXAmfE67znmfN0NsMFJpmTSBnIJNqY2h76ywXz97URYh
BHZlxZqANnZ5bYjXD1x0t6Tp3LKJHtSDa5vA2p6N8gKjZpy9E6p3xqpvcJZSu/DcQApIu74DlXam
KByfn9gCf6LhTtjAQ7/TmIDZXIDZytBXINAE4YwsJzDpYmcdB226tjHW90EKdP2fPtMDfdh6djNo
YvbOm7M86d/vWmpa2pqVNV7PZ1K/XQcm05nYmaG83kwK93t3YJa/RU8KN4ZmIDsxCKu6c4AbktGW
MaSZjsMcpjewRUZkoI6DZ1VjeNNdA7p3bDpxWl9HZsujDx+PSsoJFUehcaRTQzJ/JTE8/I2GxXAL
8x1+uy37ZzP+Ce2oSgl11H+JHbk8KTTlhrNrm1tj/7ETv8RQR8ca5OT8iXSiW1N5GMeIltIeLxLV
UaDWLj/1ZMbPAS/m3jdZg7UQmuEUh3ieOLWLR+qo2Vv5+CrHJnrQa7+c+/oWqDC+XRyToXJwEYIB
Z+oz1g+ZliY6dRD3V5vigQXZeBTaVU2e1uB8sQMGcPCAKVDRGYvQ4934WEcKf4+Bk/2VaInJNG5Y
bJA9hNMMFXCRvKdCOor8uK1ghpmEdg1z/pTDcXI0K5k7FAcrPyS9R2hrxQsi34g7Y+tbNLk/f569
pAgecZlyODr63iR3lmgQot+4iX8WSUjg8ZSyBAZGJ/5X8JhO/8yiOKicPNAvLDumqo1Ax2ZmWTrC
GcNj0B/tv0ncpUhBZqgrB7uIBQHkHcppzaCLA6cv7VanMvh6aG/bIBAfWP/ekngOJCWiDnjfdjpv
RBdnPBCjDTMR3qRdz24Id2ba7SetT7pZ5VsB2c5fVMxtBEdDElcV4faJ3xn4MBEm+SKMkF8LVMnY
2F61VwMho9gBF2Ewfr758P4L7GYWN/8bnLreYwtLyyxH0L6NDv8lPXgY+X1K6L9cb0SOCIy5etiC
H3irRQOV7VgKJe80Hb5xX8DIGUq0ltXgNF0emYWnENhwUYWfXvZWhe2FaI9rG/3lxR664JYu+2Mf
D+GAy3jVWS9dKcqxyxBoNegRcZ1tgp9K4Pje4UqS6ZRyZcWbwy7futphKkaSUIc6vHKNW/OU6bbe
4EUloyhsko4SMwl5pzsJ5b0nv1ChGUFRgTS+JG+6A+zyX0BL7yLYuSSpIhJI+QRyCr9BRxmEHqAp
oKGcY4t1gees4blI7OHtuay1BT9Z55lQXtFzvxT/lY5MrY/IDA7FoyJLlRSdZYB8u8YqLS35UVfo
AAVdVyidS1fnbPrTcvn5KHI9sIa2iShOXGiIx+98JbwqBOzl6rlTzT/UsqptXPfmofUDOBl8LcmB
mbEtbyv7JmVQgpUrhChPLCDp5NPMsnmu5X5oMW7086rnVZH7xW50dSdZfXQwGpckNsAAiVKwNcF8
myCIMnGwVydMCO+Ejo/crsJt760T0WNMGvnYyVFhrlZ8jRZzJKrKoMnxJbOAYoZsR8Pyxiktuvu3
XNlvxYfliJ5hAW4rnn0+rydUbUeYT3890g6dYdoDlHDsWH2K0TWTAQ272YNOBBeN3/k9Oy2Yn5Jx
f0R/GTcIFH3lba5BwGkE69hmQiuJaVk2C2abbAj8RyDjjDiFHOrOn6/sewxLM/Ghd+gcI1BYbLhS
efyh3RPWaB74jeI9szTw/DB4R99C7cWDcM/aW81vzuKYl0mkv6nvD5V1RsY815tvxxsspw5iAxDX
W98E8M/0TZCPrYrjU1A4o1Vf0xKf96K9d0ixI4SBuEXG7U1Lni4rGMp95USZ2Z0dZY4349xZVjGZ
JQphRQAVaw2lH8M0RfjcARmtlsOyPq1bZeujNzuQPCmHVQ0wJXQ3Tmbs7WJUVr7VB8HQ+5z5sNWD
C+q9qOgaSeQCeYMsFad9cLjz+uj3gHWSE1bXVpCI2St9X1ZtPC+EDUVCGmBBydtIniwBYWSaNKXI
c6eXpzDoWSociuV/jm4g0iT1IopgAXN8uOd3KjT8tqpkQk4EAHIz0I+8gSj3lzLpEsOvKQHlOEYY
a0sVjKTWRddzw6RhClrtfX/UQC6O6uPz9DgvWoQFFeIr88PksAwv0NrWhsj+AU1bccQEWx+A0doX
Qx0pmCHuzcg67MAhbWueAF0HoImC8gBma29Y/ZkFqP6wglZjN2OdROL71qoKoTOXLpFv8jMyWHOg
jvEurDuHKPToduEF88Xv9+81M/j5Uy5LsIMChr9Ctx+L8WGu1TF23FJZW1Z7+Y5S0R/ZdiUEp7Gp
KXX4C6VxjvFiEDQjwfetV604Ly+/E+E8JfG+PjYTmpigty+cCxnWuZOYldpTstuLoJxac5UlOLzU
S0giVjxckabQZFtIWrmPY17cbtuZJJKbMJEAc5eGWOV4VXAFjdTLG1yJ1lVJUeDSzwork9pN4YcS
Go3Jxi6t8HfxbXFFf3aoLfud4ZhwOMERFs8oHPSpa6gjaT6XNYFqpBoOBYVQ0hjVqQCvnZKri/ox
DLxzUsJHCk8wZv090h5VzOqQLBg5neG03SwniP63amfqLDs8q6At6Ooa859pLInZs80TD1TEOgyA
e8OqkjuwIo3EPjDNugTNjHcLH/FMBdNyrEKxgmuQ9Vu4NrX32/+UYBD1oxwauqgohAqPLeOjLZHB
4GvOztGKjJ5DPvhoFeIYyaDPZ0o8Rd9TQy/rWb12nD63MEZ5x4AP5K392wMgkt3eBU60Wwak5kiq
091p2Fqxjsh8aORRrvLM+vw6wkPDJUFxc3ucqsxI4PT/LVjtqhVl4QHGdFAzZn14nR/pKuimbDUg
/zE4sXYHDzQapnVdEJBFYhmRnqJPv1Vi8u8iSWJOYO9hsH3/CHEh+fDQ0nSdSGFFMIYhGqZ5V4ps
8BB+EETNeDsmiPvbH2U0u71T003xzSYV0PAP0dewjDxLxxn3uBUUaicqVj/oMEPdFyNQ7R82VGat
RMSF/dyaHkf0KC1f+ZuNQZ+rNaQpWFLFvfjxpcNCWN0iss5INwsqizkSCuuRQ0dnH6FQuRiKKeOP
cdZyA/lzi8POAdFkRDKgVhfvTTPyKSgQXwVpO/2vN5HDYAPpQDJqE/uGEwxZbH07O30PVTZu0+El
qj/vQiovHQNR2ldRAPdU7SuTejODXkZofuuiiCPX0OxoaN/0SK9fgIaH7V1hnoilC/3ObyWZuIEp
ZbeoAhaYYtxrnfLPpdzrE4UpXEir80PKipp3D0GC2aOsnSaJURQgyN+tqvg7hT3vnZJio307ygBb
9O4k0Ct7Ai63wzyQXvFxaZL06LU9wrQboh628HscPrqGariS54Haza5EpzjNem6xPp7OayTP7sxu
B8O4vOgYV75hcmEcH7vjjuRCUfmTwrOr3KshFUmbdgJwo4CUt/j2Eqr9fhM6N3X9aUiBu6MGUsCd
FDJoKK1VVsRB/tUiwh90O0X0urzRMtm8Odjf9eM54nl6knx2UFEmbHPBfcAWSDG2tbMGLxZcd4K4
e9ECWtGO05SlCSMtwSWqhVjjA3mJIBBxo60A0ca4yy7CbCaxsy4AJykThChZAFJ3yqa0OuwGnGEL
zlMNWhP0XrF4iqLyqUHpcBm2xU8sMaLB3HjYap38nKgTglWHZQmDeEwAIea2UPLoSzNSUQGGncR5
mEZLsggX7r/ZCuJrf08wOxKdF8n/z3PtG4Zc2ODpT5ZyfASyYAP3uMgT8QXfOHK7RnDCb+DRvIjO
m2ytU0lTn//z/SSXLqB4wr/1Kz2AaruYaNgCWbRMWh8heG4q+UOp+5niTRhPOfKPd4zj0kJzGzWc
uvQn9Y86mzvwv0Gz0+7o3iFLEU/OfutOGAetrpoXOnQhF47XIqRcaz3qTD4n8FA/PZa8Ent3JyZ0
IUW9f1K8OAjKiyZyfnpaxwAg98usoFh0qMVAIo0ngto7rX0DQTDGDocvA/7cWf9+5yLBWrXdCVnL
9akPvFCGY34hOheydT7pwRG6ziU56kaNvzvOeG4f4HutIWuNqOjOOnpIPt/ZOrDn9DE8b0/jA3ni
E4MpKVfHSf/MGPwJMKmkKXkbSMNDwVMJh8ozvID0IXZq9oT7sRhnrwhUi+fszyG/Q1kS4kAuo2jg
e1lg+i7nf35z0Dj3dDyM3rywPt5sIEl5bTFTipqCACHt2nlZx3fQjH+qftku6u1l/3rzX23QBia1
g7R0pbJGjizlaghrNskLYpW4Ke265TiUWmGfPT+dB6/WNzQfyle+Xp0brUu++5mWtZE6H++6JOpa
r2tBMhGNOZJw8ooggw0oqZKGKeYRlG4JsUkX/6K4Mnp1JQvyOUu38G3m/9+FcN+mHDc+J2kqiVa1
MXfq/nQhwR8o0bqHZim5tDaTIOWB0AFLu4xGSxFrAPw4Y0ToPIVVZjaEOLlUH45/wGrEMFIIX/AP
359Qh/UcVjePT23q1hgnzQVpfEM2EsjI9wIi0iNlucLjx01OmCtbNbLMzhyOtV2Chp1XytKz0tEg
NbtBSt1DWN8iD+uFn09eqBBzVHOk7R62NPW8SyOYrtd9UrQKNXlRwawyi4bWkAQ6dsSBz9CgNxmA
2Rj4zoeyMOJ6GVlFe5ad0eStSL58V/mTbZOcOFmSGJMoVjJRKTpDNyRFeydnnOSYhJ/OSKmregtC
rDmns78qjZv72k6vN7zph0YZx0+ZMCcTS7CbTrbqfw9edMG+ccEaIKmMPFHuSzlw3oM8WNTJJwBY
mt6y3MGUUFEqnlt0R5i/pzLcF+MTDsKuMNgPM4Yy34vd/QWdjoorFrn7Pc3h1gOMDHLc459iu9Zz
1+VaUy2JDoKscCf+7hFuCBKqvAVCdj2gvAESqEwC4g3/904p2xmfME1OduOZPtJtHCIbcgK22ztB
3O8WGqlVxg6K2wI7OyRACLVOLzqmrj40gv4/vh0cybqiCTmjRqMjd9P1d7AsFQkRXhTnEGsU/Qe8
Wme4SrOSHY4dD2rmOH98XYd+iJ8i9BE7T5CmeWzIhlH5noSxFMqj0Zss3kdCyk2T8NMBQK6uwVpw
QWTwnZ62YFiXfY9qsiRgBKVvkvMsZ0m/dPZp3zH5TaadjcoYDMtMo6CRQjUA3oQikHd3QvOlaHDv
WJ4SMm517FtGodAIcUS4sCfKaWy2rWG/i0vmYYlRvAz3ISNq0bI/HpoIzJIs8OKDIRjtXCfL1EDV
GHAVYjlNGM6+7jU3dQpicrYsNfFCbPynHmDcUvWUBC4Cpmm8rl92mDLxvxbyAuYzKwQ/FXmKi470
Csp799HW9z1/EAtr8nxOPaNYvLcdsZ1RCrYYK/GsYP4khMFizoL2OIthqovjmlP5XxVfDuU02y+3
bbwQI3MvP4xBwBc0wFz0U1vKepVrDVnTP2ec5MdkVsFSQ52oa+qJgzhOt0Bu3BiF3LLoBUKyYdax
j8kW9XzoJpVGJUFz3GDLmaHLcP8EYXKJxt0VoDWaySJo4sRSlrCHbNhOPmp7bW1339m72PiKV9CJ
NAkp5vmkCvE644aXLlPTFR3MzODZTNbzMf/XuCtxthfYNhd1twAgFh07YELKPCtUCot/QkRBg7uO
W7xqf2oxi39Pg7b1aKt/qtggOTxIt0cmyIyvYRFoYhHNoynOnQ4VEtOle7xPQ6HbUKUpkWQFp2p1
rHchTQnJIK//AXAUirz36QPR7hYq6EUVzxVCxhrbP/zcDaqtz9sGa9fE4qB6gyBM6EF9fPuAeQDO
x9tcmbWa+b83YpCNP/b7+pgUvsEeRxAIqVuOdcbqNiIE1l+kjFUfqy08MchzH7wXO4eRbAUxaNxo
B9Fmaa6oPl+x+kAtanUAvfaVv0kDFmQuP0w3+FJQOMMz617xnLu+rigiOgSNzASD/BNCMSDfvaQh
yPhaIX+lda/dOwX4qM+INsPc1N5i9IIF6VsHHHDJxoDCnq4GsBOpAdosCQI1obQFo4nAGmu9cM8N
Hl1lvDZydWDdMH1E8zH5a9XEMffKLgilBqYSfyhRoTgZyhZII/i5Vi+ZU4MC8Bsz8nRc9r/8C5+4
5Yf58NtpWtn/SBSkBQATRLpjJlehLTQORm2IwR44Rl8OnHnoL6zk6Bm5ohm53MSrkEIKLpWCxoLb
Wzz/fJ5LO65fuoY9OH3XhhhE0CJnoyLHLITRiQaARqbigH3olkQ5B2sQx98wHqDkrcJovyKglDRC
DSF4GfIcnDrtG9DOu6hCNt4VjKe1vfwzGfLmvuLaYtMCak++rdBq44kir30Tz+n15BAVFcJ6DuUi
qNXXl4pn8AaHDQqt0tKL3/RpOKvXbBajptejmiWjW0bQDILET4rmCR8OcgGH1u416rOLGWnLLeAo
PtlOfb4s1S+Ph0rThx+SXEzKCiMbZ88/4lwqEfQMYSUvUKqPxiTtBtukzXmWgEHzBRDovSVYUYwH
/rV27zn9+g3AjJAWZkiOXPqMsVgOb5QXVFEKAkZiWPcMSkbgd6ITSJH6zhJ9+btAw2OLKRrBWSCn
fEwddERCGuip6PCSMlSnODlK6Z83iuuK8GbVWHrr3QImJbrI/mey+gPGK5YjUy0MJRQDbMIUyBC9
sS6PjJiw1HF9khDs9izBk85pB43C4HJ0ZAx4b7kJ6QW+ivZe+JePgaVtPXkbFNNj0w4rGjaB5Uz1
2X/D6zSfAJBz6TDUDSpK9Apo5ACjmbGB0pEG6xoRA5blNXyze5NQNSsfsoVlTNswpif1SXHhBxxp
z0OWzyFivVwVBk0FF8LqVOW7Fmn+o7KZCRO8HozW6cljQf7dsR0DEZax3m5ulJITH42yzUqP9WYB
rinF/yIzeaKk0ICxGIStNttCFC2xpfOfRH8OqK1g32NSC96+sc7sikyc1EjkMAvsTD8sVbJW0iZS
PvePaAT9W9C8ze35b8bt52ghdNsILYCtVvu491QXQa2p0CyTXI5+wVfOQWWZl647Qi/trNln5FGa
Ca5tzxs7E3R1jWz8zVcyL84wZnxKavHhKPqEHxHfK9S0UYDoMFurCYyQdLf95/38yPj7ehCpnT2v
OzqhTBWvy1jMo94rpPcLz6RMOK2GR5eJt0B5hj1xGTPAIuDLWC7l3KgkcF5K8xdV8hwKig1PVvtZ
MXsgYlrvUKG5OSCB3xGDzQeNV6kiBGSoTUOvGEtORey0C2njYy9iXwX7ESqNpzi8u1MT6oRpNKja
3caRUEwXeoPYIJM2YSSY3AzZ3r/rbrEKeA38A1UXR0qLGK1Zln3MnIDTsuQpK7JK5JnRoaXq+iqx
PSsLBAAoIm+2m2W5CcKiW9yh/3f5MIut4XMOSqFe2+EGJippPAtfPB+UYLAwPIOmy6mJj7IfLHnW
73WSRy7PvnKOdnDfo1R7UysqdVu3AKG2aP3vj0x8JIUJgj/7Do6bRu2Aqc/uyzUk5bfbdRqgRb3c
ukX59j5EGN/3x3asKqlcN9A/lO0LMOOHWQlpbTicBH0iB1q3kwrsKvx5YdzfpSbUa5tHJwmgHa3c
vja3zr/EY63JHop5lMsNPIbX3mDbcizPJK5VZanSGC87Gi3/2dw7jvbyn++LN7dm/ffd9GCyPnSV
en+VOJLSiCiUOB2qNzSc/1e3SjQ0SIfoSKzWiIUpEOStmsImbp61ILYMywCn4ltFZzG6iNSvd58n
NIiwNRkRAgTNFxNfemSqSiFpkQLXJCeRxKTzZFN/WzfUwN77gzdA7drE66loXnhj9jEaRwDVr9+O
Q7PNbHdjPsqChIllSO+9TV7mTGZGEg81NxNgYgZXyTnosY7+4ZDt13Kv7S/HPQ2BZjSUcQq6rrz1
i5Pkf5tK5dDB562frAvGxwBqXwu1jB50BhIJl8lKQY2ZD7NdyaJXR9CdhsWVQT8aC3bL3tgx3geA
Z5jNrjkWNoxcfWk8yAId/Y5jzlUuWwY8Z2czO6i3E4CGGE7ABFWZQ7g1fwM7BNVZmLhMX5wE5Fu2
MWgtUiJPSbICTrpsMw1M0ZhOsjLwLK9hW77bYWJgeGCJisuFeYO+0vBTbSE1TC/S5jOOZDoyNjvA
HKDEPA9gdrPCt1AfTQufZeU0m8VzEdEzzTde0FxVhZJt/7tmJVJI/RFOF4TWDQ4SUBI0jSpreWaO
V7uKPNrVQ4E5QEQl9AeKLrLcdvokZBNdthHdE4yJbazczbYoJmih561QunY+VVEisyf81L7R95U6
9wssQD6mZUVXtxcgNShS8/W39Cek/o2psr/5iOiPtuuYEnUHB3sPf5k9oHDRDawidJ35WssnOYAs
ZLN9D2MJ+P9E1BaKs9bxFsIL0D7UCtcT28C6E5Ql5sGhNhcD6oeJpvDeTLhI7dqkLC9Gps38PNSS
wwbi0Ubw8ul/jWXDhBQrIeIKIGjr6M29EHS+TLZCNJH7S7Nfp+eRvSpA1l/0CPoejP8bDiClexbu
eVcTnikBCheaJI5HBnxOQ8YpT8oV6kRqeiUuMkqcCQmZF73oXpdtsCq9dp/kCQZ7aX8fMLOldLol
56VryK8vhA4v7MOXIlRJlWSlsL0S80idVGmhqY6rWXU/yVAnRlqfeYYK/Uc7HvDYWYNxIXSXBXcq
1ZgEdUXiCBy/RiSgtf3XQl9fG8+Jws+zZT/ffFJPGkQcESTlEzj2iWgucBraz3gdtWH6+VRqy+1M
swWf8iA74JhvJQjpVoXA2k5CKk3WB85SXv6RgkNbz4uv0d2zL6rTYRc/3HmvGMm0MVGirExZK2u8
7ln94eCh5pB4VarVG/bVLWXfYOY3agEfWYdsEbd6SSc1Mf+gUVOhaZJp0GXUWbueIh6RZTU0ewuA
ouaE9Fn52C/BTsZYt5S7wmfylyphF6BXd2PQ85IiJ1WE01rZSUo56dOt/F/G3RWYXl6vGqyZrMT9
jMK54hQOCFgFW1SZYc30+99EPYKQKRWRKIDIeO90DgYbp4wQGRhYRIp1955GF0ccVEbaiJ9orz8t
AP8GbSFYlbtOdhSgOGq2jtN4JAj+Xe1q/TE+ZRy2dZgUCGoiz/Ya1CltWy3xOiLscXuaYWOpb7n1
rGcURrqcsqhTUg8a1lvi8GV6xU8B7KByUVmELup+Y8WaUz34uNMS2orLC4tLWiezBb7GGsH6s96b
V6egmzsN9/kSvp0P9RUOoQkZWTkXQxoXSaI5pcMgTvTzRZ/Y8mKHIFTPyX+mPdYWGtnVvXIzpSxo
GWsOhvWo8dkKYJ/RrfYhwPudclyimVIC/B9jWxLOolqqeRrhxueiVE6eqU8T6kBnfWvPXmsVVZRZ
zcVLwCYb4tjfEF6nJQvvchd1l1P+hDB8c4VRIyJ+nuWMGM2/LoWFj856b6Yf8eT/mCBRXcpXeTCG
x+2sAp5fQdgZ784kLTiQgdVI+5YVJYYpWddKuv8gFRUnOIXGeB/fIVVu1EBhdqYldN9x5uIG3DLz
6kha4OypuMrT+rh0gmYCITgaIUmR+He4n0lwruUOoqgQi9Fu/mcmtCsaGplxvmo0ExI4vPZVY8bN
hmxhF44ueTeLES8v3w/OcZe4wrX9ugfttOuOib5dCRYROggsAPVllBZSuw6OiZPG7HC2RwoN479j
vklEq0ijZAgpO536INIAgsJhK3/r98f7ZTCXSclBio0kOCJSIoswHOKI6KHRb6wGS5Q5FuXpeHqy
lIRBdnIV+sPVsdsL7fgB9hG1/iLhaB/Stj8F4wVvpR5OM2psJNtLCrKXMMGmJkd5aSHdaJK0RXz2
tp52ZeKboUI4PTrDQvtUFKRHznS8tS/13XLcYR3DGUGOE3jPC3g72JlaZiQCh2+JRGG8N2MYq14x
67z5sNLnj5jE9V9kp/bh425GirOn4w108b35TRPyvtgjlJ4OJ8/atYADkv9hF4KvRN7a7OkSbuH9
Jy0ysdu8sgRidkuAWLROgOhwK8esZam9JvkgWTZiR3UWYn+vXHHvYOFC+CGrsYJ/6X8katEF7rqe
2T3lm5d8Ad3BK9ikVXtcLJfv3uBFRV1WWwarj8zwHZulIeGdo31i2WlAcs+/VbAYs0zziLZbGx2F
TuGYYoY7zKE6f/pzWPo5vX5+me5m7A63EPVeeJJTKirgGI1d4CUp+u7AkZXSS1Tw7vQyQqc3jSiX
n9b9BRIQZv8jEn1OhZl3tqzLTUG1t6KaYYaYpcfEE3K6n5IeWvDyQugsr+0cBg2MW4TB0hnvcdg7
Td2D7XZt2VckQuuiz5nnWEWTbL+ghZlDs5yplEJxOF53TnVZN0pc/Kian3ET9OsUqkL4SvltoAAE
vL4uZkVi4ps0bCL7FLXa3gyukY4mVT/KqxVc1bm5xEyI85vkbnN3UEPF0PidooxJ4+css8jw5h26
xq0vaKLhXuQFV//sVCTw4IVlLDiN8Pp2k+knftvX8V4wgqXd4fSYkqKHZDNNLVyueIgOI7SQOFd+
SJfRCwUcayK34UmHw6QgOVO7jt0smvLhTby6FGOBlos5YsLoNQVmW47DWjsB/QLsAxTOoJtK6qaG
UJwLZw01RMUg3m3WpjvZ6cD1IdlTBilL+CYs5NIL8LwAr3mTqcPVzQKo/5AbqDpsRxshVFBnKfJr
+P11YtmjqOxQrlN9eVdhrhzcuGgawMt0Fx//2bTdJuN8Fd/wgGEE8gH+TM8NF0mdrw5m4HAGsX/e
JWMtqFum+X4Pk5XE0LZ3Zcprf6GGOwyKxI2AdqdMhkFYnG4zZXIEFVHHRVB5FYwrUWVH5tA/9ePl
916OkCww+Y2eTPM0rSX9j7yacfLZewha19GFpYo9/9dqHjWzvsMR0I/CWn+fvZX6OJ+XRhyy3ho3
THP54TtB2ldWhZeKMcNZm5O8Ofu4+VxcyO2fR1fNcREZU3xuEuUn4K/QQzemWCtE2lm/+HUgA7pK
QSyaYEbyGli6pp4f8AymYvuT4xpNVWsr/A1fLC14OUxC3Ny2CXSh4im4WKO0ZBmcZLVFvC94NUa3
zl5ALsN6T2x8l1idM70cs2DC9H+lbf+gcpfUskEa4Os3LC6rgXDweNQrx8S42IZQzs6cjKPKoruF
j/QOk8rQubI3JROGJixVNU9MNMzVM8C47CfENpYGbzldp/g8IOGuT6t6HA2rvxeeAoC1PbfNW34z
eWsWgvHm903VMYqmIbDvQ/mRRBGZwgJAmfl2AWeuxtBb4o8ddiUAu+ckxgd7LJ7+V9K5OWGH1YZj
17EaaeDWVth8O6uzabGJzEa8MzgopHiQCEKQvHYiMzYp2aO3M0tqllmy19Q+Up1TTmXzz4NyUWdQ
d7DKmjT7ahaiKAXs2GxjHFtk5g1LuKahlltCTNDphLn/xfdzQQ2HXuun6eHTtbUakG744yl6L6A6
45Yc3ETf5zyOEKnTaVOVPVFFyGLFKm/HubGmQWt6aMdYskjdvReLb83ok3jU8/wojXiLSLU2rG4y
4ULu4enD/uUtDKcXQz/d9N/lESlXNZAi9mJrZJ/qCPdRgjpkxlYVyzzqw7h99b+7Ej8pJfEqdy/C
JOW/I6u+qR0pUNjpT6iNQMiYUvwEkWVuu/K18e4wg74JPyfHCvtHYAIu5iexK51wHZaHwSv0dFXk
xBzF184mDGauA1F6ZtSPrDZKZISFEUax0SONMqKxld+5AqimIEvO8gU0BDWrOSvEYwTH/+wcHsn9
uGSmeLj4jnUpB+Qz6C32FIs3sbIAUb8XFSJeKe/SMQDdUqfLA24V3VgtC5Ndn/HcypnLx8T/budp
qT/evcSkQiXgyt+uz7nFO4s+hRhUsNA0uJROnS9N/NO45XZOIDwN83XwQuh48cfyBb+EWbN0Gsa+
NO4nIvViJTuRI4BQiM/UXVqUhEbnwzUyy6MFB407OrffDbbSddaVTdEg0s5JjP1eFWHgfeVqiuPE
ic0eYivNR/HeWkKcIodJ1AJJlFhhywDdQPJT4YOJ9RzeBbV4a5V6aVDESvO2Pvc3ycSLDxQxk+VY
Onrpo/CugGz9t7TkgqhyXwJHEz69VGUgdQwKvDbzmpzZJI3ouTb+TPeXDCtpOyYcLWWytye1vbH0
pyIpNcyyYvcPTOEtO2jr55oBwkpiGtXbE3CFN7L1Q9mNkRi9ZAeWerUGPWGAC3qoigC06WJuBdVe
CbkvO5rUObrIk4g1LRGXddBfn5izYKARtSINquPJjM1Wio3N3oNHPiuu1KnzHw+tkICE9lGbhrhL
4YBP869clTPo6tLgz2Kji4kzdVLTyxdps7d9JuSTPz++0PNj5WqHq2+jqRmA6Eg1sioJjXQObL8i
dPJx69JVH0R4gyr7gsIzqhilHR9CSEBn2vTYOReal6/SkzBhUoDLX79/GU9oYWCIfxhDvH6qiyap
VujSzgj+RCCLPE4YgADQbdsqsKXuzpXcZOVB/53tH31EAHSAd2W0HSV7err841T+kHMq+GAAlnw1
xrRKW8NItVMQGu+OFJjMiTPLwik0ZDn9IhDXb5Wxyr2Jt6uQWqMeFM/rnrFAu0I/Vt5D32Ad410S
px9kruqEAKfkKA+xg6UrzuT2x1EH3ygh0cSkEB/JJ65EJTNPo67tuVT7TG+lOHnIxXidM2dhZtAY
AmG7DYdI+4nOrF331MAeK8RJu3H1bfx1Or27lHjF7SImIrY/iqzNZyni77IpzmKes/OXjGdhq4zE
cLmvnzgcNHGdyQatdahJ8drGd5JwDnXxg1+f3nbqlzY2R9eJWhCzFaExI2xPVrygLNfb2ij3T3Vi
6FAAPOPOLBHgekAOcG98xg8rksui2efzWJdK1RkYd9bMSTqO+jdLZ/n0NHLe9aaz1SDfUg+duJi7
QvvzyhSxEfzOqX/ENZX7YFu0Lj43TaCVu0kciwZVlXHWSlpuHHWNfkswNVgOb8x9lHWsZAUkNw06
1KPmWSdPjgbmN3HnCO+DBuZttUqRfYmtVsxe8w9TQ5NFKYUK/LbBz/S0n3dEdUg43VA1TzwkpVuB
kVtAPVQz+fNKzBlPeBf0bKPtPE5Jq5VUNoK53YnxXo742H3nxnXuznD3JEc8opsoT3cFDMqza0Fp
bWbqCzXHxdcIB0QKblAmGeGB4TYzGsuEERRijrUW4Cy6vLBO1hZza+dHHeeR5XQnHisaGSejk/gd
nJce+RXvO6lpnZ6Gkk1Nuqx9WnM/nflV5VdyLo8EqT9ioLyiqv1DTPttKq7/wQj0Kh1we3+Wc0H1
s/nsKZHRMwaB/cXE7iZTFqX8YmC+AWlgh6KcH9RffefJpyIWA4rxoZfxTeIhHA07iIFLKKyJVuGQ
PNwj8CarQNBkClAPbn/m+8z6NkS78o17MRdwUfbYyiPO36oWGE8HibAUXpn4I5ZqCWB3nComenkO
FPecffaA9QJJU9lkbXUsNDeLwAXQa2ynXtLmfSYwWzG2UPWVd1huuts4mHt7apE3Fq4CP/RL+oF+
K9J3Wri0/pFRT9/l3uGjxFfu+sxAP21BKKwShOKGJWA7J39pVn7z80h75tQgP0zLoYLmEa1UoocJ
VI/R0xBT1qmrDtcYCUo4YCanfOgOjOvDsp2UkUaOQvDDNMyM42t4NuaTY0F8i8PBImHV/H/xLjEH
zHzUO3RFyC40IV/rbAE0LMEV9KDuW1vF7BFNEGJtkphYyVqsWFgQEaN34TvTPPxl/fgcD2TAXMD2
Hm0Wonh7YRp8ieTvD8pcijglTtmwGm/SbO+E5+iiyHyM1ZyRN3ZdmxBtc+8U+7ZDa4REz08yeiO0
S3XqCenGx6pmpOZRzyWFvBJdrLvShCU3ejQv1xhRr9tFZCBDUgrT96Ht6WhMnE/HfokK1Hl6Nr/+
WZ8kiJ9pXH258L0RRjRXJF1n//AxTZxfcJ/bGBtXCTHDc4EbUXmCIJxQUDbTNjEfT2hHNng74tay
K7GHll8n58zInvyrEVAqIZXJ5IDuvqBkg06kIzGsMw29eqYuSIXx6jySryQ4UEgOY4ihbpcLz+wC
c9Qiji+tjZ10XoL35+huy/PxlenOifOZccGDOqC8S9+5sF1BkYUECsI95QZSAJQoMoM9Y5ioxT7X
1owQTMb989bMWczaSNMw8ripfukwSoJUitK1mWH5n10+syMSg3TJZskFxQ8k0ZSsz2TvzLuITdKz
fUngAdyKAboRAOlVVJjMsWz1RbScn5BGuR2dRZmEd/O0EZTVG18MLNSOa2xdsQu+VUNsTqVbZjIJ
bp2V25FMCn2B4nujLEdP2VLrwByaEjgIqB3/nMHc89M+cToMJT3ejaCvkTXF0RmDwyk0kK4/+vNq
n5GjQCrA8U6xIIDQYZ7FgTdsSJtKqiWlpqh30jGkOVHvpVt49p1YppAkuzZWdyd95RcVQv0mdJKc
uvEcN9RisRlGEwzD6HgZmHBgYhjFxSItD0QWqHsLxEUjJdT6fCZb+/Ce/XxpOWo9CiIWmj3xbrDP
v1UHs9plzUUVuXbqNJGKvxkuHWW51ajzlhdRtTGMNQGStsDA2z0EGp+4pKkI16ptL7hRbW9si1iW
gJRxzjC6hpm27ab3hoXDk2ND0szox9p11SoFPBhjzj0UFx3/3axCqytmYp/HGBGemRy0DUhNXRLU
zFEYYUrzCkHtl2OjjOVOz3Hjf8soFEJPxK7HT6YQwkSR8eIEX/FGByno3ySL2/mEtFB8Ohs0W/+A
gTC9yWY9XVmgDjgzNdlRhHhE87PZrmJJjf+Al4+FBEOzWocqY3nALRAzlML46XMX/15UJ/Rye/DK
4giMeN4CZoZgZYjIf6qb/eJaSfRK8VPZJ//RJTMsT91fubM3wEmt5aop/jib4n9E6CoGVxYAHRQX
+dE5GuJB+2UwDAbczPn9bSZqkwgLEAPbIvMUen43YWBITN2bgij8QKY2FYVjWv7xQQ8lmWJQrv6V
PzWRZeJKTYtxcW40H6CWGmhuCCITCWFWON91Xk9CeAbEKQgaHuOF86+ex8yZinGtPZumzLOpc5oX
OywI14GVy7g7qy9yedVGEwoOEQYOIxclV6Bk66QSHzwqkXPWO6/UaHQnKuiowokpbObnJvIkk0f0
XlT8RIzh6EInOFjsuKza3HcxLYubBOdDE6xEaw1aNpzfE49DyjWaje2FfVsz7EW+9mH9qk/7+NGA
Skl0gRgmMCd4A9dee8oiHjszfF+fTrdNP5+juNDQMDg+uDw0dIlyAWM7FDrzigL+LHnHwmbWtBXQ
BWYTcAKpSuIEfQ4sdTQxfNAlTHQMywctWPU1Z7Kz69t5ZHKlrdfP7Z9OZGM5n7AZSU3IBeQCw4kv
Ym+wME4YWFdDMevFKVrtDR4h76pmDietI0m1199D/mKX1qU0pbktSsmAcDrk5CbdZtgcJEXt6iHu
r68m6lJwXQKEYSC9afVGmqopIBLc7LY+9yBUMz4PH5FvT60nwBm1itOR36KeJUhAPZKXKVz6Vv5+
yWrQQ6nvYQ5GmxD2cR4GzwhRKe6A63iFS1yhduLrelDykPnKftBGtNfqLYlRLG4Tc5UvpsQD6dQq
rCvOWJGvz2dbQcQBijwW2vycLn83m9qmuHJh4ENa3oWWUwpcaEqOzmelbVRmEXhsLOLPqAZafVKz
rChBVa47OBCYp1lTXQgUiOe4MxQ1o+qJKwj/Yfvrg9zJ9Xjnden3h5dsaO5XEUQk8jLMvdyzAc4L
pQhdwBaqY46gyVHF9hsQ+rMt09gyH8wEmPMRX5nyHLoW5R9gzWKhCC1ljAFa7UVT68GPI4qvsv3V
sjH7Kbx4cCw5+tG2+CWjUu1Jg5DGhchiWxqvN8ISZAmLuV031cmPYfi5RDoK6l25AMnmYqpIG26g
GI3oSdRE9N1AqXRkkdIQPzNqmNTkhYRAZ4LTRBA4NoVD7jMiZTVParWQYWZP9PURkxyK1HlX0tGo
hj/Rif/UqhlAG+7h9QuRctyEO/XJKlGJr98qudp+Ua0KfzIy+BjXj99mA54CdHJedBsRzJkmPrQf
pI0ABwsbZydFeOoBS958psm3nzClYRsijUO7dzKAz9+jotNd+OSPuU0Y6EsGO42IJH81z2vePKbf
991C5EQOS6Ou8W0aHIir0hFLHCbLRZSZnG1qVDjGIdV9Xd7TVctya0w5fXbQ9R6Pw8Ba+iGx7dQM
66o2TWfNi5Elfy8X/9ODyHXpX/u69ncar6n0e8xfUdFaY4usarguHj4OSNP+46ReNTWCBbNBoFSS
zFjWsIh/K+//E3YeieMQo29x/PtFmMDvb9oAVNnuTlKu0NT13Jj+U8TOtrT/eNy3hFDWG7xgfQjg
Ac1iRFPNjDSzQGEZevCPEFEPq3gg32ZJb+5PQBUfpao/UW2mSvtIIGjnI12MvUIRpNyrqz0f/efs
9gz/PIKKHUWq5JB/qQ9dhz/Vghor7zLCOreB4MwnbuG1u2dRMQa0S9WnJWtYrXuFxwiedbq55t44
ilWBCZe+eoZJkGGP7DJEc7mJz16hw4OhblNEUMDQzsKv1q7xN0OkIOOLxphmuG3DkS7VjvWT+u3L
+T6R3rJgZDoohpNDFamBYbB8M5Nv1IVAWbJnNPn6Fz0+b1zDYWceWdvgX+Q/IvCv+A9urinzA8LN
rwyRieVe/1BSk6/Qowj5BnarhpnjgzvGSd5WgsJt3xN2nDiao3eP4198+En4k878oFx6GioCrmOY
LoWwSQSXlH1t32e5PrLsevTuyPZY+ge60q3sx9T2N2+HrIgRAin3HltTCGJzlPPfr/Ng7OUYgHvu
lwT/8PpGO5LyMnO6KyFfNIhIqLX9s9K36rBN1qZiIsB7MSjaxJCzspsEGtspd/EjFOpLJ62whKYc
pFHTWCiy2pe5C9SWvk8PU0yeU6wxDU67LHHuHTLMr38UyBEKzP8dvg7yKtgFiDXYBbVZWoAbFOHZ
nTzzhVSnt7OjIF1092HcZU9Pc/IXVjR92oWEUGSwXz/Bm11W0HZ3AFDUGcwnM3OlUsZhgbLaOcVQ
LCSYrrRdeEzztaVoAsa2xuk6SRVJ2KlTvK+19/7Egdkn0ft1AbfoGltDlPAEdTSKtvH6VacffxBz
zduPKqUoV7Qqzk7/HblZprKcCIVa90t2bhuuHaLAL4dEvvDb1xnTN9fGkzlNaJV3Rq6xQ7AUpAeQ
9XDRyeapWo91uaSUt0hStv6PdWP0x49yuCqshVPTsX4ckYvU3HNW/Q3pTfh+iqWYW0svvG8z5CSF
hLAXc/pJgTlcndNbnDBJHAIbRWmL7sZDOlfk4MjAPJIzgOreBW30g0JkEsmiGHRWXmWnlE9PY/zY
Xz9gKrfCz6vtM1vC6imsz9ADHzkHj/vFa/7vVtVAdfDduVmk3xlxjF8Q8NX7OF8kZ3A2B3QoBiiu
20+48Xzpx/yOd7DxMouLgNMdR5/4HARaVHvx2FBUh6+KoQ6uoExUxKgEtd3Qn0k0SjKwDwEO4DVC
7AEqC//xW0x0FMPCtnJ+KU13i/w4hu8U23M4NBt4MUKUZQLbatn1lDHjeGGslPsDnXdu9MjtvMre
Cw3Y73q8iCEUXKAEu09EpQu7MqC+Ltq+2JaIeosU4OsgwUr6JI+luryQXf1YgQJg8rEKmlrlig6z
dKm/FRsFNq1EZnAdCdmd6RlI5mLaaviBCQP56rGTY/gx64WUdRN46yn0p3r9iRPD3ZNUZQ/+QxwB
Al8PPmqZc15jTUqZWx/nNcobzI91Lvmz37f4OwYDt0W6c2HJoSPVgwRbrTbjh7cs0kDZfI1hBRR+
KvKFek/2yUZfZKX8dGrJtmjSAzkjpkvw0j6V9w/qYzkMcVZQCear6m24TvCJC/QXCdj0KN2P8Wa1
SfGsz/ucv/4DD+OoYTggSpa0dVah57K0oCydwbHdg+XoTLwQJBMLy0jXsjuXxpZbDD1fV1lzElAO
xsLlhfJPK75pZbI1UluKu8KlexWxTD3xWzX2ZaDm6Pt6ioM+H5gtxCQfFyidWfI+VLJY2AdsXsL0
pedJkQDuABsOOgEXRYi2cgzHNamCkHkXYdFaa+7alquLRdjy7Exn1oQKOuqvw8unhDXx501g/qu/
bmmoPneG4uhRBn4f0F5RjR0C8IoSzHUUrW2mpBZLOVYi0L3O6zXW8b47KtIn/xtsVOuPh0FSZqYB
9bj/Hp9uYiNNvleGblYinEiuLsk9CxTppJ3ZUvAFjo1KVFmDRYJExqKH+Jk6RJ3x6N+syJI2NiCf
xZFNjXs7/5LHilfy9xDdgERU4s9eK0dQtpD7PZtHcT2i3fhKlagy44Iz5RKEAneJcgW6Gwh1LKMz
7q7Gdk9MjVwlkPvLjwVFotCtvZE00WzynBtVvZfWuovSOJhm6p/Sq32F2qSQ2VRrTIHvtlNHneJT
BjlvTOEm22b3cibw4adPrhX4pBFvlTAs3qEZVZ8x4u/kuUxapnZM0Q6zTGCzG0ke+8xn/G9bXImU
DF7SuFrCikSnlg7qLSymZSWNSOdHkXPn3JoTCTdUywnuwpiJg99PnyzyGAkEW1iOQzR5meKg7U4N
GZ+UM3wVN8xLaD2GlQ/DkwNUTHh1nFxsi/5ngOqf7P8C0q++tU3HivCF5e57jAM81Skr8CHGUldW
cmjzMO/Kkg57XgHb5jPrawTt22PCvsnvKCeyH0yVYStEae6kkZzONOBpOY9HJtkf83uWvsWwIC2t
encM649VDUDheOWKbVt/oTMqhu3IIAMntL8/B6Ux8uXBH4e1Yo7p9KhMOUVGrqQk33louJ3El1wn
q8MJAqJjkNF5Znz1fOksmj10ThmF1iiOCACiExiZkam1RBRyblqcpnataqtFvQkkZAkfZga79ePo
SzY9XigPyU5TKIciWDKhbyPewRPNYuqMHvsd61jzYlt0c1iFYCFfHUNnMTbMf6rMlBwe4ql0Q23J
TSQ+SVLnmJxIdAN0z/7nWzFHLlOVdrFrI3tBFlW6oQ8AYVFdTBOQYlj2cp8mwlhRsw+9ULcqoZ5D
Iln+oNUdVUoAA8I/JQGRVsaU8eT5V03dB6wjBH7iCpUmTCc98HX+HIzc9dh2gUz4edCRR1in6+Ky
QIo2GvsEf8LaI/OjmQ/avcHtuplwQnVwK/5D9mkc63y7kOLQUkBRz1X7Xq+6m8yPN3F6wqz4uC6L
ib/GxI6Zhy2C4KOo30kYSbUXt6UBXfnu3ikCNG3Lj2nhJyv1wquNSZE7Rvav/4Rp5601nm+FenbO
G9i5GAW6fBtna4+mR6Qdt/KXypgZAWDwyINqJ0ugiBfZjPKV1u0uBrtxgpftMS+O8vAOArGSxMSX
oXpbr9hNDsR4nW0S4pxSJqKcPY+Kd4i5mGpO5YmkL79g3WApbu0/LSeS4c95gl2MYkhQ6b+d4aac
tCU6z0tlmVjexYat+h+gT9gSPI3DGX7jwK0X+glcTd7aBgaG51Q/e2w3Iqvh7hLZKt6kJ9hTKiEs
Rs+CynHbiTeAlfFa66Fe5dumh9+zL2NFncDIjYs+qVM2RnvrVW0+pB7h2HxCjnDI5nAdr79xWsko
8/FBOXCYVth/XxpKrHAHVx0QqrB4dq2gJk+aii64tMeogZ/vlnwv4y52bUZOteI15KxoSq9HzVD7
urpP0LOKUpQ3FXaOTvfhwS+5so8PUUtFsc2/Nb2L79aIgDeQy+FuEy6p6XSzIS4lV70EyuQJjAko
yKX8boX51FJbAt5ZyoF25BCN6X8m7tbDsLh4CLIxWCIm+gsjYXszMYpseojp9S2TePumFAoqCy/W
Jn8Y7wQ7H3ZzweXF+hZUWfXkEka6kfxOTpCyB5cmet1JKX7Jvkb5+YrJi1sOUtHPXX3NLoVhVuce
l47FmUOf+wiO7N4d4ZivCj/ubdDcoamRQ1Jdyi1/SMw2ZCqnhJ9YovsTy95SK9mcOEx76uenmrAb
/xKqcAvAj77cJE2vkPB/PRGzS/cWETLEKpwLxq0TyYmKnBRrh/uoPqDztwqdRnSvik6NKGstHAMn
W1Enm0RztE/saWJwG6xySdHmECgomchJokbL+dVXDhDmPl6SQWC8zvsn5QvpwVfNtTqI5kH0esaM
SgGKmZDJjxmLmZwibISUgmJuaxV8Z0E5+D7yyoH+aOeWAWerR9k36XNXtlUQXGbdY5cUnmPJPZAY
CcP38qJS9himSVoJm5rP3gSAftlG95IQ0/Serq3LgBnZ5EToYnopk4HeABAwz+WofEoYj7hZWmhO
IwUCfpLjFl6vS+4VGtYyWZ4YQua7+4gIVEl7FrmPcZWYXCJQvtJcARPZCuHZvS6VueN3MrAZst7F
6Q/QRDgsE9XK6knrBHFFVT5v317wgn0qS0VFp6x3v43qbhUtZ0eNPm/FsOLaHvC6L+ca7AJ7Oa2C
dxHxEPcCISeRbriMprT+St9wkcBSl4GjTT7aKs0iKTU9d7DFe9S7vHZa+HvKdMdweHOBWhNaX1/9
TxyRjJyD9F3V3w/cKyTCjltD63sQtbfKT9Jn4WCfwH8ynEhKnRFPbfKrDD+b8ZDWMUgvkSUE9Kes
eh7+BAu4g0du4svSvwbxtPSE6V7lKtm4o6bSQ3LtMics41zendnWGCVoEgXU6P0B5ArYFpQRANuR
xcVxQFij+uU15P6nUkWCg6HK7DeQhJkc7+32bzVlCW9YSd7ofi5T8V++hC6QRXSi99QergF71rOz
cCbPG8IhChSi8cCdrC8grgnAi7GukSe7JXmY6ZKAi9t/cwbJcJjq5zzMcVOZOzotITfBZCDTkUow
J7PIgBHKWriBy1QZRdcZmOv6VtgNmcrGsUUVULaLICnxC5OE7NSfnn4+HF/I7L6vk8cqzzejnBOZ
bHVwRXvtniugc35k9HS6pWrnZj7DxewyyQGmSm7QZW4ijaJMM1TmK0L6eCkynQRDiJ8mKjvV2scf
Ub46zSC62jbBh0gxpKSDPQCynf4WrM+SmSl3N8M+UrdsuwZSVe1yQpXR61MrPGpXOC1LeyObNk9+
Mt1C7JYn0Kp5zQzMMBQCPd99sBHLOh2qSd+MjiPPDhxbA4fGnxg2Stgcj2hSyvMvuTZrFYuw2VDW
w5IjD1p5Lm76w0x16x1L3vDCSXwAosjEF5IJVaA5Tncd4zmX5m1MykXFL/0j2VI9954NZUBZPysr
L1FcemG0QPydMYt7GbEE0p+j+Duvhi7VWqgvpYIfd2T8FxzzkOorjDPAn/uzoPBhy5WK78QCjlUD
2oE1qQJG+NY3+OAq9Jck2OUbbFqIAaZms9C/qPu2OCeB1h8gOnNZIiivcrhGstRafG5HaFkl3lFO
42HfEYnLvzE3RsUB3awZBBYv3p9ixG8lJ9WDi2Hbfi8TNsxH/lBv1bVvV7gLupdaGg6dNi9PkBIS
O7jUgE2XrmKiJ+YOdlKGvXa52kEIsZDU1M73wwiLYj2UcivkWoocNf1LFwOecGsDnnxyjdoxIIGK
yd2kBoTHn4YaLqZSl0iNHLDmQPdXDc7I6OoOLbVnaOUAup2rOknNIZVCfxnMV2U3gCDgQHm88BbZ
KY0H496cmqX1Wlv2tNWh5rsQEYH5gzlv5x4dHh18ewAYv0NIfzFkzevVEInS15qMA9s9PzBRldrj
hQDpJ6Ic1LHd2mNcblDjbFHq3Be+TXn3auzkMkOYl4puCn/I4iE1weuv8VxZN3H5eNOhdXU6cLwf
44L0ZyWKq22WSn3UJMHfXwOZV6tB6Pd9d0NuGI7F7JfsOB/e8WGaf9nB8G4B0Lcs+YY5Ct6XWRBf
QQLjpyrrxjHaLutb6m9A5zaJBpZhJVukVk/x6AzTZ7HQFQut33wOlS0MbsAle4f9obldyfXPCDah
yQzFph9RIJtZf7RbYUBlyrWvklGmKuBJrLspoinQoO71MwRb8pPzVQIRsUoEpdXhEp9T83uBVY9L
E31GN6AeLkeO4y0a4Jc/nuBJyof9C98vsWhSthNC75uGWhqpeNMxFaQs3RinMfn9mJK+zpgfUKW6
dm/KrWSYu2kwC+pLGXJ5bDdaVRyM47qneaw226W4lEB78XLOxCqEt8Wp+jk195AOwpTZzk1wJaGg
PuMTJJsWmKcWEgUbvPcEKdgORvCSf+Nv2rYOrVrUgHKsbkucVQUvUTaz7Oq0Nopxbis59mfg2Zdp
y3GFaliNdOjYJKG+ggq30cGehOUV3mMtuRoSBGxfGem5wctiXRVd7bxHfsBu5USuuNeQFFkDIeYL
7whtITgKyoUVMx47E/dwEi6woT77otGPKaM0U0XpN9PXdEgt9qQlKRkeTKLkPG1d2qYttuBg6yBs
yyYtMrcK0pYTdRPkOPkvvEbfRwj/DnKchNEQSVOX6PEIpnRebACDb4Og4ox5pVy60M4xIKWZDNSI
D/YTaYSN2JyIrSePCZ6LZ4bMjIYgun7gZEQVpKSe4eWi6X8cdt6vB0WWrAwgZgIYD/EHDexccHJN
21Oj64VMIfX9+pymdbsd3nWUrePefe/S6v8RqamZgughKRd5i0ieamoDvw1kKpFdR+FDJ4u8xX8+
02IajN0Qk6zNCfiQTCfphD5YSpcutbKzZCQ22YpFYFQooHXWgGR/7iF167oDvUNvaFD/cW35Q67z
xPud4RT6et1xsOLCvW3GQfSG+7tXd0q3h/oS6pjC+nHrC+hnlivVH+ovQ8wr4ZPovsO7QdKgJ+Xq
2SwhRVKRa1Vdc3DPoVPfOJSNz0W2Yr46sjEjEGzsc5UTdYp/sUYCnggsVbmPnvX3el2JoCoernqZ
wwJx72DelhM8D9+M6OxK5QBywnEHtH3L+W94ejUOeMKM8BLBEkHq+L2+jnthpnKxRGFS2bp9DNUH
s8QRJ6Au7cVCdC28h69/k+02y1MCJLTFtL1jFoSpjl61Qj7Hig7k13mzHy0alEeytXzHgPVAf+Wp
8H/Xi75JV3uILTC/jCt5jugWFnXHEAvCMsiw2aWIQkq3tcJ00M8PUJ62ojLvSfi2dm6SmziTlqHz
4wfeeCsL3ptFvpgAQV96VKYN6wKl3NcGVNDKOuZFkfYVPZEqoh5Ge3xdquNZW6CVYgrGvE3hVEmy
MSWhytBC2sEqXNvj2KcJ7rTCOBPZGY6CqVJ8KrAkleGGeovpwMkb5MJvbogVdzYA1rozlaporLTg
ILcS8X1Bl1YI5+GbTryznpodN9+emwIlmG42MeyoWH45ZisBvXDsfMSTU+TRVETN9yEDYrzs4JTL
L3ndOOtzFBxghEQCgBKq4gLelg3g9fGbJijgIlDiK55HpdkjNKa3GJ7oJKbZpBWvHtk1NXwzTDUK
Ptw62QUUpjLHpl7lHOdbKrpYYYfejmsleKwC1q569VuqNVX1Cm4oQpwk2U0Lh7lW8oHmB6yd+jMP
/h03NiXDosEA2kD5Z2zSsm6/d3e/hqzd6PXxRup72VS87OQsBwGx5PL3IURqY+MB5gQq1GnGokyS
yrSiWe/ju/bQXWXRbes905TsiDz/O8nBN5QcuGVJm15F+o+HxD2LKZAxXN3xXm9S7y5ZYA4rUFFq
DfeA9h7kiolHSdlACMGr0voOIpj45UYZ+e6q/q/xQ+DMKPkvmhc3n05WqRDJJqRE4On/pmkloys/
X5S1cAjtBM+e/N4GirYjBGPZj51edQq/hCvdmWu//5riXJH02yPPQGu2yLPPQObiU83kKSWiaeYk
KEfK6IuMdfhtoxoHcRtt4tUyan8QhWNHCBaPIgyzDCsYBT6hCDqKFqoBg00xboSTx21e3KHWqUPf
TS+DZ4xznG3Lx4HPqnSHQ+Ja3DK0JW/4+gWZElKuPQeF5f/sJXHx+FroLAXc7FPjIfzGevHyEIO9
tUVWkh2KMPn7VvaCcSQ8ZmK9/4T4O5k0IjO9gQ7netTbyCqugR/Jfr6N7/8h7tOSZlfa03DnAUbj
AuIp/19JgYg947CnxYrS5T1D6bKykFkb/IDr3mIuSHrnPJYuJi+OxrZlmHRlSGvG69uGETeQN73f
81JEphiCJUaZXqHptbJYmuSwIY6s6tvAL+33cQaj8+Qj2eIDrwPYHwCPQdrKnllbxIaSZgMz9tMw
hBZC4naovH4Jz1hHSwWvEAPIaLBTQmTE1SEI/buHaz48m2YbS+X3P0LJRKxZ1PZ1vYRv2+IEWzFR
cgJ3HGEESu8j0rUJkfmUEo4WL2jthFalyADS7ts1OS2Jd2Sb54K0htkDi6HZx3QYNB8NpkjZsXwQ
Fkv0NR7Hz6pEvjO0M06mS0mJ1pfb6LbI4kGWbXOTRiVkRNb5j9OnfdOZx9T6XGEFjGKRwO2ZNW+v
fwsz2DkQj1HfS8Id2+93FIPQJ0i+4sESV+z6mm+SHx7dVOVq7U6ygaEAvxWkVa5k8dH4+zMY3Y5a
gdAgwzb6G2ZgEJjLu6yu7iT3nMMeOjttTbZs8nrk5mDaKtgRXdlAi9nuu5JGcx+KkxOgya7eR7IW
ui9AfNUVh+XLHsudeemgKz7Q+TibeWHm1JOup+HbF50eVMZAe7t8JQuqzlFWMVn0Vp7Aro3e3EiS
UzXyUA8UATWWqKHqqXjq99/+1VQ708jW2zWZnLuu8ZrqqUoL46cXQgBvg4xgZijhMPoB/xvIC+mG
TPGOjbIf9fblXhUiRzuXe/dMSAvOqO6bnoH+lz1n/xAs1umjCrRkyJKkeok1oYejORVdj6eUfRSa
KUyfOo7ug7WSr/MnzmaIy9FvEH7Szb3FjP0WJ/IlqaQN86RNkKihIlCZtEDxhMHBbJinfRIGl651
JPdSMiiXNmbpdoY3nazKcDfFfFGjsgwGOkGb4z20Kt0+/SVPz6mG3zwlKva/PAohCnmNWAqKyePm
xbZdP84VEPauWTQZpeEscMhSe0RsvQzZOsebJvBnlT8RCRx78yn5+SMIrInCo/yKNzPhNz8JgACr
vk3dsVqKBAoz8896JUe7EcEzvCN9+atcvqvv9EPHgNcqIVnrsa8lsOvC8SNuX1B1J3Kk3UBLbo1b
Q78s5bfd7GE9igaH8GQyopZSCu1ZGwXvKE4H3E0e6duZJISgvgl9MMV1Rqq6BBgnn7crYlwT4d8I
B5ob8Uq3NhviJVM+QHPneLB9Xv1uKF8s834eBA35G25R+ouzaZseIg0zJcixVSdxmbx92qaAP2Lt
0FGDg6u8MWqqNzkduiGSxiwGE+mrJF6IKHBJdsNQ8lK17qdHdSZWp5x+eLkTKLB8VMJqJKbVOy+Q
E5KVdFeiOESFybf/FRH7os0H68Du61EXL5f7OVaEVdRoMZ9zbueFeJWlKOPdyYGRhw2kQmaBFuFY
4FH0PNlpNad0Ee9Uh/hQoXAo/ec6Cw0lr97Ivsib6feMJEEHUMJzvy7o4llXiB0p/TCTjXkTDCm/
2ZspW5nKfXWlKsc+xw5xOrEScQG9Y9Ms+vXiUjqgSV64fMFzNqLMWJN9KemxEP5PhQfGvHrGDnf5
lCx5ztBy9vRFRxK8tr2lvj60tTpLGg6WytrfZHiljYdYU9LNTv+rBUT+sANBOtENwcR3hfpJqBM6
/igd/2F4ZqwykLuXUXmRlhFlJsvUJtjl/66N1RZttOgbY6YzlksCTd6uRuHKivhRdt7ugCJ0ZlRA
FZlmg0UhCN4urwifnXnB9HkXM4pM2JDEd2i47PQTWScEDS7tWqp6prYn9Bwdq1RyDHDqkibr+bKv
xDZgSZZ9s6gNjG2Sex/zELddFUzgqGEpxwf/J+U+SMTcpLXznHH0yhfDrUaCUwNlVFHSsteuHv+0
9DAZv73zGoAs9Cp53oW65/mejgpdmo/Xc1SEReqpHyfD8ZANTTn/n4DZOaSKDt0jgU4qR2aoNmDf
DT1vmSCHAv59mN3LYDxgmO5rKtaJbREDmKB+LkfDI/YQc8tRPwa7j5KscX4OjM4P8ghFUvZbNHT1
S7Xd4wdjrCDEBfAZb3k0V9Wt8eLcHmOztW9/zXJpJxMfDP/mUtHD1BO+F16YJ4LoqXql8IiceLJq
5C2QGDQK53icQaqmpGEmuSHmofwCO4sevmImLQvnGJz3kFPJvlR/OBCFHRBFqytl8RRmb54oaLNH
3Rxu3udapLqJT7e78siCbAGly/QTFZwDpFwOosBs4p+u8cd9f3iRTglIhhIBWu6AL2zsvCHjpSaI
2nGcevqtemAHXK0BiDB9nBvRCAuntF5f6kbp9v90ViKqvj6AK3ZNAiAbsT/Ym9nhFrQApcwX2ner
gWiCyexJ+fq+xDYz6js8gTeyStL5xBxChF5mS5l7Huv7yNpIQ7QZK3LNJEoTmjh07apeBykfUB00
j1+8At5SB1wtr3Dnl5i3jdgEFnNdPPHCTgWCmcVHKor4E5brB6inEeo/G3dxlkEhk2h6TVQqT1+h
2r5FlX55QM2ir7LcSkqENe6aVqZCZVegBva7MuUdIylFH068L62L3Kdb+4wePK36WjBZGlSa6huC
rdjzOqeCh1CRIa8lmFIpZdXvG0SDWJu6ANePt0siCP6eIcyfyQsGpFwIo5hmHEL5V8SJAX7QIyBI
NTi2ENGQn24WueMEpmUD/gFI3uZ4xuRFT7S87Fz0+P3/C7ic54sWddf4AxBOqzLk2Ajuz61qtWVO
KThp5bmcPNGlcRvEQAy55xbjUiH7OeMXVxRLm8QpHeNh+eI7QaGm2XHTZUnY0lY0tH66MvU9zTg5
NXz1fnbrKKtm1jT+Fvka0J6vEra0dVusPEaZx1PIiKiROc1Cy5RT1an5Ubtu7NJqUoSFabxnqKer
3PQNDHNB0IEvguXlwe9JN1mIqgDzS2nr6TqPFRfDjPCrtCq67XCzqfBh8/R5WWIG9eMMq8XcNlRj
3HkfMce9IsSOe8KzzggJtkurekvHg9YWooQw1iXFTrHcZqLGw93wieY7jFb2w/BA0Hmbr3xyL4fR
RGKfLWPjRERom6FaokelYk9pj/Ltu37Ob2ISDLvoPvH54mPjpNjGWbYgPYTgEj2GIikMa7Byfr9A
zNr/KcvXnV8Rtelf1LGlnKqF99HSCebUAx8d2agnrf101j8bAYcXbEQnoZ9naSy+9nV5tqLqwLw9
WEOa0SC42NL8n8Cz1KoaSEQCDUlGPCeKh6fAfiGxA0XUgyyOMsh87YpvxL8vGtm7OmOs5taggImr
ucxc99C5WFmdnUJzIA/lzgbLt06tjwNco3P/oxjqQPffR7ZQmHhp7eCWhkhEyoor/+H8Rf3op2qr
RK7WjI6yLzSyCBtKehZwhD4qYpMQ2hP2MGKOnDoPsQtptD0/1Q5acYvUBqOMLeiTRcCXYw6Y//9X
kSQ36Ka38SRhd/sxcDu/Og+BglN6TIGt7vrQuto7LB6519CJV8qqI2M6p6fGuQFdbdIn+J7HowLx
dCH0SHVwctEhZecV1PmqZxG7lgREQUHZc6aUMROVxDxa4nC6SxAGvZq5UjvRki3KTpVhJFREQqyF
irqV8m95qvJPpSOnHxnLWkuSv71o8Cu0TYa9h5wcyNFjuNdUE/ElgE8dLDLc8axVeqJh+p9hfGBq
3Yb8wQDVCUtvn/UQWOufvcLBA+CS0mr6xwnQuxjbFlB61T7rby00wfleEmwV1uYiIEthGPSxK+2L
Bk4hOTFryyajTFABDkgQu8CQ/t0v3TeDcQ0bsW7LTfXgVUXxOGvFwwYYz1dkcNLJ2w++uhJDeuJQ
91Vxg//oyycfith1MgXAxsrJFH37OnP11375iUd/VvIzHD+8H0TWOEWcFc0COZZn3Sqk9Sru6eGP
xoMf7ablFGoLMV/vcfuITjPxHO5m9D7fYOZgl8GH8r+Yg93pPu2P86PRq5ZIrgiZbjkZse1XxS0b
VFmheVAgtpB6ggc/8JwRhS/MlSlnIik6KYnKs3LB+sNKMEg8hVQ/4qriCJBGqe4PO0QL9jmPP//z
3Hx1A8s2C0kmFQ0oTg0Ka4RJ3Bp5I1yU1piIUy056lph2hpmY7hGTzqOTuqa7aGq0X3C2ZF2W7jh
RE4MFyeuqSKupnPHQaIGki/gqaSABSvepRRgjnxKqyZtBsPRtJ52lagu1kKtNCzIG8Np2lLVEB18
Eo0Jh0FfwczDFff+qynMfZAMYiom8hGtr+LdGkjQ/nU8ulFykyJfCVHaPAkV65+ZQlu0Ie/BAxmU
IA+o7rwF3vJQen/B/QEJe+83yatCLtw0CgNUy5yMY2fdzpVFzHan3XLT3CwFKBaNbWX8FTfqPzfz
slssGre122cYpWQO6FwaDnctBsXtiKcsKNt4klE8/o/weFvi6n9wYmPGrFaFZtp1IxUsjVSpHrwV
iAy/HOprR+RAqBIXQLPNK6Uqvr0G1jCTwwB0oEd2X1G4YqN7ayxXHm7u4RsaMWZdII1uC5Hte6Eq
82T2B9MjAx0kaXQivlsg6J4dkd+73+8G5JyWlSZzhFYWP3kGHxdLcz668RsJbVcmO65PXanB88Ri
ATF636sCUu77Ju6G0YhKXvgq+QLY5ftYPvxdmDweABPz7pl1BNWHdOp7rJGM1qR8q/3Ylf3FU6u/
82CO7x+hOhC23w37OGLOJ164zawficKGbtFhbpys5q6T+2pKpHcQIGuie+41ood9BHEWztB3ygIt
BK+eNzWR0XkC7JNKBif+qZR9ixSHHOK1VIbcuBAAJuH4TyviedoMsnA/Q6QQAQAAxCMICber9wPX
uaW8S+HDbjs1bogxEbjrYNK1aqltTTJnb6QjW82Mp28jgeNVzIRAPL75EfRMzQkrzzaj+pHUuSpD
q2E1CXXkMKYL9/aDdFpynUt0jW08t8L1fOkfk6flEev+uv6whr2LforWb3jOsxssfu0tEUczRM7A
A8b2gIhDvecsrz5p3EqrCuLgR4blJqHTV8zw32MeG1bbNub+kOpgGoyEDbrpiJw/Vv7slKDQQFjl
ar4JdmNND3HY6WtkLJB+KVg+3mpsyNMe/MpO9f43A6VMGqv/bgdrgILtXYH7eJymtmAEhC0t96uk
FHmqrT+TwF1WbtVP3STNzlKjkfbJYUXXf0g2MOTyfbZiWDmFFto/SrdDyS1MzAmsQDCbXG4CM2lN
vFECgPn9+DXCPd3u1E8QrQp5YE+Ao7MXumO8UowY40KMwoG+VcNEnjkl2EXUqwwAexaUX6b5Nqvx
8To2/Oi40O+iObX6UrSgJipt8syAEQ56qDiYFW66uqGdQXXT5Cp16EPcFRbA82gJdVVokIbOt/yB
v8TIrt3xS2zwK99mcOBU2Xv7hJafFrsHIScc7bpcJL04emw61I1ULk2p7eHqduSYC5uEv9dVrzgt
UK/2ijkQ/wBfMwuISXlESj3yP7WZbxzujLC0hqhOm1uVWRi02zqk8bD8jIlBsOaTAP59ivwJC0iD
Q2x6ggmgrLz7kkWfvjOfbC7Anex5DRWehIPFI2ZoXCjUAydYyMM6UfsErr17T667JBPJoLw9WSN2
CZKyOAjXpNHvJxYOg8TT96PPU4a4GCUmJXgpBrRDXEhmvMS14hPWTaFvE4XpwSIRONXa4suMzq6A
BX6xX8Mj32GI1y5PEu2SRJYBNWNfiDxyfdLM+phdXhVL45wsJ8frDoslsiMibeq4Uoc9e+zuHP7p
5kths+HigLpSOMVuaq2Kyvn3JCKqhjYPKanBSBbP3wU3jSZUcsyMQ/ANfAbgp8WdMQCOOiJTkrbG
N05QZIS07axwGk5qejvttDloC/aA8PLHYVQdJEbffFPkLKrg1p/ir/C54HegLWtOAxEef8v6Ggds
i5obguRULvxQLbKT+92AnKSp3wzJxzwk3vDX9fkjbI1uLZeAKsuavp/6O65bvhNr3MArrD6wAnfu
JpJX6A1qQDgjBTglS5y4/shlfy04COOt2+xVa91GoMUfgzLirQ0QtnMFg8Se3wlx88BLXFtzWiIm
sl4fKPcsrqE84+HRWOSvxbBeQBMOY1jul6eXVUrGJPtJPWBJVm6bKB8s5CUrQs+4MnK/xn67BNwx
uwFpqYaOvdG8Skyc0W+c7yszs8ayqRkGmi0wo0x25dE060x3xZLdOhaaZv73J7+/vTowxTOW9h8n
QUm4kSGZB6XRsLfh3OcZa1Gu5jEZSHpr1zt0kz34yyYRXFcrmU4Rc1kyJ1/0lwS+ukCoRFOpTjJT
oatm6Cik4SVs50OdS53HfGle5YLv7JdVF4K5z+vGGrTNiiUEJEh3H9/YmKICH1Y3/48jDvSQz0R7
blOg02MYNGultQHTq+VtAOTnWfJYr40PfPerJ04oTpozo6/+WDUovYwSS9NGVo3cpgwNG2ADJNVC
54AVtdc50aZ6AuO4AnfJVkH+bMO4SnTnhnyjnzUhCt7XXGtA0tanC9kGAsNNfwSfMJaiYV1PZJok
0zMaGkwe2p2vT7BWUot/9/fx449SCbZpwK8td/SXXcmmWF1X//s+bQ0D7tv5cZ+OayJBxaydIKe6
dzJV+v40gW0a2kNwLBQIdDGfleRTMtnrWhOktQHInm8kwcrtKgGkVtaBa7o2PdyC9xpv0KRR3oup
EkNLyqs3llt4Tzjaq07bYKWdUuApZRmZZEBGjCy09nngKnX/Y91g8uyTu6g6DnICelPJCYR1jMdx
AdnjOyZvjxxBjzvtkcVOvfz0bwpbV0rBCv39Kww1Sy+ZydRGcfN9NgZqoMQE+Dmg5jN78RUZBQhf
Px//SYdzRWlAGBS9nlV1H7HvjC1cJxVAjw5BYWjU/abxysEPU5ls4TbEyM3D1Cx2HUdh4+jr4YM+
alaXNNsh0+AAjdmLEcTw3g17kw6O/GkDzgDou1SH/YEr/DAZnb6+0arKFnZ0RP5BAzooyWc6PjDU
HoKca3ry/0cecJ4ePS1MiaW66bKPBxTAhVi+Wg7QYQxaPKSvkOgpBsjfXXfHXPDccIqB9KmOES4i
702zXpUW7jR+SxKbJVIsWEgKe4fBHqHDomyd3TusVYmeC8PKemmCK/AAdXVQk3SOJ3Jb48BTnQTj
Y4wM+eIVnElDFalv21oLJ0lav2gjbuPs3Ub77EGQ9S5zGIgbJlsGR6S9ruEi5DyNX22RYdjYAOlE
AYvr/42AZ2FOHLYzdB69qqLqg868eUCpMX7IGC0ffLWRw5bnmfCkM8lKm49u0uBu7nNSEcfouXTD
2ZFdxw7TXoxYuMoe6guxofRazPS9yUmzGiyUV78mKcAQONoQ0M+BvPvN1jQfTVEra2X0afiBBv7g
yiAH605frqppu4C6mGETF7oC6Jok0wcRPNftUG6el8+soSUsvQC3WzqXxtrsOCjbV1viiHt3jXBn
mV03/hnhBEsHdlyw/k8sJLTwdocSiX/A74K7u/fkncyKdt75Vwz/2AM72TPNm5qH0tOg7mqkt3i4
oDvHDHo8zB0X9fOCMzRP3XY2M/JLGLUWhW7iZNBmgoMkhpRbOEh3GodWjXt2DFZ/mU8mETw1cdlX
4W7ujg9HL+5EBWOp+9/S97iEVM05se5shFsqcFec3oC/gRgoBqKpV7ixBJztnK+GYRodQAbqkVUf
sTQJFdj+7qKs0xntd5GHkauyYFR9bszYv+Ai0ZjKd+Kq1towjW202jFDyAW2thOKuG5j40cGQlAI
VxTj8JpNOpDi4LP4GCmBC5XYvsXSAIw8xpWZZz00fW8ztEPN02IhKMVhiAfC+SXTToIFC8xIbx+Z
+8MwE/gpAybrg6ZMSKyWvH1so56Bj6+70x9SIoeut/E3mpZ8aTmZz/Gqubl4N9W98s/fg1oGsPIK
XoNlAG04fFr1F6us/eJHdiqTjmwkCXArEfQQeDwjJiDMmaHEecB7KZWXZnrEDM8oAIsF1CyozvKi
4vSekvlYqiuV+FANDi0avuR+qU1As1Rco3p9IMDZlob6nPpnsY1dOYMPTp58yEL+l3Vb7S1Wahgz
k211eyTNq2YyNaBIbjuwLVqQFChey1BdRonCfrxtzoB8wOWMvt++kxse1SgkKoMKzuoYBjAwThUQ
fxXhQg7mKWYcXgJwNNeeb3/6YBYtaDcnODOGhFwrYpBIlvvhznHI72l2vAQNTulchnUXnSZw0TZ4
BMdVHKtI1QiiVvGr9Howr++pW0kDPtYPF2PcpFl/Ir1AhtcFrFagOPgKyn4gkhkPyuNCBBkSDltd
26LmxxBE/8VsL23Fj47JSNDiey/oqxkKrIXyfV4TC2KKrikIhcd/TD1nFJci0CgCNe5ecPt5woys
saFi+85vU+cSINfQigxs4CpufRkjfWivd3aKVtlgHv8pKcfXVWUSYhNPG6UIJX/PG01C+8Efpce0
utmTvTmyvOfmVSqjy/UMtsz+Uu/9NTmuxGYWXRkUNmB5gLKG75NECupzlsQDKO39/MXEUVBijsrC
5bSK/X387BO/WIksgbH93sGoh9xaT1NiHoFjiGaYSHUTIzdO+pX4FMbyvRVoiVfJ8xdcAeC10rZ4
KJ4BKLAOO0TxVMf3IetNQKQEvook96vENNw6Nt/IWngLRnG5XKemdlSXN5ntDqBblNcT2qO/GG6S
+JhjJZ2+XwGaqhH3nirrEL2WZimxGaRsIeqz2iCL14NX71l7OelfJjSQ6DUlGWweAg7PmUSoTM9s
Nqys3jMjKLtVrY7fiMWUrYxC2joN5O/LDfVRTjYmYK0y0FFNYbEzcRVFM28nHb3aCbbR4CfH7X1O
Ro/JKcjjYmj9br9JfsIcAeZMT+xWzx1e62ZXeTSEa87OvtK7g+ML0x0M+uocKwBZOu0XyCXNvfux
4DHYyUpzAH1Lv+6f1+3VU/Nc9sJYdejBa4DmtcpKuSEUdFLcV55wc4ECn+A9b6hyU3OoS7HuuSZs
zj7IFCNa2OVId/M3NpcAGT+we5rRrn2KjUGo4SVb0JIEOdPqZ/nNLwNWQbdyxriNdjalLDidL3dS
C6skZJfn1g7kbJ+3v2CPzAymEnuMFcZ0mK9r/qsgI8sGvdnXT0FHni8sOWsZimhSQRo4WSY/ynTK
jFoRVmLv13UHC5LV4R5GMtCjq9AWZX1s4XiflZ38s5zC/wLzb8BMkf6NNCS1gWmggvEXys8o7qDH
zxm1T4kQa1NTOgYiJT8jNrviil2xAkJ2qStihEa9Jj/uFTygocR9bKd4bXNXyJbAfNhv35Wb21f/
zBheMbT85BXH+nQ+F0d7BcarMWMzJI6P4AkCIXtuRzVppFsyWNJwoaHEzsR3WAxZRXyk7DeWVCun
RSXbcToNnOFDlBwL/u5fVfdLqe4Uc8mVeQeCYYaU/1EtrUYWP2StOSUStWZ1wQ3/N7hjnlj1LpKl
j16QlAh+kDanrebrbm0/nBDeUCf6FYi1GXiG+B/mV/3k8+yhz1HxOrlZ3xj0rhqsZ98/Nz40rr8F
7XlfJGN5qXEYub11VEDN5l1/gVbZK+DerOr8LQeo0Z/tA2QbGvMbJMi4DL3osDzGaRg80sM/Li7T
wz3/QhKJIYVsoN7tAevQNkTqPbVgci0S4YrrAjx4GfEiYlCzNxcQ1vNcYDD2yAgYKZlsiTpBJFNW
v21Rnrd20RcadLbldnWaLPp7OGKipyiFVA08cFX0eZS3mYzFXHNEobf7brVtCbBAkCXzAiEsIjSM
AhrlMA/4ytpXG0SN3WJWsIaT3fhqpPjekw+X6HtKifdLeOQPEdnMC92Q+m8bXdIsHrmAsdFc5nLM
Na/TbQH8tcUnIqJQo6FcoOvKgM7EaH75jajxbIKY1iZvhB6auOm/Tec0mM2QsHlCwmTGQGJGX54S
xKhWcDcmkaFbMo3Wdd4VDmrxj+/YCeYCSHaXzWw5kazzJ6B3tqTA8NAc+pmvZ26Tyw72HwWJqWFk
1eSajXEDudtr9Ab9OQJtZwH/u7OWnsM4278sU2OS875uteizRgsmZi3ujZbQWfai3eOAU4JnLK3g
Z4jg/N+gmlyBODNrGA4nh9TT6hDZfyGpv6DPvF+BZVO8mNv06NAqpY1tvAieDDySrE0IU2m6a4yW
EJ8onTOAhcmLSbHx0MgtqdEGUIcA6idrAHIpTbDD4yMgppRfZ04StNnS7+qB2qrlV7qaAd/0GWcN
PpY81p0eyDof8EFHwazScltJtge64C7srsP4/qURBlvbot6P5qVgCG2lE8HZbn43Pm6B/nT+xCkK
2bVoYcL+N/qftLXvpd7JDSeYARSVQLFJmJff3quM2jA0C4GmH86qSQcIfdvrogUpfODu+yooO1L3
kIXgvy1M5SczFUe0qz/hyGVSl/33uPWf7dJiWGD8bbhqPyBwjIuHbgEZKXX7s76DATBb2q7lS0sS
NM8MUPTNjI69XJyI/iR2aArfPUXFOR+k2tTN1freUFVGjJA7kUWhO6FWc7unmhO55DD1b6E+LCNP
wk0XXWJUUz/n538YFqjoreEnfz5Hddsc9MWadutBZ8vmbx7+5Q+jVDenh6XC/h0b6E2eU/M0FXLB
PY4GfzrKe/v+JsM5w0pBf9o7R2cqybmDQSGPWQmIxlZF2j536MYP+Cfv0YpvyGB7cof83qlFIBle
jv88nDdki8mhFZX9+eaRzJvKubqSJYeqLLyKxGZaFdgI0sCmKPNJk2MdzqTilX7xP9RDw7hc4jCf
DbFZrVZee30FEhn5jG+7cwf9PEhEHursCypxddASAK7np7tloR8dBOOzXWeP7G6tPE/Vj+w+vmKk
EggNwbQGjl/nINsa7/EX7EWcYslXqpoxKN3cNsgoO7nj1Hligb7U4b04SxOTt/8zANuN8rEwCtVb
6bU1iCDLaJmv0wdp73fhFTHCnlWUcTZNRE0XbZpNZaGl217LTzUv41z3IDzCxEA7pmC2mnzY4fnC
bTIRyW1EUORJC0SUpjsvFyYfqcxm/PRWMQb0UF8A9LAdVn6dxi7ODjdmWft3lZhnKy3rgd2yB7sb
6VQuzML3JXBKfPAl4DDPsjoi8GrNmVebF4odper9plo73UxBkYI5Y1kTfwZVFlfinxCMmxtGjEvf
m9Eny11OvVkZeKdGcbTscytQ0Odv/b+MHmT+a65Ndk8wB/0gJ15+6mVmlIVId/wxhdCEyVIgyNS5
p3OHuLXbTEgbJaV8G4y7V5qygcB9YAWyJp39Qg6PcSrqh4UEKZNwnKf3/tJ5gOgsLY34z0t6zkr8
6zWM42YOHsUqhQ9pKTXAZOu0QnAnW1VrsPCbNKITQio2Jrks4u2hPBUFCLGJdoooHay88kTuvsmf
geBANr7oKrMgdw9ywonLmfAFjrhazbyKqMizKwSKyg4bA8cg5lcqnKhgRstB8M1wHF8qHW9eUJud
rugY00VjcBomciEYy8OvFqZ2rwEX0ZcaSC+FQ5yb3XP85W/HG83ftL/ZfbdtN6Q4Ts3GhW4T4nUY
LyTYoqpOkZbZfhX+r472i6grLCQN5HBsyutmYTh1rDLwJxRZon1yaU5S8AinziZOzfssc/j6BneI
wOUQLGNiAZSlMZtcVuovskhu/1jBL1ZHCzw6cIM/Lj3lEtOJ3sfp81y4DxoTZEuD5sdGK/2gWsIM
ZOukdTBxS01A/qr6006YCiY14TIiW5iQCRIbl2SNXwnDFCsaggiySgntClGr9h9VLCxH101GgnwG
elmnuyPizTEPWbASgM5IPEH0PAyXsOMZjScJIyovUxAvNYzJO/tx/3NW0a6A+Nd5OPmX+2uW0uLl
i8csjlVWbGNuRVbSl4IcxzG2Pea55UdAl9iSrKy1OeO1bC0Q58mZYBYIY0k+Zsp31nMGnU8E4L+3
pPhNIJQBKfTkoJfB7lW9yNOdoruom0GI1ICYx65syjIfhmVF+hJIYZT7ALkN/VnodjVXPruPfIWj
1ileA3j/iMup6C/QdCoxKI+z0ZAhkKTJ5G0OBBvKR+qMGp+t8bC1bPQGkZtInuTwy2dvt0fjV798
5gEhc7EuZmbVZT60rAM9fWscTozruzF8XBvO0c4FVeUgcp3x5Xjyx/mz/n21wzRC0oGAvGMpVG/Q
XBdbOe8486hk/LtguKLC+JLy5Eapf/nRwOs9rcwU2jHElJocp+a9kS2y/JieAmOKNVplugWCGDyJ
B/mVDA0ZE8QOkMlZ6L5vxHPUxed30J2TdUuncy07sNLqxCbFQ9LpuJvXj5r2CY0MMOM5gqDtrafx
FlTmIJmPvfwUjmRuJ4W8JF9YiyNvtqz6DQIhmJlEGB/J4Zgt5zOiZPuXXN6oFsQ7ENj7Zfl3urHi
dCiiezURyznOYcTvvWJNOBrDmi9mWj4hdJWBzJdpb5SUa13epOo0l3IclLxPY3vrAjfKg871Azlu
IKUIRL8bfkVFEA9JjXFhYvPmzfNbSYicArHhK6Emv4aZPkozkOAP1mZlXiaXLv9iCwYC7KyCjfFf
0GyuIi2l7zggLHsVij7QdRJ+rwkAbW1VmvDjIfBMDBsXhoKLZkP99JSwFpm+kF0CAAIt8GVUqfFN
Pmm6HQExKL5Jp4kjD0V96Lx8HGy8SKGObp4+XUYaGbHeFgYdqMrhpdGH/E+uoIbPEu4qH0OqP+ri
yMztBxN8oUt9/BNbhsi1qbQ77ULh1t6UNFOFHH+pYJLreGShIlP71SBJWdjT2x3K321wJObJJ3sd
pshhM8wHcxBDu3kVo2XP9it/MH1ZecWVPspXJGGujVbOufzS67BWtrWTKsKmcqDH60fam+lCMyLs
Ft0dUpQczhsg/j7us1LY3gd/FpYPzVula/PgFA8KkCGSny+2EGuScASn45LtO7EIMU4bYR56Ks2N
B8gK2y2xu6P5nS2KI6+BblWHwH77fxN1SSeC/U1Y/vOWaQYu0U/hlcSxuyqzPU6r5j0zewVJhizB
lQlVQXVQlr65pq1Bzk75R44A0Bq8qYjzI5/6ozzU2Uy1PX/VSyDsmvLijv91RCYCy+24cSXlJYMi
UzmEzpzefDnEIKYApyJqni5dDVvGl+4oHkQFPVhsIjN0Snfg53XdPnuB0Wrvaq1eVVWUWgsQQEXr
kUggjSdoBtJsyOH5WarAu1BoDjVN5xGvDW37RRFZ1hWrOTkXVJteAPkvpuzWxu7KLdv6peLclBB2
YeQE1ffwdRDCq/DpIpYuGDou9k3NDhdDa/1CXF99rcUhKvR709KAtEVxNzzoRss7oAblGubq2Y8W
/oKplfv69qa6F3cTN2ITA0TddDmNkd1hf+YU/aJR141yifUC/gPfXEpHY80yTWKDgV+wYrD7ri2R
hGV1te+cnncYXgtV/Mqya3IqtIzvWeDOWtXvrMw0uKoyF1UF2+2u1rD5ra/lEJSGPSv+nktkEz0w
pHKcIHiA2jS7gtRg6Uqna+hPKhRTj8MkGMaixMGw9GkTon9k6MAQ/9TynYCAiv0XJ+vYrdDddqn7
lETg65qIOTFPryOblwH2p552PA83CuKbKb/H+Ct/yXy2Z8pZ1TNQN8Cmbws0yhqYQm1U/CYceU1m
weGZHV9U4FoZ5+1Par1wI8GjOTDW39WyGnvbAe3dTk0lwCKngWSB9WbiDvUXYXl3BBXrhKHqu7LW
cdYX0CwbFfkYTki2c71yKOKc/rcBEJOrn2M1x0gVZC60hbh25BNVIZafYXH6jNs7h6p2JnEHZaTD
dlnMB/ZAWV3+5t+PvhAw+45+pwaTYU1jkle/m+3YE3o6NSfOGYZccJcjhNeIOqr3cDAlXwxfDaoD
94peY9lyhey+UVUfDhhhsxY2dJC6q64RcMyJLNHsKttRI2b9nmVsYgHxrat7s+eSy5St5mX6rxgO
AhGyfYpUJNo5aIrcOe+Pnf20fB0+C5HzgDnPp/MR2s19R7yCIt9wkrUFzZR1HibOnKZMHjOdB3Xy
1cM08TDqeoY5786PLRwZiJztGHDddfjV9yAiPCI0LJDByiyRZDHBlnfsoE/t+V7UWbkVQeVC4DGR
/s0RcflpVm6K2HoBZcCUumcxhEzOWf5WBD6DPHoZip1HP1A0/rKWAySs7ZwJEWSVj0IN4e+LVlAa
KqIhjfi6LhZCYyJXlzIEJ2pKAQYHPI5JcN9Ac08Oe5BtK0tLWmRKmO24cxBNBLgDkYZwZ/Xpd6rI
DRtipFO2w6SQmyDWZKHzvifRhGhKK0/+bv6yP5I7Fpr1pqOqIH6N6x0t55F7LBPxWx0P9OCmyPQH
3dCEJGBb3m9Mq9l2kqsKT8TGUhQ+xs7kLcRyU7ng5L5CS+o5ryYZ0+MyEtSzDOld96JsigoK3jnR
YZZiIBDKlxr2qOUCyoxDnSIvV+qGEqfvlCJY8vST6S9CW+F+HL02kPp1t1VA9LdjDRy+L8Y2FeMu
Mu2ky867q7WYWC9JyUzXBzB/gyYeQQOLLLWnM+5ySlPkpuuAQVaTpIrMOT1DaOL8OkkP5BwsyAxa
8c1b+d7Uc5KvQMUPlFLtFr7PgdTup4LpdGWYbIFbM9jEBa+R9B6Sorwwv3epW+1JOCaixbj5GyI3
rN5CzsoJ227lXy5MrGCQQi4vq1cFkOCKjhDGc4NP+oidfcKDM5tGYh47CojUqf6QUFJdMEVyf1lk
q/V9T7gd5QjpPNKVDhnfmi1LprmrMfSHc7gTfKPnXLipsMbPJKJ1MURqpY+C3ZAcPqzhJ3jiqw6u
XHy94tOxCBiMnIbYoGZ2LzZ09v72yyn/qJvj1iz/kE01VSxmSFmJ4JFdJYgYswVPkayWOxEG/ZGT
x55RuFT9pzWCnpTefnVRxW+qiAEkTPptISkwSvY7X9r5f9p83XWUsxPMLZ3PhSzhfTpMFk/q+FWV
dQMqt4cLwrOSd0YXskhRiT1EDx7UNe2YQnSlwNj1MOLT6SfztEtptmiaOQF6x6GbpxTOPDZsk3+L
ZHHcFSTkRa4+cmCcgHjnG5PcpyyLZQiDUeZvzh7rfJipOYL67UMOHzHlfb6WRylmEhCP2pITRJvz
Wy0W3B8VxkmNZ2YFLxTmq3Se6dVNVnzxMsGnIjKZsPnQdKk3WPrl4P+7Ckr4aX26xyQSlWG+f7qZ
/lhHG0DDM0B+/86vFzRWBaD1drVVys5vZHb9n0k9tsw+o+veZQtfcnGCtltDxOxff370Q6uPZF+s
sNqnQqxz0i6rFXt7N6jBbp6zXU2YBMIRRj6yruguxwxpnWcW89GuujxWoQALteS0bLde7kSdBWmO
9EyhuDpxCfM0PtBOa9d1F2wscID20zDDQcSWBx4sqV5I03MeBbWW5OTo8xXTkgCaJhy6kn7AwPWR
71Glc8A1AwvzRk4NqKCKK9K0RoI6JpRVbQHV7ufQGxQm+ThH1SuJNmHC0IV0DMt/8QCz8Xu88iZ9
bpNXgWkYlNvfwPXu8yYdRXD4lO3I7U/DNQRCqb/u/4YILQd6Iu4YiTss0s9rizjr7vgFdJZp46rZ
Rr3dp4Rftq1ln96yC3Hy/dBdOEZyNvLM4Hub6JnE4U/Jac2ith0Sk0JPCiJ22xS/LMUmKW/fvprL
NY93ogmsuC+CYnc6LnEypPOKMSspkKrsR7/tnsD6WI+JTJJSKWMWI8muVkl2Y4bmMvJAL94ZqS7c
0Mm2U++gad+e1eU1H03O01FAwBC5N8tvn/v0N6f/CRSFFHiUk+z3Lo9rJf8RGxLznDZvWyJViJnz
xrOMaVH4eyg797Yhgy5DuoLBRtDM8lqdz/qWLilRRVpjo2MUzqeD17KDrhc0nc0vyXxcGIuDJbNP
zhR9qGS/AnCl3s8ok2f530aW1kzu/1zV6llaBYsWHL773KWI7es78tqZAaxGuDHfN43mFPk48S5j
B/UanJTlunWYR6FSqpHjnJe8SjXgYDs4UzsPbMCOcWVDf6ro8NmeBc8GiXjiRQKCleIlp/J+D8CF
ZDkk6Q3QcNTVXSn3EugWMXYlCrYnuQTui0UOmufD0RSqh1Qi8Gr6JQ8FUxbjC9IDFtUaFCM/pwtZ
jBukpeg57Qxki+Ecv+aregxY08rFOHfLpcNEKZGJubj6bW04bljNO09TVVM3nwNeMYJGYnCvxyXN
ak48ymYXkCMvqOoS7QXivTiNc3jOBqX1KqXfxhXjUBjyW3QP9HpwZTwb9FuSMhhZe8JAQ3ISdSaP
+GZbE4qY/0kO7FbsgAmtKWaIXS8gK0u0/c1HJHGjlDb6HaSD8T5EiFXzL8mQ2/+2iSLKjZv9UThd
lJPxH2LUcK3FlUBA1ttAVeQfq4P3WC7Id8NX7NVDSSR4I4Zmy4p+nMqRJW6eFbilYMUj5U+MNM9s
gVzJQxnvicEhpDo6QGeECyOHnnXVbniH4Z8mnnICnWZMULxIBQRz7dElGc5r1DZw6eexinSARMh2
/MNlMe+x/E9b1uqXxpigPQ9XLCBtJYJi7DSu647TzPq8yjrZGiuXoBRlmxsmr1Znj27oXza9eR0Q
kHBHwvm5B/+VG5Ox6EWtkD82maU+617VmtWwwYdXI8Jf3wRJCnTXusk9kCBWj2vQAnreKkUPR2jI
g1JMrUBEKorDmg0GmZSpPn/SsRqXn9kAskqAGRzBhIF2tyfn+ST7yFM4LHqQ8Vqh5WP7WljNG7jX
oibqMhq6K/ttzRBOB+iMMjjt9A/GX1ZkVy6tiZfxZRNzzsyGRHnRMK0ffoCjd2R0idk7ytqsJCIC
Q0ZzcDzQAB5FQy2diQg39v1lYENAiaCER1sSXMgNqiUsCDqnAvSN2bWb676BMGq80Sm9eYtW3KWc
iS05eIcMAMVVmHp8c2DQUtRiyDS+0PQYCgMp/HbBksYm/LbdRzg/2jUNJnuMdwTGrod8h7R0xOtG
8NuWhwvff5J9cfybImCXuRy92vFt2bg3W0VcwE9RSwHJgcBaRWlNtxHllm464zjXX2gZCqJEBtw5
rC3SxU6fTSplxlG8JWaq14pcyNwpWuZbgxXFWvTkCWjninhhSVfcUgoIL7Dy/0Zl1Jqn7jzpnUFx
OBx49NVgFsTnpbT2nSa+jY3Chhl+fuNLJoodmNp2dtrSmpcWrY7FeZ8ZEEGYGe/SnOA/nUl0l/Wk
qoCrU6IY+qmJnrpmEdW+ZhyWv0SMUSbIkuUq/J3TVSk2qIJpk1yeUL+2O+byIZl519okrxSE6SmF
R49MN5aUbODnas8vsH2/0JuEXYx+tFgEfIxjX/NS59i6YxYjPlQyQDjEKb1a7jNSHsdGT+6B6rqB
C6wN0fM5+IJgq1/aD7QrbnmOhLA11h5D9GV7f7dSOm2HtKMsUpYL3D/qB4qEXtvA2RDFVTM8wiea
y0vXySE0pTx8VnhajsVL6GZ3gH+x0KWdz0VRj22lLSL7+qXUdyhUDOX8hbc0wWhS6bwqZrAT/l2g
TISY9yTiX4aWWQMxX061jCsqSQes8s19bD0R/L6M3sUofVnB6Rhq/Gw8uMlvB7Ns71YPdVAqyALP
L/JqfJ1dko/b/lperBCz4dDzVgYFFKgrP3z4K5Z3W6pYuE5Ce9jDTnWEcn34mukg10JOQzrZXWql
Meh5zHns+GXdX7+GfkcsCAeHe36U6sikY2hNp0S5DKoDNUlph6sHnJbgTeH1f/V0xDlx0ABhdUDr
+olgakD/PiJ8rPiaeHi/ocZBv983/pBxPTzwWm2MbAlSEGUiMac1nTSJA2JFKQiaBAAh2EJH8Zpf
4RUFRkLkAS6v1av+kpz0h/h+7ATuTDitI4Seu3Pv6LBa6wSkl6RMPcnUJsJEwXeMyQPY1gzw4iMS
t+jHnV/iClUB9ruVPd4+ASlC18cUDJlE+zmebSp1uwuegXznqned2AHKQzE1d5ZJiG20yprJYZqU
1n4Ekws2vo19zb2qZCUj4cVSHKZn1RNkCPoPu5bHt+beTIvyVC8s1VhVlRS4b8Wr7l7q1OPlB8Lq
/Fwg/8fHaJkXsw0SJVMRt1ko7kBdqb/pEGTqFtzqMKL8mfSCVrUv77cU9/Mc/egZbSbA1ORuWHrM
nz5qHemEZMWNmFJwSsDJ4bPrup7G16N0LNwMiXO7WhmeoDzCJ76v0YB8Iwri4vidPK7bEsBuTLrP
bQyXC820XPnUiKe76joxJtmg4qO5xl2a1dhglo6NNhxqOwZgLRovXsDA63qA5l5bD2UEXFWMGP0l
LCMoOHSWCzgIIFCpFiI4QeQdQDra6yx82sVoWlvgSxyhEUhKGEeWxLfAyc95pGJUDsvsE5b0XrMo
v2CpR7IcFebg1W/qtEOrjvrOr7XHbLihjCTK1s1nVMkwdHY4Jz8FMYtyuPQsHoAUUoeMk9KVfgHI
BYk6D3yGD51jp8NMYvigVRAgAkKHi5O5/IZ4n7h8QCUzpcXbP+1gvqCDwuc1D4+lCuxEA0P6aiNK
LAbnP1hkNYSumYntJDXRC7Yu6RVp8Jw/XnHsMjC7HB0aaqGJommBpI/YbeILTBhhDSZyQJ3Yx2vl
4Dy+ofPBDr9w+3YAFdjbzlgfVOsgfW919IudmqF7i41iOmB8Wtrg57GseQN8VL+E3/6tuSYsf8Es
+qw7W2/TtYSfk9dOZcQp2ro4+MZk6JFU5+kG/wB9kLFQ4EBN/+j+5v6BOth40hmmIAFxc8luPOfn
DgIRWM+OQiksh/qozc7tGCGn488n4DCdmyDYYhI627OeSbgjkpPVgi0TZ7iOAQJVYp6RJ9Q4E+yS
mC6nENLWwXylMhyUUGyS5/LL8cSoS31QNi6WqEuUkzxkWrrUg5InJwVjfd2CLBkUCL7mZX25GQa+
l+wX+vgsymSzdX+kEQ7E65hGxJrcD3NDF2/75CvLowJe4CSfRJwv/6woAPyWA+dYiNVrOGQqJmvp
PBLGcP18L28z2IQBNjL3ItKTjfWW8Ws4rcIxu2bYG202K1KpVM4LPkBeHrgePN1p481V/Prn5l9Q
eI1onZGs1aYWWno51uEKHWpd2RpQXOWn4yP8/MSsdSnujhL2UNtgvuRNKVZ2B/t6b+reOSNaUWPp
kZ/y1dJ+tBclzE24mhZ4l48pEabh75Rj7mMTN19kVdntt/Q47UEZxWK9eRd3OF1w6aPF8XjcPkNs
FOry0Ew3M4WoDUFX8YdGUqWbu28XBG2ELAgfQunoPUhjSCkBz4xd/t46k6IvLbLqG1nos82rubft
nXawV04EZ4u9JQqD6INlxfgKZCwZTL6NRAJP7UBTQTEMhuizE9OOtxa5ZwVEBYgmCQuM/Q173L3o
IDfj7ShAhbidz8QiJ2rMmZ2PKTOU56IlAegeIDW5LLuwHMjVo2Hj/f0Z6d0hSluNc7tdb4zHwTVd
hv/dqEtmZgxI+t2CX0Yy07N3T7FrDiF4wvJjv/6BG4vSh2rrtfm9/n26Ws3jT4YBlOLDSUqETFLc
EldKZvQoRfO/jLAdgpaWx61mTtvnWeLIPJSWz7M7TDddVaXfo4RNkB5r/J0LR/yIMJPnsU/pkvvw
8aXbqViMEfCf/AopQpCixuRnyKVxnVdo43OGrVXaKzmUZq2YyUNUxOhaZCPGHpMH2eqgO07IrE/P
O1H/2csVEnsBNBpwJD4KQ2iIsVHaV0ld0/2gUgsyIuPGrln4+E6u7+qZ8bv42PQJ01rFvz41Qs2g
r4IcLbDjriPrJ7v21SFHeQmVjSqDwFUqGbA7nE0oKsjStSYHXuAC8p29e0Hyjyk+bqZXdOGxK6ia
U8lT4+J2d0adBMfjYO+/ToEj8xCy8Wya1ffBTAmQ2aYewEBml6r7eCJU+QDFfxiEhaVdbMLHTO6B
dD+n3ENh8+pWPxcBTE3jMn7lR0lhI1kgR6LhZJHRNfcK3QPBGR+UP7bWeI1ByLa9DtZ5BfPKuTB8
l/4sXnBX6bKzUyzbnM0lwcd+WVt5docbEQ5u1FB1E51WLBd+rdoNuz11DslT1Wcg4ArQXiHqMR2i
twr89ifxkTHjkKqKrymqPvjA0/CsIrdd6lG12KFKAOTmaz9M/Bed51rNDRiSBv1pPYj+Q0a9S5KI
HDrH8YvuTqzap8aQd0iCCuu+M6XyXPBhpnsZPQtyR934e5+o/cLvRuOhnKLs3PQM3w0mDNiM4wcG
yncMUQQZ2WHRD7vCfm9L37pBR3P4To6Wy64Q4/BVau+IACKxVMkuKQc9pYEH2QKQug4FE7JDweDF
D4XiZZuqWoYq/2ulbvA9L1Un/sb2iohezMPkcXTAx6zNLH4xCEPTj1+GA4qD3zH9le7UlglHbitx
pxaByrKmG0Jvt3IFoegnYX0rPJYOS9l+c5BHUIrPecWggo7MydEb9koWLkHHCDFjRWu8/qXSjFWn
uw9k3a8L/5tc8c7cJvBQRMHnFrb/KmZYuXWIbAEP+dw86l9JIv8Seb/26TPkv8bCDxXeiq8CnXzP
2OF2BTUUVE/ZKBxlY9Ys8n915l9tqjq0ye4QNspKWpe5H622yDpwZXkE1+kKA0HGd0IjNfoS7ifb
nTkXYUirC5PgHnsYP+iGAQbIeq8Pdn225ysqRJtJ44Edjp8S+Qi0MQDwl1qzhgNOPYwhOeGYkx8y
bQgQyYhayKvSWsE5SVRvHi3vR346aFrF75U5xMNWNFkolQsoVe8gcmjhpkruPujf9coDUwQq7IEO
e9i0r462RWNG94ndpttBQjRiLaiD6egmk8P8bRMepDhD8o1tu1LmnF2w9ZM3e3l7A5sjtU0JOzki
2/RvEYvcWVtaMTKRx8xhgNYqZ1AvffjiVwv089b06AZHrIpohd7LUXApygv9oDr+xgoq3VIzrUOu
zMWQTji4VAUUM9URb6P0qT20nf7gjgckDLcwUYiCQ3O+WQZmst1avueloS+T+F55GK5E1p9Egpmn
YfQZ59Cu1hm7ycvBVuzQoOvYzqnd4UO+m3a+2IUmo+g2HU6BLxbe0+Yr+AjxjdC/fg1MDquub1dw
7cGbnkZelkGyBh7lNKMEApAV5+e8csG5FsfgcM7JqJLJEO8TOWfsepMSUiM3f+WkaoW3yyBXhXBF
8OGR5iykcKD0d3K57j7svyg6TY4WnYfMQ9NHsVf5HoRdIKe+8mc9RwO3wbzisqJHbebqFiNJXtgQ
c2G6RVAUXT8+5S2l3zo6Ei+oSujwH4Mhs4Zsz1MrSyNpotEm9S7wRahQhug3MaT50ELL2Cc6qFNj
WsybuzAi7FF9tEHfBdyjhH9nuPSvCpX1kQO9kvocJBfSeFRcr9gNepufsNawJaYswhxWc1LICESR
E9C22kbcJmk2iLT0pEnIWROM+sOyYp8sKMH17I7UH/pSF9qMKa969xy+jNURoYGqriu8xHf6qQne
CVjxgkYFjBtQs37kFnvhsWopya0WBfhKDgKE914DEujk6dkwg+Az80KjAtpYE5LmCO6p1O0ewg3Y
3tcY/8LOrGR2vQKLgDLXj/1RtKUQoLkynvAIRzRxta6ESgvFwrFz8pTsZ2aHxVGgFpjR/OkkL3ZQ
mwuj+wH5K8oKn8Fq+gRMW0X5+d/zCmAkxJDindq5+thwPPXTazYZJ5RgDQ9cZdNvse22S1WIPCTx
1vmm58C3NPLsLPRazvZUTtQLvKzgWzG7dSsg0mRxojUGoL1OaM1hs4zQbvhobfGHhDnb3lNxWJPW
ZuDoeQvRJTLEYTEc2zPbjXyba+G3seUmr9T2SpocjdLv/G8nNmfI5FM9bFLJBZNX2nl4M0Q3avZ+
BZE4kpZMYjxMsQkHny4UKwCZxC8P0RMzed21VJmadMOOFxuEO29ApKo1VtzqisL6Fft3c4hmYuRV
eemjjporbj4tlwPQzMEMzTqVFeDyMpdjgToIYCVKT0WN+aWU1kAHbDavu1lhbxPYIi7CdpYAMU+8
Q0vo+Z2qId7yScfA8CDyE8k3/uSyedFx8oKWy4Wnr8qdPq0aMkYlxNeCctH7c6qb35cmpN1fGnyQ
xYcKoUxdIMD2755Gyojkep/LsMpawyUyLlsuzNUvuFwvXTQ6mc1CeJyFpdd0S2Jcvf2SR35TuW5y
rGAJXfFoiGKf2ZUr9y9hEAFoyMtscH/fyWmvaJl3Kcl5CCluXT4trS076Yx8vY1oEgtI4MCSUddo
EcQllTDGMordtO4fu+B5+kQdgh9FaFmhObj/2LdRVk7++xFN7GySICuPHB4/lf/GwcYt8qWQ63tK
faRIBKS7JH563kIVxXWuUmLSL59VVdHsuNKObPD/HNuUcD8McCMj0PDuWis00PdDEgWv58BKRyUD
8mpZzTP11WpL7VUm65WLfDMHzqRO0dh6pIWuUReA4K4faDyil94iMOcV4A9NYUC5nZfYnwE884fe
ZYTtYWDG77zhGKo+oD5rUfVuZ5/qrkWk/0+wryICSAsEUOQJjFi8081j5H44d16Sdpw4FdxBHD49
El2rtX6qA0/gIVzb7UUUWeU+yliHQ9CZzU9PPYlibAkyrCyE+aK5norgxx336lX717vd9951kPpG
j2BsG9+HD3W4UG061YmiO4GoT4VG29HmIGjAmoYRsYIYIgDLKTKYJc0dEaZAs2dGOlmUtcG9q8eH
UIaasumZAPHoU9wr5idKTVlt3UfznwZcvpzmYkGIAV8vyt+M3F8+jtPu7XtWk2VEfioIHI9IyH3a
4qERjJpjs1m0a9vElkkySPFUEablETdJgCGYVFjZVI6mCR6/rtEUIdqmNkoC2Vg31yxjX6+p1Qn5
cc0H5UJTtudOMmZRWzqLjlP+XvtkrKFoi1mrvBeBynGBj/3Gld1pKe+6P6immEpWzJrgf4MkpSSz
vjANBH0/YgL1PEiaL3ZpHQRKaSa9GD7FCFJsWRn4dW7y86LkG/CX5NljmLI4hCxjaLQ/FeTsOViw
gblW+sVU28mXZTSpzONfryNKVISgQMxjSog0HCkFIIbnQCQ5GyhooZ/8M5+oYz8i8I8uEalYzW+K
17w+JbLEgRk5ZT7SJu4pmE7YPGQsD2XfZS0XNLC75B3evY9GWACw4gVG8o8e52Fa1zwQl+1zZVqA
yzSA46X7dCHNMXj4MlBOyf4Sa7io5GoQhBFPttbjMGZrfbFdv07JdUXNutY5SXe999m743Qccb8I
ue9aPoyJOC8nbxejLad+Np7tqLxcAnpxyo7ehMTyte+WNHePPgjPKYjlu25KQnzO/rmtF9eTZPyx
MUzHPxDRW1sw6fPUpU0VJCPHVaoTKW4LApFSQ70qUcEFXbsfpJsQYKW4jdkRS/4BE14WGgA2UJDF
1X981MSWFlSJOy+tleHnsqYbdzhr1SI5sNEn6ZDgGudiBUX4heXxM32UH4uK6pc6ddJEYHO+9xU5
l+dAjkmGzKHD6JnZceMyqC4Gg5zVQNUk01zsi6FNzo9UzgMXvfXOafwngsOwlev3XZisnXFyYAFu
f/vhU2TI7gc4r3Pk3Ea0o1N25H99ej1y32a5NeHdz6f2IAGAQL3+wpkMg2866N9QDtAj5vKphPZg
V1yuT4BVK0I49Dtj1qNGqhFbttvC+Cv7+8Cf52ekUX5wv71wBaJsnU8fX9Jomaukqs07KmBNWuzF
dsZ8sOuBnvrjy2+q/FLxbg2Xjzu1hxvjCQZ+sVPK4xtY+hJmwVklypw+iWMD9GLjsRUsbg//KUHr
reD7d6I2lPsUytjSsxNrrUVJw5LVl5HFvbivKvCy5BCWjJz53BEkCerVrTNEwSaPGy1C18nVYDpZ
Nntb3Cqe2ToUpfyKG7LCOa6AQRDmMXESuqJFPAK37ZWvh0AuvNPw44JwVNQXXeXRyDX2rLzjh3KT
wCvaMBWpIW1lsfINh9ng2wHCbV97taw2IJoywmZtZ7Klub7oQZsYOj6ZT2uhi2ZGOYe7TqfsIHOp
mq8LPF5gnurRtOYPbiTINm3g4lMmFYECz1wQVuDsu3igx0mT7Ep53qfX6aZAQywgtlBgAhVgJ7kO
owlqjnguSztAOZLtc8obGKpQmccrP5O5eUvNN3csIeZxZswbgBTH026SzEJRIyDxZiKF0UHoz7iX
1t1jEFZjhzYu065ACd1DYkH3NpucjoEpNfeXJDldRpA7gnMDds8fdW1QGeDXSqiCTUuo61KbX0yU
RDcbXxCltk06UQqQ97za6T5FAd4Lhn06xuMhhl4nyDGPgAiGDCEYNaQsdTgXb0jUOUru1uzSDCIX
DGRYuAtAdNo4f+fRY1O78sKGguM692OPZjy+6LMSBppAd0hyWRpriC3CQ1RGv+yByn3BOHDiauxx
4KBQTuGG0lUYr+hc8ey+RJcWjGQ08h/+uyOWusYbkbxbZxOLOuJspf+pH9dOgH/Exgo4w9KijaEC
Uk/1GSXFBayBITOWaD/OTKvYV0EugD11XK88dneLMOq2erJYQtchScN9QeASwWAknEFoZSTPM7JH
d6RuTafe6HMqpPm9VwhP+mbY8pODA19NmTdAtgGs3SZzmnh+Skc20ij42mMuBrpinLewxzcHQ7Ru
6iTd9kbuCBMnziO2z/GbNdJ2FCR3bD3jQrOBQqMDFyQPhKW78nws2NtE5mETfNhE2uoW6hQutqkn
9srP/w7121c6n/bil/x98iUHIqJird5OUcwDoaX28Bivj6Uvp6Y/aEOgOZgc/ZSs2e5Rkp1I2dyN
fADh0o/1elRERQ6UMXs+rQsGRaiOPNmlPXnixC/xf+Ab7ERTTPYYuBB8eZPVIzLfS7trS8n1VkxI
aRJ0WJEPj3e7z7kZ/XgGviWMYg096U1a6L+C1g4glaII6oY3/aoSsVuFkg3gpEZW4cWPzSbbcx+B
ecXVJ2mynhz0Fii/zu4AaOltzwtzi1/Eb+YPIxsyLhAHIeDqsQlMqKh+59d/he13LW+OorQX+wB+
rV7hsDrZ1X69J8Jx5ndjujkyDn8szdg+1okOOnVS455BaZvM23utpqRhlBmOx0klFggVmpyYRT3i
Ufyp1hyGhrErwsAhLFEd+/7Bg87r7mAeiX/9jXwAwRnvKvxein+MF3uRNgpHZexpu2DjoLD9GOt+
Y24hdAF0lphttYdTvaHUQx0+4C+H/7L5gWMrRdyodJYBSW/IQSoJUQNsuBjgA2k2ujja7Re1bWRI
8YjRdA4OzVlIDJ/x/s+S+wbNzTHZBbx/JEOl+td07GYj9SkKiwDBhtU4y4nZKs2jh7hhOuj24Nd9
tBji+tnDTR0MtHMBLMw3dhsUuI0UNlIXXdjmfuKuocW6jdeI/HEC7PxM6fI5uTBawQOcuWwrIpeu
dlDy0JbhN/0exJNKSWajAuE7MkDdTJcDMkQMlNvBWB1CfyZiGKOcIjqlrXoccaVPgZsxT9cwGHWl
y/B6QdZviEXoKDjiPthmWFdvmSGVSec57pWkRjTgqWhWj/zrqYx7bqc610hBWFGmN/QGJgwSnlhz
Zr1w5CoFg6JBb52mctQwhyEKVpYUgo5yHlQUWuVIifE3ov87ABCivXqQEROpXCAcogr1WZgq44YJ
eVQ3Tj8Z/IfcJQhCbNuKAFyp5kHzfIlJbQFtPJ9dpFOLfCjZZ16G9bLc9akb1JKU5wanqKcpdHmP
608vz8qxOrdNhnmmjIWK2iitE18KTNAouqaNCzkfbWiXEFQtos08GqF3xPfnR7PiMmcA1RhbRBDA
L7+aG4MzK2dVfHZroql7ReBBT6HEhlQCv3ALuLlh1sc9Cj2gA1rbOs/+wAsQ4Upb4MQNFeacaWZ+
kRLqFr2MWQ19KXnetNEoZVAv924sdYqgv5ea+T0VRzBVOu+IDocYIZUxtty7cBR2OaJLPrr1mOmZ
Ds7P9/kp7biAxMv+VuGPNQhUIWVT/hShoIvN4XwxTAtqVok2esNFUJtzRcjfaXCxzRB5viXnbRgA
VkU4JgmsSxT3RgevdLJoyfEUc3fsKKnIg282btuBdnORYxHmlRNj9NOVOmzNZcTcwjxUitInNo5l
OoUDtA0NYlxj1j6E3d+xhdhVumd/H8JBD741fEoiAHlSr1F2faxdQVW6KYq+65LE8mG8pygsuNiA
D64BppsoDOavadpMSEme0L5UFrc0Amp8JQva2g4Ln8kh7Vt+sxuV8zkGQLOp7Us9bWV2Fvr4DPUV
vpPlNEh6vMSUf5RY3Z+O50AYKPaSWf78ynqkug+5zzTkAOnzswzeuxuU5GYyeiw7sIURmbqGVsL3
zSfYBjQ+ytdvCaSRbKTlYZ2dTeXg0wcIhvvWrJQbQMpoFQNvQCIS2cwxj9oj6E61xiAzpR7tamXA
9O/k2qO1Ja5eSMRZeKCziaJwdp+pkOK1i7ar14MTNrNN8ZGTZp3s4cX5gqdFX9RQohNOo3qVupVE
RuEc20PutnOXmp3ReWmOAi6tfs/zykqom47UT7b5T7PGdHPGy24N3LaMyPpHgRJxPeBqvVwnH0Dt
0UZrqGzlrWs5I738SdQ+ADeCnZ4V/YfQH+4AF7+VfgBOAducFsq8ARxbI1/U8uRePNtcGeY1qxYG
8dcf+ZxaOKq+9wLun/UsY+dWt3g1UtMa/udfm5Als6ucAi7gYVxnhPBVoHtqSrg4fuA0Io3hsoWI
tDS5Nz0JKzCTLkZperDf5lDGhCZdZOQ7PIkoYtiIYs9YkdHj2my/kAsHPTL8eRtMQFE916LruDp3
MlK4NwPDOMUPr1cCliysPLEOS9Gx6887kNSIenHEMkIVEINN72chv1VHjZ2yV0FXdxef0GzgtYtL
EclhUClsCMxY7JS8oCSz+ADXVpsj3avwG00PaxqGe7mshJ+JnpA8iiShGI4JfWHswnlzcf2UaunJ
8jkED6KNPQVlu22UTQsyXnPF/aGCSTl6nl0gut8eZhx7NHvbilJZrmzWuWPDPwLdBIh3g4DH3gTg
rRXNC8elpUWhUxf3Zz0T0TP4UETi4ygiSRo2+P8IJ5s2GyHM93J22XBwgPf7l4nPgT9cwgVdeItR
TXUYaStlOySRLfP2lmtHtoJN6agDDWaTv1tj0yO7ZzAnTY3wGdwr/W5DVlrhDY4cQtE65oL6HpX0
OCunnK1+PFnI4uSfNk9JEsyizgemOUk3j+q1k3ODdzsyzzgZHEwR+Yi9lxHj0+m7oUI86CvAbaOU
r0Eflx8twXjfu3tY0R+6ZANA3NfbNppOyJz8BE54qm1Fepb3oTWbCqqc9NJ5ptRz55m+tr2aNuSB
hp/OydOWg9H6pfmBiFCo6BUumxs6IH1dC061s3FlpPdSIecLNuz+wwb/3PA+BufxDp+yc2USC5sF
dxg4aoX1GDn4pdSnVzYOQ66Ml3q3fFTJjvDLzIMMq2WqmnxAJUNI6MqdQTgsSHyxeFfz6FRXWnci
MHisOgdi+Kr530MKsF9/Jm0NVb3bNUhS2HJo93u4Tmml04RTfzLOj0LMwkqotDhYLJzjb4qmSxMj
jmmNYxLb4d8xzMBfyJUu3CK0AtzBPkuz/HfhAzx/+OgIoAbUQiUsqe+T93ynC9JLa61ghkREdshC
BPwznpL0Yb54Uw3JV0O10x/vK7U2JFUH1Jsx86QET1/1Ihu8DBXlV51Uz2IGd6nrInSYsNDONFUQ
F2a8VTOTnbV70iMGix5Z5ZkpveYmtp9lSt2Y96sFhDgEh06Gm18yfm3Qd3LsQjh5mCoiCqMAe2Dk
j9+ScD5kY3GX0Zw2LzcW8qYgNHWuzUJ+xWbUPL6/JpdMUR1zR6YMZuD6gJ+cgUFmrR1xFKlOvwwF
8BEQXaowKjSeKH33X2OU4JHLsR+NvxGVHdaLabmOWxAemePvcdya8+kukt9g+B5FGo08M7D91WkA
nYdFLuxOjfugAGW8mzHmnfaZnmtQNAiVYBrHGcgMf5s3kt1GswTpdq0Ro0of8H9X4evTi5tRK/A3
9l91fGrJhp4VWB6C2YeYDwL4QW5Xe6J4+6qZ5mKFIsNYwHRlTChot8+TVBVFQ8GOnI1uFk2AY4He
IMGMfpLS4tFAufhmQ0q0U0gFi7tuEng7RBkMeTpYrEO7mxohg0D2+6zuflUICB+jJKzR9GqGIzae
3k6t3cL7I79lhGY7enjlMcAc5oEUhnMMqca+zbxlzsV3ZnrXNEG1QNCd//O7SENLng1SlRgGGas7
N0ULe767STG70gJB2CUGY54dcDLkxfHZYrrYqRvE6QZdglH1EpswmTQTO7YD6kNus3qMjb4AIY8W
20wFtLmZ4lLrlo/Vwekdhi02OmVO7IkWGA8nJdS2ytG2iJr/S5SXbj4WUaQdPaf2eDB6nBiwxmFj
hnQp4qUvExL7vPdgCj1AMP9xHbKesgZgqgmbT91tRVsezTfHPGHdawnanAxuLtiztdRtyLyCflOy
KKWQ3sI+W3pIPOYGLLQlSijgNowpflaKuY8+Rk+cCt1DgHaqeOZdIcarwrh+r0pbP4OMac97YdCh
4p1CV9GFplqyslJYIxxZjo1bGmH/q8RzuZIYIyP4a/QOXCrznux5UAPcdFAAv8jkiedx0+LIk1Zc
U90J58Iu8BXZK2D1R3K5Gh91A1igrHb5u5niWS3dEjfGPj/WzB+5pJj6t1c5ud07D0DSaexTkmfn
r09AaBpNtMCoYHyY/4ebDXmjlV1RRTz+01r4hiaI+N/mgSCHYylrkRhLgkbdrUzzybxo6YB/njiU
K+vfUDhsoVeeHThjv7Jmj0S8ycyD7hJcsngx9lXTbJb33nvmmRDMCx60ye6Qka9jAQFne8H9nEh5
tJkbvxdaT7vLChAMUzEA3g5KsgALitNRGKQQw0BbJSLifLA2z4j0LK0jgxXWxj29vI9hldGlvxYR
huTQXaklEDG+2WrEwu3NurRl7sx2t2IboN+qawm33Zo5dNKKSsXt0xiv2VycujU4C3gWUOVQWWNk
EkdXztwuQeMGsNyx2TaojnC083RK9Q3FK2wHRyk9QpCCnJj5Y40R59eajoqMWlepr6OCdKVWUuJR
fVs7BtrAjkO89kdoP0inc+3NxLylm+snmv69qAX5sV7mnBj0eVgTjTd1Wg1Kym/skPEDW4ltxV6r
GpBbOuinkfNHePKNl1zJ9VViAbX6UmvWh+xdy3Ti2EMfPFBWw3rZT5JVihcNdNCZhsF1Ob181jmk
w14WEOWjjZa73s0+qd2nWRJHxH1vGHn+ap+RydEl1iyoE2wwyFDjkyFzVIQNcCDdnxaR58FLOT7u
Ay8o13AZazrXi8lF3/T4oorwB7wS5sE0UQZJfs03ikg94RLDpFD/Vi4ttrhwZZy9ft76Rgz3p51y
piYsoB6zLvH0Lms+hNBKg+dWJwq79EyhZqbl5fKYS+DoVzr7iE7DHID/FPdPdRx02Cmkye3+I9ev
kezbAYyjw94dED3foSNSqquOlQLJ/jOzReVF7DuctLDsKKwuV1Z890LmBeSc+l5ejClBQ59YeSJ/
l8o1buEJGohFORlIPATUuUe4EMBt+zU2eLhUER4OQBEBjG6cJWAV3qxnFcwEMMwdYdWIrWFDQ8k0
Qg9zIVpIEV54+YbuVBt1p+nNrQ0SD+wCoBuFgErWd2MBm+PT+09q0QyDCRt6krdlePcEo/tos3iV
lYiP2P8X+nvJhyvlHp7oRXSRDZjriX5jw2RKEJ2xg3NfhxVoEBgTXsuNQmx0T8pQOQaT8HR+QN3G
DONRySw+2G8HDqNk11RYmiUCV8e/6iwrTgBauQMSWMm/tLYLx02i2K+DLrGeUMc2UE5sWG9Wl8ju
WjalMhzFpxfKv7gBpzPolh7zIzQyWWMkFGk4RluKQGgufkHPuUkJGPMl4I1uKdc7fCTIq8m3eEDC
Fnd2mHcS4nzwL9iaA/ske4N/gTqnXoAJ0mxNsmROn4ko8Vh9U10U0lXjjjtfVhLqVHb31bvzIhiW
gqIJrz9rAtyd+BIgiKrfMgjMVvnI6xEy7mG1CFND8pN37j9w9BtoNc84EdlVNrRBLaEwvSbFk4dQ
9SFujblHcjCAmq88TpMtyQu4BSZgumxGLR/T3DRMKkaTvgKkScliewUNqOE47ZY3IBcWRLH+zurS
qQe0qUNZmZqFxc5RWo3EC6cU/OHObT1Hut0ub9WagJs82Hq9MPXLZmajaDXlWQjM47Sty1vn/zNW
PB8qBagJ7KLWRUDdVHM8YLyVbJDI3KFBqppGZOAds7imlrYVXrn3or64U7rutqjz0PS0o/gj2G0/
ogOiMEcbsvL52PmWgv1O8iW1G9yGexMe5sv5SHJIeFpo9EHSNL+lgNA8BE/oyHQ0E9/yVrgtNrL4
qC6BqZdqFqobxAs4oF//jUsTnJasCfvb6wJd9r2eYxqpvA6TlvnoDTkv4tMIg/TspLI64KlFQqgN
i1wJqvhSioo8DPcer0GTtB3ABeXO7yjn0BqLAimDqvwwcDWbrLbGON8uPuVZnlqC1wxprll1k4R7
36y7yXqSBxXFhY7LzW3QuxdgaLjRYLMTGFJvH46sU22v/cUm0T5HLyCYLVHin9F+tmpAnce4OSOU
T8EHpes8mfQ2wo7fcn0723sa2ot7BCj45kE1uh7fWzK3GRSR11bimP+YC/GfR5dSKUIglrkl6jK/
G5fdVVo+VVlFi124myFZjvBR6UnmQWQK3xaJfjEqVUNwanHXuN2zwQgX5vK5m+aehbWC1zoEjjSY
YCCQDHrm0/ju1KrS+WHAjD/8+mbg5F0oGIU+a+uRsP5k1OOan3gWEmNA59XYuS9dzGnZmxCysJaE
LCXWpd4zNnD9JSAWcZD+qsfwdwVxR6UFWgtspnPxs9FokllOjghTiiuqmPsZQmsnbT76w2MSwmrt
+U1y3DQ2APLQZ2D4QDER/I3m9KgFC9TUwazx633TXUgsrdm+ToKUMDxbWCtXP6FvT8yhn6b+t2dG
UnsTk/LJxNi612/QjMIX11h44nTmboXq3Qbk1g1hGURQ52GlOR9yJVXsKLFDujcbZOfS6NoeOqJy
EzRmlKWvkw9Z566m5muhXbTpzgq1UO9Q7iHqHiwCDgnRq+nJmnuHho5UPvDo5ew6Wzc1KW1TrwkZ
X6/pfact/WcvcFZ6C15awvqGU77KmiMkq4PbGK3iDkLOpCnjLhAtjvDU2hUynZk+s6k6m8MC4O2q
U4uQPcKWT7tYO5kA+mRwuI92aEgWIFDIKsrwrlHVmHtej3dMkw0IqXW7EHnFeenlc6gbojUDYI7a
P92kmlT8xgHFBONRh7xJPAwhDj+c4Kj4P8BA+dclMhjivevrrN8rn4miQ1Uzd80DACfkmakPfcLL
hdbjCpHTZif+2WVcukaHzNr+s0fBJmVvCnwRQvl42nR+wUyfFy8v01zJmpUWn6QWW6udxDGaxej5
0clH+mEen5wBwLf6NfBrOeM3Tf4HVeRB/sHqU84X2QKodU5wbrYYCPNH5vUnuA4Q6Td3wwN/RujK
OohFFMrSM3njSj/f3a7Mk/LiCT/mcvQ2kmivMF1H+2mxwnyPrVSgzpHNaOJHQq9jZnJuTDlUgSqp
oFMNqmdKjXqQNTa1n9T94tfO5hH2B2IaQnDt5JxCpwXN0UkAUxmNJZD9ClXzykMovZPPQVOUO9WR
7ZbOnfB9XOrQALtPENbD5mh/a8DJz30LF7cOsG69OR4OnbxqPPMZicAvtTjv0Iu7Y60rc2gPu7UC
nVqqy5xlRZegFKoQMqZ8hS6UDj+MZCSoij6u6WzI1EtpR22QNkomRdt89z5H64ICLnb03FnjDzy6
uXNriyjZtHTkBo1uXvvCuUiv5YiSaDpYIPFfduUdE/vVYuCBD6fEumgWGmrJhnDE3dkPnEYg+No+
L37RUHp6126qgu4vlDa1NNT4ntwhzZKvbjRFGGRafxukZfmKCOemU3IXDpXrA6A6ierSCM+7Z3/m
hnsPFXhA93FRCD/7BNvdeMLJQ6cBrDQ2cPKISb+8TviRW2UjYsbEbmFtqUrDPhBFXNiDUwDuJ1Y4
t4JwHHcGDmCiO8CtHuKNV5zXeMIrWqkTy6sd7pACdze2jlTqrnip9eMkUNDGCsjQ87N42MNcOHZV
ouxRk36vQ6oaGMOlii9CDvwqC4rNY1GU1Dept7cd/ibDnjAs8eJaSoiVaVuuXi6BI6zSlhDtq0r5
dqbTfq2SiBi7jFI70SGazDAz28acQHqbHaQz+V3X6ADNSDGLEq3tYz+fQhEDXc9R2D+6JluWSo0D
mHAkOHnCTRuo0R37K5oaHjbIB3k4rxm4iSKdpDMS1mlbtAbABrNmBB8iRNyOMyuwxHyRwVcjcOUd
gtMkzOc9J0zUD1NEruLcwO4Hhq43+HQOmM4XZ74XOnWs9xPzvxmoeFpmNOb1D6zF52CNzlnmsLpu
sO1B0k0o+pBT8VXI3A7HvEp/9Rm9EG6hjtA1Xg2TkSwzYpKpANpRsg9cEPGhndvrdro50Q2wzkLP
LVWUml9hyQ+mwwPyeEWACiAGSuXF2fr0aUSnRxwQ3dBZIlnCHQVQvlIQiefJG3QNDBE3OruPnubU
ECOPHvjiuclbSIkA7CJ6gAE4i7aHg0knWkoPT+PZcdclFBZ1PltBBRlixBdKpy31eIDusJC8+boX
9DiY4zkb+3YeWe/WEt0f7lPsrHXOHtPZ/A8kith9uRihMvVjb5yqYROA0j/481Gfai09s79DSLHJ
R/JUl+6crwwPfRSFKKTHb6jpOmWIgI9a6wCuU84s78l9JsFQI5U+6Ef2qkiIG5kN/OUIq2Xz3LJX
LXEG8NP9UY52iOtS9Exi+s0Af0eP5/dap8SRa0viW97caaZBeh5snAe6i9vA+pc2RoNJKdHvJdbv
J4PjJNTf6cY7yahf6r+E34Ajhoj6rTrm8aJRtW2ex9TY8Zrr+12Sqqh2edUuih4HYFp7miIN3LLj
HKchrscw/pQVRRHpgR6cnmnTsY3TsWAdij3f4SZM4dMYI3k0qU8gguaDT4i2LTQi+4joJjDme1fg
Qi2Chpy5/SMJS4GpPUReKT67Ur2Po/jtP3wC85dxVIQs9bLaI+uC9lJwOHtcHiG6fqjmJ2PTVmfm
77/aOPKyb7qH8FmMMS2V7TFH2g/baLNQmgkC8DZ5sVeHDgjceWZlKLCUja5yXuLqtJStlVrd8QAO
r4GsHPD18y/xNvYCgmOX7ZPLFs2jsQLF17v9kuwIzYHfajXarNlOKo04fthYyBNYXxfwkDGXRlup
TF48NjmH5TiW5rHz0/ZnYe6mk9aeKMM/Xt0p3Vqh9vcKxBfaDFDDuzB5E7VI9d8AszPlX8IOREaG
RbbMZ/PEBey7zAfjBeSAPLl9xOmMoNmmQdDfIsuV/sDmlMsFRNBLFzDAoOFmgA65aus10RWtHcQW
dt9kkO9o3dQWtyzcBkG8p8omqI8h2JoqMB94J3TeV5TuyIM0vsfyClbZLSdlwFGAu6knEhC0Mby/
37QUfXOP2BZOvSGlpRg4SinTlxSvJWOplHARj6lsKczIgYfIm1sFENCgBK6osrnm+DswNK2esTFj
y7kM50R8KSmh+M1RH5KUZF9ETNtNks8b4D59VgndJIeg1fek3DKBuDh9Bkt4Z72fttIIKyIgpjU7
ykkTEZjmKIKXhA2YtzBN7U7UatUxB28fDce3GnU6CsGHehmTLNqWmOEdpTAGpwXyu6U4a5Ixhb/v
5Z6vAqtZqmx1VdtFo0tAhu7PLFyoEURKBdi22XWtmADN2rNYqQTcsby/A3ajTwTr5XcTW0hCkcOd
mlDWDhaSDxMHsaneC0Zjfo0uToedC1t9JZUc/aGakHjjJLx1Q0x8V+M1goqQTNyPiUA4D7Kui36C
XjKKEZhTB648UQbbNVAxswAAj7cpjnk42QuCK1r7acNGdwCOJ5ToBN5mlw6+2kTXsod4BfP9PM/X
t0Fkn8tVrN5r0ygrOS4pZfkQddT3NXV8Ap/f5vhCt9nwKAQEqRdCaGikoqfath2Gt5J1d3kdJ3Az
SgDG3g89f7OHD3xoRF2YoNckpPtSA36OEHaGI53rV4bwJfrHIOG0cWnigLgKKVMHMAEaFaelFY4J
+RMb0umDR9zMFGgxmQ4QWtyISrt5BOM7qS2ZefM27b7TDVg/lSNNcC4b/EyfW+JqGAicpUXFsMII
Yavuh7eSeJP2ccy5m+nT3aK4LX2kEw8RA5uwPbrcsWe/joTtmf7slVrr6pADv07S0frqFOzyy66P
+fh/GJlSnqm1QkMV/6cN/tYv0a2+8bmslyNG1l1UfEYIGgi1KF5C7aDgXYLQiMdviB6Y6VzJ3a0Q
w7pKgUwIslIGTusmWY6L4/91AtSORNCLMhyQurkt0uYABw+3MNUWygtpTexaqLWYC5iHrHEmQcXs
+mNi/I+rHRUTh0uQ2iCTjQjvfuqMhn8t+danhYuBGMct1caPrqwPNsgyv1pKncE9Pc4yLAi/fhdz
9RLGb7EmRZ66Ulgut4SXch9rot+Hu6jHb62xMzyNv/CdxBPBUVs3fIF0x7UNIGJ2/eOVT+0z3WT2
9wFAQTtwW1SFwWN1+ubtsExuUTIqg7x/ZnTC+yk8t5tIvr7B8MbVOSt4INr1mRREMhCvNrUPwR7/
RVwTxVNG7y+YkkJaEUCURLUFwGpmkQS3Btj4OR4q9yy4yvTqxTAjkx127roZSVpXy0kw8CNNP5GG
pHEDltkvslPNl/Zd+5MIpApvkPD1BFmSP/XeNMYFG+CvvdLp9yXRZz9gSghW0KnDaDcwWBZ/jwSd
dRvTYZDX0bn+ddXEhlmoAWR5BNlw5DEAfrNbP3oQyDTGIq1aipLHSMxGjcOXeVJlZ0y46yGd81au
gUB9uujedjw8JvLuC+Ey+On9YijNcQ5d+nABnRtaka+vIzoJMDMqdSCvKkU+PKXe+Ccdy97tHpP7
MNdD2y5ZlYad7BoRGF05V7nTpPpAYrw1c5+Ns6oQaD4KPr7Wptg2i+s01v+doRrpifpkimdGVZsH
zGzqQh5BjZV1HgjL/4Xs5biU4L5O2GA0l7LYbYnOPWdebu1QnaJOClr0ZcEZCJ/BYXWcJmxRHs4M
3L6rnIEKcXPE1QpBiBmiluC2KoIPllbAs5Kni5d8+7PyVRSgv2IWb7eGvHTrneaKVGGXzfCXvg6Z
IWTnVJEWg8+sWt5z1Tn1v377fVsrjPU5a2RqRSKX7a0JlNHP6Itipq3XypMTb11x3DAIlgD2N8BJ
m9+vU+d7ZCJog3IK2SINF1y1FVHHJplRV8oDTOvGlFj9FtNrtUykpZIyphyEAaNpilTKTQjKdt1x
AfPhDdvW+nqMtr1adnn5NoH4FTY2rG9z5Oh8UVAzXreyhhWJ5eY+0mTo4tzoL/xYPWhaacL9oTLc
/ixzo2AFlh5jPQl3rxcwFrUtB17JRv7rVJanBTOrFogZ+3ZUxwvC3buFbVEohkIkPWOZrq1Q523V
HmMVf//S/VhtWSdh/HcLHwJ6mc3AGxK4WqdLohqmRlyL33w629BBXSdCqLwXDJmbek5knfV0jarT
unc166lDn8yTcnV7Kv7J1ssOYQwtwWJJ5U3EoRmSRgInblYsTM//425k7QAtj2D2dq4JyJUxcTO0
q2nY24/WOZHH5TioJfHwVWYbawsB4hxYrUyXM5t8I1qeoVHpl8nKbcpG04r+eB4bL2lyfuanPW8j
5L3wQmWS7ngaVZMLlsnTFtNwVL3gGzMKobCQALyVpdkkN+OApEuu51luN81aB6bNLBhrL8DIYNMd
GJoWZnr6QhucUk3Pc6zTAPXuBPXK/1/b49oz8WNkGDXKxqZkOe4lCCMxDdKiOX4ojVdl7RSpFAVh
LAokfFF09rDG2WGStVvjsytmmbIpIxk0uFPrpTRWGjJW1HVG0UH5h5JBU/QVKTMsaC+Mu9bF1JMr
it1sJoj3z+SMbPuamYsYMLc/NO9KgRk0aV5qufvIP0EMdak8lq/PwKND68JqhYY+m8qC17zBJiR5
tEM/pwXrIf24x5kvsAZ19EqRrpRByoXOjFPA+4HH3PFYj1+eFebppsa/wJSiL2k7+MmszfKlB8h5
vm9JwTGpzWB6S9ivbSVI/31/DCbnKsSzivZGpHr1/l+jL6sM0YSNfKnhpExKKW6J/StchzLvT+/u
ogOZx2puYf69dZxJcefzNuHDs4nol4WjyqG65R4oiaEe6/vS6TKDnFlcZlLpN8rITpEOhE8vhK4j
Nr+7vnIbu62HrgLbJnkC0XewyuB4z4yiI6ZLeoNfF2tQBeVt6Ux+5QPABa3HFSVihZFZP9rL1xVq
w07ak8I0Vrk04AtEZr7sfOisEZGbWR/zzs6XiyILw4tFCswAkfVmtzoEe8yl2Pkuc0VIa4OouN5F
P9QcoHvbAcd+6P0mMGf/LeRSV/omK63VU9rnEh+UkGzVUIPK+sXAhgxhCiJaAbkhnG5AqyXMzWDA
xMzJg2dJ3G2Pyi/2Pjll7p5toh51fIr/UnUrFLkNk1Czs+GXzbpMT2I9e8b6igPY4SWRdODc9yC2
IM7ZEm2C9WhfPpjvrcfQOhVeExpa+mm64uu21y9DScplLPhLUGZV/sIyXwhL4Xe0ZfXFWGgCgtHm
wen4xFnizz2Bikun5jZfh2+JCd4OeaXLqNHQ2Y+Yf+wDFvgXQz/UBj4eSYmnZZ4i5HQ50hpcj0bH
vZTHA62GDc0a6UJ5Jbo94FYWvRBy+4vPaSXLwZgrRrGpQdKINToqJPCiPNvjnI1u69cgE9RGtbWO
qFEZcovNeyh7/sxkW/E2m3ErzDK51E7wFwcaNkMl+F7cw5PSg2TuMDHQ0SZb7pWDypZ9znvo2ZxV
IDCB+KA0Tzn7hhOswNKBEkeSJ8qHDOxbkocn96N5GUb4vtdeuH+sf7z4GOtWtms+kUI/I2gx9IjY
HFFE4AAq/40wP9URRoVlPqLJMBbI7L97HVn1eAKvhUKf5bneU+vK/kERNOEiuk3FAs8YOCa0PRHb
NJLJ1rZDrHyFnGVAm4+HIKIQASdccly6KUeH6KvtF0EnGp8EJ5ZfHERXx+m8mClF6Eg/n79AIG7H
sIvlVCnF4rvKQnIBI0bmRLb9SnrnStIBxd/zkSGoCvzhGPN89+FbHMs+dgtVpfoCTrqY/s8o0KEm
j8//lSNGJsix05dDran/ciz1a9E/11Bznp28lcL0dNXGY+cw+Q6ciHDI4SFWEZdGHFPqbwoYajpu
MFFOxt1rnlpwmjMSc8IUmpUq+HjZ1YUuhlaqqenIz90S83B7Gg8L+rI1rytqv4m0YekQVyLfWt+O
+a271Uq6ufrZwAMeXVhnTxiBTN3JzzA3YT20l5PwCgduGcO/h7rQI8OUUr3j+BT8E9hFQNRLrh8E
Kbv0bc+TuPg4AEoqQQRSJxzmSbQHPzioOUeiSbTPSOPNJwOMm/1vyxBtb4sBplTs8u4M2Z3ZD6RJ
q7V0TUg5ehsziIKFdW9JCAsRN+REdkczH9zM8N4iICROk+qmMNZTXcpq36x9+yilnA++Hfxf6v17
kpn1n7h5OD/P12S7l0N1R5ERuub5ohoM1GcQnR9M74JPEnuUsCxcYK0afiIaUp8aTHIltSvIVTQz
W/WMyRO27pbHYagXj6CKMA1gVnoLT/XSpo8Szb1H6nf0FLECAESqTg7QB8T3dVCvTruxmkgogFCo
sSE5wqn25cAvLGfUX/XTd5Mwjm2cfftaBSLsCw9o6T7h9wXH+CEakjxT2QzTgNWUzzxJvNImmw8Y
MEiYQGajV3dRUJ3BWhElKMSDrm0DJN0rd48FrQKUsPyUGegDJYdHiVe6GCOYa7NQSas1CYH7bqeY
7YqJB+ApH5G4XWM3k0ypB4FopP05DPeISrASgMlLvNRKiSt82W24Kdg83hZsZaGwDGzeLCZKTA8L
7I5pSWJZxWsv0bcHhFDFZcQWaNxWrxIZpLRXkFzkrzbGccP2+2Ti8/H0EBjcj1H6BYqmCuZrtyx6
4p7GSgV1SqmtixoN0MT0D1e8zu6GXzjxtyl900e6/HjwDZsNV6BB6igd7j1VjAqS2Gcyi0pEf8RG
F57tgMXz498MHK6qO5nnQQ4zdai80bEzinEQedtiGOGG0IvzLoRXPVfPTxk1OYZ+uZB9rgWuSZIS
4ZT1L2+fZvWC2eBZ7NgodMXfe8P1ZAUryHCOdscTWAsfUdkseIF9nCFLlbP0AgCH+VDGF4D4MCR1
9GzMxF213UsHnx5n7G+B7X5Ufi/x32jyyR6Hsu1zVKOA7jETORcUsW+2h+dkyGkGmCyVP8+9g1V1
QvsPFiY0lFBTG8mljr4F2JGAdDQT7/2fTCWCU7gq2ek3uLFppTQC6CbSDFSpKTs0+S3lW8S2/jVf
Rq37WjB7a2e1QyFYDQ8ik9JblMiWick0arQsrnMw+v9lPq2Hu619aH5jRKktWwyHHHPWLNUi8H+F
BnEVNEflQtudy3/RGV7pD42JvEd4OENlIqL2+3Oc8RSx+3XOIqavdt4C24wjomeYaMeLV+1wlV0Z
f9mgsNz6TY+nPPXf7pmjVehcsu0PZNoo7i4ZOdW3Z0Pa5YfPB7YAkV6FoMMz6gXysdYB8+8uZ6H9
hM0Tfk7nvtHYZsz39rLHqIeN1utALGEVi3kulpy97Q6NyMpg+SaJELdd+83xr97FduWyTH95qobf
JQqmz8LblVeYpT1MzAOa+4+91fQzHxKyT9itVAibGh2NTShEkTpF/8jsYCMmKaFz0wRQ+428jFtK
TqZUlY8YCDw9sCvGkOLTqMkdjaiR8D/XNECwIhoeRR8Ifbt+c5RRaytzjATt2lxQNCgMwBF6AQ9k
XILIrfycU7FGaeMiJ97ihbQzFupXMt+qUuQ1wBAB9JkasJobgJE9VT/uhZwfK56OGkCx451u6gX6
P28Y4pFoYmHMg2eJW8rSeqEjh2NSs3OB9xkKX8nvZwnyJ1X9o0s3VZMrQDjazWSyOwMXTnIItQAP
0yAfsaz/r2LWyXrdB6J+T4nPPqZMZga48zJ8jsTGZPCvhFEyA1hOw+GGnDrXB6ldj1t7ni/WPCNO
RDVyPFJzeybHwL3tcTzdrhuushny2QDTb5zzQ7Ghf2N3ba/HrB2BWRVpCcxfRrA26JkzpBS07g5n
YYQiUiIHZOO8TQ1ZVfDcBIfaBNyX25Jm1kJcVR6/ad4CyM7p/Qdol88v3PQyGP+35ROBNjPdimDe
ku7e4qZJe65hJl1DEsylKV4t9FqM1+ml/IfoVKUmSK+g3JoYTwgcE9lpmojk1iI3obgHSQ8/dLGh
evCYp+8mrHs4PbmlosWHxJaBR84B+QFh7YfBG8+LV0u8wq2aMimvwfN5+lOFn5NjoB1av759mpqy
/DnCOL4RwkSJ6at7ETUw0/pth0DxV7uxVxLRvgVY2yvTK3DZTPhczbbzJzxEyotbjg21/MtGxySH
RsaeV74WSCp/Dei/dKfVtsqcYGmlKPpHZAjyUThQMjHqEmGUowbkgKIKFWFy703kwcnEd8eBlee1
qgZCeoZnRhHym0Hd7q057bvCzEEmbXodD4ORkPTfatmjpLqynLTBzjMc/zSTN/RaRP4y5sS1IQAw
bThuHbXJgpsefNVRC7NUh/ot/k/chrN0sLvI/RYId2Z6++ZfFs3qtlFagIXr0106wlpPTEg1U77r
CTutk7ttpMqA+eEuBElMCByE94zICYNIQvMgyJhja4PT6AeBJbayVCzpLv6zou2wbc6sOR2VbqkS
jmAElSd9NMzC1FbapogvWWSMELU8bYHuAnTaVSLe7TspBTjKgmdkqKrFueBJS3/22H/fjcrVaTdl
bm834uhRiVSjgSeqLcPOoQw8y6sV9zvu3H0PrOAOLxWuCx9nTUEiULJqKURDSDoP2bR9r7Md6XLg
eYZlawSzcnDCj5xSxI/Xbncg/k1/RkGhBY014ExO+bkwhf2WMFBGGi3SS8sUGQznK93GT1XdAe9+
1NweA+hGMkitAMYRucGqGCHHLLSXiVrvDhu5YlgzHa5CWjXBOtecdBb1+a6AiazH4UoadsxvIF+J
Q039yhal0i2MUkIUkLu/tjPZpBmanRbpVXIHBKplOMBibz8FLLaVd6ReYYoluNdbxfwrn/7ctdmQ
qdeBQO0DeBzoiRkUTred7o6r0oQl9Sw3OZn4taSaa/AcsQiIdueXAjQX4bvQYZpVKgIchfVWJcDt
AgMIOg9Ylp+OSEJ6ISzYvaKta6EGNhb8aUr6LPZYjdXXgL646JAabk4b2tu+w39z4EKwy6tM9PSY
vA0kYSgcGfTP2LpqQ3G2onaEaSMaRJ4YRO7PGDwegbyzEmciME7PBNqrOaxqoTdQ1OvZy8Lckms9
CgD9bSZfGCf3qzB0KZcCVDaPxrtjVNePnp1J6yv6GNhSwali78FjvDvEUH44LiuyNSXpJrOEsh73
1hjF14an/RG2CEnjVQ1rtx+C224zWdIcOTHo7jpWTIYiVWdPYqxZkpjzhkIkPakXpBgfKrlo44wB
ktz1K7WzYM2m2DLkKht+RnJN89agsfXJicZB8ejo+AobrV9YjMeaUCwL3FU6OJQqATh2Fs5mFyPU
NR2qI1mlY7MJ+k+ebANfWvwH7XtP8JUKgl5ztHUWexcsZ/L/xxZpaPLgYeIr7zFsxTheoh4C9vtI
vN7Kfptf1a4qMLOkSfY4TUTi/qdhoaCQoENOHlwahOuT611xFpRRB/GxC0RxyRNpqb7NyOTnxess
bbVM53Yey8pYiNbsWyU9aW3VGt37gdUTwsXnuOBM9DmZSrJIPbCv9vYXUBTU8tBsqQ/dEPxTP2p4
JbTA5uukKqJvp+PxcDkvC5oNIfpeVaK7cWQf67VHNflBi5MW7gPGRF9xMCqb/UP+MwVobxPLWmvc
jLOxnQC9oSJh9XHcxTevIDdoZz0NfsUh/LL+7ZWlfp3hCWRnxv7jC7VlM0Win5vaBzyshm7M1Rr1
FinRXxMauUgBnLSsHSimpbowcSn2vrmiDQKeyu0poJZ+9ivfz0zKPFsWw8/ZSykmPqRpE36LzoOR
AgsHBoOK20phK4TaP4aW+PcUowb3+h+Y2S07b24DAxN/XY5iMG4ArcoA+W3DoTJwijzetH03N1Xm
blaVW345bzOJhWPFlzlqBt8/7xkBkQjsTnDhmzaCDxBdToYIJUqdkVlfqQjbo0HwTHs/cOBFRjPb
bEukCmKUP9ZJPjizISja9F1NqCGEYJodZ3oYFPU+Gnyrm8iJC64PyhuKSZqVYAaFVriCqmoLPz19
mn53oUvXFzl4JsGEX1mnN/gL5Yn1Fkh3vZwEZkIFDRCl0Nk4zdGpwcL5OPTpgxlqRql626D9zw/G
x+vvO0u1QBuOezjUvxQfgZm5q1PTCpS88KdnmyO8Cip5Cl+GSIgPyDDCRavPFG9seaaT1vzFLzvT
hGkDM1Stzw16OLTY7NVJRZ460JPOdisX7Iw997yurFRUwYa9HoWz9FxeIZy+XcRl3iCtb9Gc9oia
lvEhKg+uMJoBe5VkVPTsqhDAEt18anBsSAy+JhiWiaUAycNtn3qp3ywwJ570HBiaRPBZ1b43xZb9
5kkwVVne7PTyqFhXhSbKXhMFA4k9+aIvzZ2N5oNCGRVadfEmLXfhflxBiNNxCzzCOXA8jYXXDnQE
uEFNshPpZM+lDroyoc9w8TAC3Ri2CF0pEnQaVvJpwjEZCxJh8mcF8ke6AUVePKIGT0dIXfKWmWts
ZpdZyH36+mVrlbnw8oTm1wrqpTnCFHHcJ1LH+PALHu0C0Wa12RP4JYDAxAq/w9qbUOlkjKBRE8kU
iBdnVc5XYO856YofrV9xuo4P1msbBeCDB/cgFVDb15Co6kaKFoharRzu//shTNnGgFTwKHNMpgsb
mUoputnGX6adrSHzoawkpclR+KVPux4nL2fSb3tVnEZ7DjK8Fg9GZel1gz11/+lSoZjIoI372SO/
W89D/DGbiKTxPJ4gF6Eb3yN2oBgNqrCLbm5yzr3jmv8zM6zhH3dMPxTKzoUwSuN0AXfK725pkmw1
ETmb/lG4BGUocvjZE+QpUcV0tXiex6wr0Y+4jlRanCb52lhx+sGAccbygIW0zrYs+Y6Bkc1sTj+2
Vk3MxKWGxjQfc+lRE9zclnkMlHtp1bMdnDKQx7BhU4+FgS4egsg2Eo0cihFuJMEVH9GAUw/CiE+1
/HHN1NamXqx2/81BsRgRwaEa2rfzqlrgnmXxioW8s2XhNduyut52BWYEaDjvd4tR8fnfj8gD49hb
jbDqCdAO7FtmasmTxXJdpm287rVo78DKZLePYh8yP2YHDsEnvR4wCkHcVflo55QHGWq9n39po8b5
AYg/4gjS6a6m69cSN4bmcJXV+NKZ2Ur1WFQh7MlRcmp6d88BV8hT5EzPB6cxiOdyVLVcIhtXZdPh
/mbRweVXJgbwKVG82ouTmgIgHWkC1IAi1Jgbm0/Enr590dHLzBI6zi+05UtPWKmuduMGstgUXBhA
GtZHxb9E0i+74LQ0XEu6VHb8D4oXbk82isgK/TyE1L3ZufHUbLuZ5QDOjQYuZ8xfPg3uaH4LfNRF
W32oQ8uv8Yg1pTpgzyuQs/VTP+WHTiiJveU5Cs0Yfxz2ei0qlFtCM8sbuXg/5CH84rQkXKAizij7
G7IYZjSjjF2h3uUW4dmkYYqlPAYS1SEDcU2x9CZ3v5KgEQR3evQFFVGZiOYVU+oNdoCg9cii5A7P
Hhu0VIYpP13KHp3ZARU0MQMz29jO5pAYDZ4ebV/b9q9iaC7iQkc8T0zR1ooHgQZMQZorthO2jbyV
+HgzUw/2hUaE3smn/BfD5e64GrMDXrY8JaqR48LhBGgwcs7Za39UOTt3oiLnXhQ8XUA/CS76mmPL
cCYcfny5zckNtHYCic965kyOIwgEUt1nkZg0IuDyg7Av32o6LFmK8BrUEa9E5GGjylS7NiFoCprP
4Fn+hzcRoylJT/ZlVi18awQThGT+xc70UR5P+800ArYAtqWl1BwOSl68BvqrpHbQ/c4G8kzSlQe5
zWVkCBndnRqYQhkR8i3bbXdfLU/1qgDT3YiET4WR4XdREuVZeIcLouT0jILwWPoeuk9HgbmfT4+c
sTDOn84erdGRkn/PlZLEL9dfoSfuvqlcdb1GegAWxRWr6ihaq/TrIhJdvmQO+dMFpSXqDAMP7KYf
x17MfHqAsxoTEBz3B4mVwpdlpvnf2N6NKHOgOnf+PksiRI7/jltA9VJZXpfFrBIutSPvmByjoW5W
LmqlSk/1JxJHbVlzQlj0KXmM5IBfKMIfqSFRD5ZJ3ULIgJzcVSobQxGUMnhSQr5gQn42xoZGgfED
XjZgc5+wYRqVzOHDKZsQwkiI3yzVOSpNk4Js94doXy1KaHx7ojEzJLXctWtI8d571Zlxt65kyQ17
XzNIiWqF028GyBO4HdPCG4adF4mkL/tDARcjcez1SblfKNecQeHotiXB+aFW9oGdoGuIZd0TL2EX
bkZmg+M8VzkX/Mykwk9aFSbwQgqgcDKObgw/uIoDSJHPSv1Hv4NsSC1DN8Ah0rPv7yk2p3Yhemx3
U3m/dCktOWVWhk+f9uU44YslZdnhk2EunBJQqzzylZRCFuqPD0l0RqrkcVrFKLCkzWfQUx2dqc/p
C+wflKljvpwSVsl466qy6O6EV7r3F2lPn6L8h0dQWKaDU70QLD7FEHEzCKbZzDx7hRoORWdzW4qP
jrEq48VLPCqn9ay0U4n7vxl7A0dgtEa1h9aJ459xoXzYjwqJYQtnElWnOBBsUg1PgRR9z/lu/f1z
quhMmq/RCLPZBJ1YHroAeRFQXTFQ41wSv/7YCTY0SwW2cCDGS/nUTDlKdxPuKk8Tk9G9+7PolXSz
cZUF6IM8bgapcQJ4ZnJ21KAlKGchqj6QcFhVatWw6JWpnV2IaXG7rHJvH7IAslVvUJLnLYQlX7ND
oVW4zjZW+ZIMpQdBbtLqqEIQtG6cUGy9F56D3eJNamtopfHc92ERMxpjIIxkpE/OJ1QN/Gdsi1PO
0kSmFejEw+uSKzjyTAPW5TthoEDsiVyVFFSd4i3KZiSO8QOLJ2fMyKRzC9QD6aHZPxVkeB6gyDtl
SWBFb0RRfNDKKg2YgZ+B5ONyWIQtQcP+Uh1cyxN1zLEMNkoaCBcQy4+g+59TDtYA7TJZFsACfQeS
Gt/y0vxPuHEWBbaf1RbpBAtRL6YdoqdPKQ9xXOio5ByZX1ZkYvWW3lowqrIQZipkh2RMrFNkeu2Y
QXff8Ndlk4sGBgAG3d2ry3RadBKJpVg1iNLm2eSaiJ+jSOOt3YlmkJGLQ1zemffJ/kfgeA9f3yGz
ca+m2hPXZulp7ZgQuDswGq1dtQTPyeiOeK89TPHQUBDfzboeE0ks0tMie6vYS/Y+BRXjsOWuh+8c
WjYljP0CR9b88eZR6W7aDaGlyLZql+ar6kwN8xDheahc9zwwFPJjRWOrWgEdfpXtxsbCqvcoaEp2
ZA4klcJXyosmwHr4bcLPsThWixyxT2fy1lszwyXNHxQ/ZkLxJI3P4CO9AM30pfO5PuiNvlbrTVww
/MvqXZ4OCiRJhYLp2HyCQWk0A/+04oSQxwbIsHTKkhCni8JA5KOABhy5al/cnhrbs9wwj8RcHavd
1S6AfFnnb8OfoupcbOVrgv6GbzE85SeHH5PjdWhTpSZiVBGLdnBukUaob6ADuOrEF2kPaZMY4zzZ
0W+ugSkg6jUDuuA2BnZC19SzBum9QnG+UQTDramAn2go66ilM9QSGr/+HyqOLHamva/466URmebp
okDXhy7jVqg/A/zitCpPBEcGOFwzIUKm7JLDuyWkYl/eDCnduZb+vPS93jv+6kASnvYJWikxYXi3
t+zlgF3SF0lHDxhS5o1z/Shq0lnXB3wNzi4bBEDtz50KgVzjk9oDx/8Jc9E+/756QTgZevhqgrMq
vdpSPq/BBlPKWfxiK9GZhym/NU76CkaIxNL15sDYzMpf26Gr5/HBjNDVrY1hnmb291kewNDb89xR
KwtOnBjcEXBBryQZMrEcNftTnyN9N7d7T+22K0Q6XWBm9gDEYTCfoF+sAZJN9lvp3MYGZfeaYDpj
abtBAz/sd+fg8nbYjkVIbQZuiiovF0TTnvprWfwpoFgfQy0iDxQnIaojsOLpuvRcVsj0QeNQ0iWU
hv4QGGOS5VDBQZFPDZCD8NJrEPXudkLv0p6gUvMUVVcOpehsskclXgBtn8SO1IJbZK1wUgMxxAk/
4E64/6AhgWUOQnGdBgxoWg8qxZopnUhNU0w0QA+jTLFBUzu4m444/xljW3sYc5SVG2gdVhTxXkuc
ozhlypTRZc+rF/Y8kB/XnS7c8IXuLuqz260KY7nN9uIDMv4tRF3wRIIZh0OpC40MK9dsKt9p6x5O
yItngjlPlCY8m0JAh3C+6JFzHjCu5AjJfHu4WUCIgrWV3Lo4gbUlM8ED3pgjYxUHTAKiRS3+d0k5
TXL2bHiIM/zzalpjgef1/am0R+pN5+6ixXFQ8hsXpjt5+N+YW4IMttGBhPiVDGA2t6082IPgHXNZ
Wu2NTX3l8kifoLnO7k88f6Hin4SAyBHvExn5N13I8YgOtmeV8Ka6TDM2400Y0ZawjkpSlgX6IgH9
ntJg08xZeDVv2TXhz6d4O/RwI4Ny4p5LakM4vGVf18pxI84nTv5MypJHWQTKYSH/lzb/7olp2gjC
Gqy1kQGdrsT02I3sgdlAS32+a5l261CDmyOTLk2EOW2GTsh0APoyAn9zuyt67uZ5RjuFLbn5jgXI
8E9RlrWO35HcvNj7sf6ZT00XG/yXBaXNXp1JfFienIjQJcBd/2nQ++gAOdBzNGl5eDc5aX2bGxcl
q4LOI8ozJViKkjVaAVxjn9hy+mcRu+zUk3PfTD7bxpQazf+uP2IJLylYFUUC/hZc4pBsbT8S7k46
JLwuazLYs0C5/4roBn5nH7F0bcI9PLu8RbvB0mE+HKeqU4saH9X9GhtFFA9bsHXRMQX8fTX6R2oi
s1RRlowj0LDDUGRdEErqHkkRWuJaREfVlg3c5VAsD8BsfQ+sfU/4i4k9YuytLNUuTS5m0csx4tns
rk9YltOzIEmT5JxAWm/xRh/7JMAhnwTvwdxFmGk7NtN3MdNpE14qT/iWIsg9WLOKXkS9SqITViP7
Q/+d3dvjnEPNmJlmI/x6/t3M5XVdoDsFbHtjDvZeLHgH+l3yM5pShr/Pa1ziSQN+OfSG3O57UW81
yfYjxpMUju5UjzGFCBcsEmKd/bLzaZ6ShkQZCHmca92nrLXL58O/N9wQeYgu5o9ABYF9bATGpVRT
2f5U1qDCucat1mHMy4cGqbx2VODzc/1/eX9JD/j/4nzfPs/QmWcJNf5BztC7N7koK1gCDN3gLxv/
cI6o4qRlQOrP3oCT1CesSaJk1BajJKBY6XpXLM7JtWRGWpiaBvuyfA2N3lc2k4sVgEBrgwDfxYCh
2J+3akSVeokXPg7wZGekBZA/6Dpnfgyt5Ml+y/y0kbynN146uDL8bfcFR1kiRLZEW5yQMLOwuC92
2dWGF3ynW6wGDtvnflEGjQ9aVBS96av/FNrGs72LKeq4ywJ/XCSArxnkZbmL0IN4VkrZrdg3oHu4
AcqbpNcmC2LXVzfyJW0YRC18+jJVU5nfCIw++k6YmWUbpluvNn4CI7uoywHk9NwQdpzfR8EY8HPb
AjFGaeqdW9JVD6zg7LaO2ycTuDxsekyhYQ5PnWtn3oCchZRBSezZqZyfU+N0jWEBFcnkUCz8Yn9a
IAxynMYB4eh42c79IXJS7kdm2eC79RevX4OTrVICWIDRpvAA8+XPFr5ee0R56mvwWe9MUHz6EZ+N
73F7Q2xL47zE93zN009Hi/RLNh/CCVy5QSPY1aLkl7WrFmZcSyGqid04P9pzDXibX0HNLJZeyYiX
RJuH1wxMHdoDF3tkhWUNB7Va8XcvgqwmRQSjQOqaQcVoccRpXgtic+IzKa+hsEmj4lxJ59xVMN+4
Vt3Ax1hxpx3GOceOOrb/B2QPIRJwH1bXlrmzVj6plh8XonUnYpCzXIUy1wcL/0yJ6VP4RZVMcAk8
SpGtxnLkb6OSBR9L0honZw89xVlhOG3FMowy+34QgToS4IyS2Nl1zh+feCOifCFeBRD/gMo/i34U
Jk7F6PnKqCUaTlTQZmaiA2Sk2HtzXB6/17Rq9rnSziwxnqFQl4HvGUhCLKtYPaOMfhXqHxWCeFwX
prBFPcPwi+D1FnP9kjWTFOLaYeYpjKxtLO2oMohwtKKIRQeDgajWNprllPpKR1vLT4JFcvyE7084
f7W9Ilpj6WWWF57jsiyD7vY9jPoHOZbsGTWV6LpMvQfj/ovLcHWi9NIhaLO5ZDBH1fral2bre2rT
MJQwfX7ob1+olGZ7n1D61ozPrF9IctF4F5x+TjpvO/gp1CUWln3zY0N39mfOFFgakiir78t1StfK
OiUZejP1ybd/ywEygpX+6Ed8/1iNgx8MfWvbvzPeMR+epWwpoDfDJGkw6CyHbtOYsxxJ8GUGA7ta
QoFODqeEVcf5ikSZUDXvnry6peiBIvN3fdHzRx96FDgEd3+eo8yXb+Frw/qMHGSqBm0ZBCv36Kd/
BOImrhdyhGdo2SiH6hb8kQO2pdtUcqCOHF7CiBfUJN4QSo3adKHS94O5vLIU+Rv04bNBDJ+oY0oT
6TRD2r+RIMpw9tpwq5WB2vtaZTkByQ+hGL3jf31oBQImUbncyCfiZXBXXXQP4MelZGHckwE58N8C
HCEifZPhXDjKBQ7gpuV3WRofKo0J6WSUIYxoGxjVZb3QtTGdspwxFBVyEe3erKc3o7PtN6yML+VS
WzwpKmIkngXlQ6Dlpq85Hf+GVALy5LFFGA3OpZhTfSHIk/76QY5siDUv3i5LFJjvscJ3wiQxkIfB
nobcxfevqk9WPT1jpqILAi72iRQ3t/Tphzn/foOQ3Q4kvXJ++M6xJikNTlss+GaAgLJkbxwjRtIQ
ErOYyYu113UXv1kiW9AyPMp0YVqbcJJI/7bMMC0DQFb088iV27U7KRBcnLXetzQ+kBtiD18WCIaY
Xw0CedPh9krPZhugkI6c/K+Wq2gtHwJMHGsNXyLKXUEXfDcmuC7Q4zAB9Hr6/PHVkujuSNBXYEjR
hZboKHs2q+gmdHK/GSNQr9r0jvCKQ2GUlfAd5tgWbzVeyCpTesBGj73Vc5z4do6oiQMgeosYNu75
iB8tamP3Tfzg++7xrufNZ9LB4qsdi0KrgKkqX06a9Z3oDUk1XTBmFKQU8Xvrfcf3tXFuD6bNItkB
FxQ9d9TPtieii6Lom2WRciLW+wmDT9rN065rBVe4Nxg/EGPU8FZZSa0nNMmXbzIYD/l8XCChqP41
+f/wbjWdCXXt3+257qGsF5lVHcNlkaE3Zf51QaDiOhotcecJfFR067Ql7felckxxV7aYmBwNwiKl
1DwOvWwkl6ULCIh1neebQa814peMuxEr/v4B8/rkFpOuLiuIPom2taDP9FfQH7SLXmjhah0fyWn2
G4k/cMfouU6hTFEPq9007aZwHAYthMGKlxPfuw2uWl1ccixAkjkNl0yjfQSEApW8qJfVUAbsSuIp
G3wJ9o+eYpv8KCL5esGhi09/2UFa6lWZQNIo6zpYG7JerL+3bMeeyU46t2xF85GMD92lTVT8xHZT
1EjDQSasN3SRltdcanqXlFmsxTAG/pITEZnwn4c9tJrAMOHOQ1ZFbogyoIkl28W0dQFI1uZ99nPl
cY4enaLeWHD06maACW6qKQQA0Lar+SAM13XZ2fnKwwOzucBkA7LPTpE/nu/UPc2dB6sQKsrKeypv
n6ozWRxHpnL85NR/9Dn3+KsaCD4aiTWaWnlc0J0occUSAqmp25yN33zahlGPG1okH2TBL4bgRRgg
dZsEc6sYyRWFlnpa38MXjX3bJ4Jwp6Oun/cyKVUMY/Uy04RD7JDvO4VoNEI9F00Ycw+CvM/6bOKv
Ked0Zt48gZpXzTeSGL1GCmgc3+4F4/K3juxqNgI/riFdvWK49C5ROFMaPcnkXDeVDcR1bQkMONIN
2s0qGzuNhF9+FB0bxZgPwIVYdzaLkuWBFnKQVnJ82eSHqqWpQNTSORURjPsYzBlzl+Ci88Bs6ucH
ohbjOdoEFPnft8y3ssE/GqJKUUQfaoWeV6v0th7fLJutuThh1W6+S8Fr3c5EHYauM7cLZLBzolyA
owmKMuJ9LqQo7Jqg2wdd9pRpVEDcYeAxLP7EDgchI1C5OKtrLA/9XnCV/O9q5hSfbF2kxmpwi+6q
ZP1fJXISggBdpUN5WNW4SJLXdnJb61gemBGLiZzndNiovm1CiH0k12lzqPBtcPB/oqwGNtZeBSFd
6+8Qn/OuYNjOqPK3dC0UsOQjGfwlvj4FHuRq6mBiWxswAr+AI6doqA7vrr38EC3lO5YEQYJrkjVS
p3QNovW78YyvpDdlUhcjnBSuNZXpENcn4DOfNpGSPi01K9p/NSRArvlBY4debXl++uSONsEKKXAN
Y2rD8xELGcxDXrhhH5Ra5o7e3RQIYJLIvkt6UnKj79cw5FK6NnAz2DkhnzyDfSPxfOeaDoHrh/Bn
prFpsnbC0lZP6WoPs++B9o3yLE09/jOSVZcf48S2plfPUgb2hK25qHbLt6c7qY2R6x5yL5G/23VO
CJgJ3QSt6S7vyJbbvhh6z8zNj9vE1XViMnHr7U8PsH5OLdGth0BUThhu5ILTHHBZdjjLf9d6tP7C
IJw5Od++XW3H3WbYrIzWLP1kDcMlsgoVCN4MdJ4Qrr0hTmB4mXV0eOCE4/5leQzP4fQybmcg34Wb
EiF0C9nPK8hg+N03ww0W4kO6QpaLGLYTOQ4bXAjnAmgnzdO4xNiwhJdLNJMe3nbKXsHmdtZp77Gb
Kj+XrWF/ZnJDXlHxd/747LAAf/lH/yz/n/r3R1lnLCKPmL4hkQfMxbNR+JfthcI4MuRehGl9YawO
vS+/qqeAuTXZe6ibKOR8aWiP/9y6jRusA1/DRqumOptB4i/ZDKqyJtggNaK8H3IkCUDgVvF1y62L
W3dUsn01jwbEhDLSvzAFIzexm3RDyY/6F6zQdujYI0chZHb25nAoW6HpzEhTtlzPOMNiREXEEqOk
fFzuv+Sk2jwHEwtwmWuDltE4AhtYRxMGhINLYHW+3OHNYk1+F43nRdajvh45X+QXTFSrv4/CBRll
TA2QHHf7QlY31BHmYJe7khVuGKU6tdQWzCFO82kKgoPcwfdb6Y+7EcMzGjckNZjd7s7YBwZrtgRy
L8qOcQ17Td0DAE+aztUsWGHePb6TYXP2ZEOU2yr83Vnuso8bHKtIWaypF4BQMfn7U9t5vLGSRd/x
8wG1wjMTXJRV9khx8S8c4oZwB3xew0ReNfqYuQKY2Kyz4vf8ahQAoyOVULwXbirB87rwS0nbL5tR
SmQxSZvP+YeoB3/HLOw6/gOeebrr+gSw/JyZ0FvsJY8bqHe29kfBNcnaArOOUyZdWsSFIZQLo7pQ
3NPs9Tk16uACWzZBo3M5JSuzsZmOHPys4xoUeKmNVBqGxvYNKeTXKlMtNvEh4bdmnrc/mByzrmDe
n2epS3zn2BQycZ2aCKcHcXHLwR+i4t2luhi9tfJ3D8CoSULx3MMtViVPBlYq7HAM9AQV8Jbk84m8
bTitbohUK+BKvKNmQlhbXspgihXQfS/ggUDDQGCjPFH2eptyuxuUgLrprLVAfOlJwx37868lKQFL
8C54+1nJZP4YrWzbRv/mCLQ/gbAbxO7YcLvJ2AC05TQ1GtL+la0yzpJJkgGGnMHaaltNokmzZSaN
W0mBxuTjqBglyzaZaaiVaPkNpozW2jgm7Fij0yKRkfkhSvjIWRxhMbW+bmFhJqg9THsh7W0t6s+j
Kh3hIJqh7IABXh7SxgCLrWFp9QiXWsF28TNuiVTRrojnMQXxNpalPVh0MfOm3IQAydeIwAI0Mv5R
iVYRzsyrGePgxJvUqasaZunfILIefO9MdrF5LtHwINw8aqUi+KNb5podfGipd7Hirdz/N7QMpqTh
3HOpGFrfKcCWEXC99w/UYeEAwbdT1R8iZ5vBgod5bmzZqQZlXuS4mD+x6aZP2aKjzX3ir+VMxbCy
Hfnx3iZ0O/qHqUNypBtsx2893fubICFkhaKxC7iDRWt85qD0ewFaQ8Lx3z4LYwlde8tt/cZ+yUle
0dL5vb0dGqhQHRJqNKBkQfXj9ufV7Sr723Hc4T1nc7e3mG0ld0iuKGt8YqBNzXz3+lK+X/xXt7cw
pTy771eDUWJAYEfQsSNETBNbKteQN+yMwHvUHwM8v0X4HXVrmnMtn9TmsGxl1QmzDnKufh65BOvA
pP22MXj/ez29af4B0YEKXjDuqVw4cS+jbWgtHNXFglMFS8bLK1Pg/zX7fjy73kQ+KfQGhny5NzUl
fn5244iSny3Fn0wegBNovxY/8PrxGoe3zR3z+3r3pOG8MBqKgl17lcU4wQxFYKwcw3erAO72DzNS
SUuv6BpqdL3R+VOkZLAO5SMEazkqWZYV8zcasZvVDbNT3y+5ycDcDWK6xu4fEQ1N4s17dbuK1eA5
oQu5htyxZD0wvKhDICKG35ilF5a7rrGaFpvAtUITSVNrJBFzq86wSq4LVMRKjLRyIsddns2gupTB
POJyVBruBuVG9RP/8NoDGaLkdU6MiBuE9FOjwTVWlBm98tse9lWXQmYZb9bSLqKUpFWzMcQk17Tb
+nIMARW1z0FtObRhx2+vBpN+4D1s08bCcGkc7OLxgWmSHOHyOMkYH1va+ZPRF6VJ8q5gMeihlcnb
r+wpCGosj7zLAL2DxDouYliD9YNZHyzUSaJGMKIex/0Ji6tzgM2HLrUvhispZSfoITjv3XME10N+
TYcGTWv8LUxbR8YTtERoh3f/opCPQZhgt9V58U+wVRDEqbl8mXinhrHdnsxYiqRoe7F8HVfh8+jL
ts18xhuNbWn2n64Y0q9tF163wzqUqe2++/NrGYQ1r+8vLOoI4BWm/uXGWkuqnqVjv+ylHF5CXzJ4
HZAffnzuotKD4ENuaMbonKjcdT6ksUrJ3TKzU2RXD2OYnGxhx+/QoYGa5Ke+v5zzimvd2DnKTzPi
1R7JAvv/i+qkWh5b0CqTb9hzSzlBZINGVCffds0+YaV7VmH1WWpAJHJAbA53x3ln0XIU7zLJJOL0
BmbPMiYuxw++EznO5H/oCf6MPe6OzWUq8dPLRzgkBIpA62Jh+RMh234zoX+HK7G3YMJwEkxx2DhC
ZYuKQIOpWCkTlabnS0B6Yxi5LokPPA1TLYjzAOQcnCIa+iQPEcpItISWqnYZQSzy8JaPyV9JesR4
wqo/ZRY1UIahRj+HDghCKXe/DjcpNfXrBq0r15DM9gg+xQC0r/xeUpVBMtbApUEWCf6u6hsYLZ+B
t4L4ojHECscH1kFK70VfXBtgJ3H2iFH6tgskmEHqJSyTgymi9Kb8hjykl7d1OP5Il6ObXqoeOE/u
caQX0dCoA7BuE3TzHR+OkmW9Bt2nR0CmO+rQ+NqZ2JbZM20AMvVXLb0y3z0zJ1PghmOVqqPhhO/F
hi84LTx8UFr9RbwCO3NZw1phdwAxfrdXTVc5ovKW1Opt+XPYx40w1/mj1OzGV4a6UftqhaFAh58T
/HxsQw12j0GgJdpcqxcA4KzeWE3Ppmm/n6HTG1lDv7nbPmy4rxKLM8AeH7iThzE6itARpFQ3S7YK
UHlRg4FMULhewRvx7rjwyrxmC5bKIu4Z8Q5KehJaRrTAxBHRqM0M/WY8wR88qTlSsxleX7Uxfd6v
uE3EHJb8ZiRN5b6iHjBRe4uZHdgCOHFNsf9mmzqKbbBgp73t3dCeUpmivVpvdDzsBjA+EMVpfviR
qR8563TRpa7751s2RiQAGzLE8Z3ww8MzHmyuR66fYLs342LS0IN5dwTy61iejDOVcoFgh8TG4+iF
mZd7qzaR0tNktj2+kp9HH9Rgpdii2i9dRkqsWfpTB/iAPPDWgiteFZrak61NZahMuKnBjL/IvBl0
F4YiBUJECHTo+DgXzuBzCqZNLICvxLFNfurUVUpvsQcj2OD4I2M5D/vyeJkjJaiPOXV5m28SAdwX
POBylznV7Zg5eLStb/pRtYO7YldwoLcRkyuYR42hTZp3Z+U5fAOfR01JXh4cEreaqJRSVGefzd10
HjCN21IUhRjYpWJgbXOxXtusZ7/bh0P1PDEBE4vn6dPv98fsptvI7OZ5ZASWxzI1+8NqPRtjk2bw
/f6Aeyw75rUPBeid8H8E7n5LUD/PKRynvdQQZyXCFTR2ox3w+U+WNvi20r63+oEjANdAQW2gBrnd
k5BV324o2lV99WSYvuT3fgtt8pkOFj58v/8i9XkEwqOIEEOHTdYebKGQL5hjegfC7m2x+i0ynjSw
lCpvUGHXIZj99YXGb+KGnYSCEBzbqSxSij9BXXl9Ng/RAj4ltYulVPLFnRBGiKpKPLdRx8NgAmfW
jZCjbmgIMCDMliUZmVzO8Ks15nELzlLmkHxZ2FghP2UnPSsaKK+9ZTF+Tx1hcJWwEvZe5J294lhN
SDdsLSE5y1YovmTp7nfW4IDL8vzkk9pOfj9xAEAs4GSKlAMmBhN1LlhZZL6rZ9RmG2AwIElO8aLI
wT/CsIcAFPrNrWUVOytnGktRFH3Rxlji4XWU30R6OkHlCJp+BV9blCL/CfTI+eNlg+iGTNQFhmSd
zF1BHjJnp56X5mp6ebO5x8VFBZccZN5sBwEn9OfsPk3HoYFsC+PT0KOlo1RXVY2E9zz7XDpd15yG
WBqqJ1/ypGcXYFcFvgn4B+uT/1pOrotwkufz42DLh1JwfAw1wp8IRVfK7tXO9cxIqgBVPBdvlVxx
c9IJYzZihuwYCRAZ2iPFFuFwT9HjGSOUIVW7PVoLzVlRswV7OUv3Fm0M8bW2fsnU8tZgDixiyOmp
lTlJxdjGJDpqkXizJ6JmyghRPlF+sCERIJe+CVhlwLKlZ722Oz0rbOQ/KQGDvUA9KghaJQUAO2TW
iIAkuf4h8/jw7oufwJ3IBKQ9LNipP2CjV4QOrrMZiXhQKbuXp9bybr2sakSXYrYnd9qJZV5G0AFt
vZUScZ8kTCa8uY9BjBFiaOId5gCmOMOOaX+uFFM/DD9jix9HWl6AVLmy1Ncj/m6+tqV/ozgVjqrk
k8tcxMKw/3pioXpk19waWC1QzNbR1rq5034Ci80lSFHStqv8JB++xEcsZWrhOiApSUPiguLTZp8v
LCoSYNoIY7hT2q1n+Qpu7CXI9ceNAC+i2dHmmvEwQ2zniqsPgYrL//b3DOZkKJtLGtNADRr9MMkm
GcZvw1KNyHclc09uy7QG1XBIpMKiEggllYrxytNlbJrJmjnqK7F8N7jQa5cJeoS22/lpexdKGmOc
O4d18a8Ru1XBrRQy3RvJ2CJYz5JN5xB9rc6YoQ+wmdwHmDWgy9s5bEQFW5QpDb7+UsArrnWdZ2wM
Ia58BtekiBtc050ttV6i9BP7mKh05Y+F6fLgtioEAwSnbCvp8hQncX85qXhrHsyjyi4Jw1082H3z
m0PnGqOPppvvbHmsCNnh9HoiVCB51Ys5N76YHXwtJWJTUYc5VAAJXztpT37XoyE7Q5ZvJ012ZRkN
4HLSPc8uFv9dqp+m9kVMGKjLXBai+9LM1yqVyATxBv5lre3CZK/a8O9pmwop11SJ7hf0QBmeXbzj
2gVAk6evkKuP+p4X00clfsqpGSYMTnQkS7d1winKQOVIyQUW1pSUKn+KBxf6SajlAgZ3zXCjFwMQ
EcPTYzexh44McfwkziWVwn/zUMSkeWDmjjJzEDbGnKn5+rg/ueTtpohmUn7c8d3ehPjW3vNYeAEo
0rcSYNiwMy/XM41tnPtIwrEnMHUD4/r+SAliCvSljK523aXw42T/mcJLhx5qLyHGqVqX5m0BExpC
0jODAITctZ8EwXIB8MhxQiZzjaE3MYcWwrALda2eKYfl/AyjL+++a51mb+EBy7R1Wba2VOhjlsJi
JSy/BDwStr/wL0wzTp+Rhpixr1Cx2qHWKeYMi/Yil1LX1DKu6Yf1iJ84pB55a1nAplDu6CKgaqcg
CffCcu6HCIgjNHPmw/Rrv2AjjheDPiYBjaPl3DtG97OZBKPiGptPyxbM9KzfMFXP8sC9MWignVr0
2oPcrnj3n3Sm4sB9dWn6RiWG4BDxHyyOTGUYADFg8oZuwHP8zQZTe+AFhE0B6J1tZqp3z7HaHvCO
UvPocZ7Gok6V9d3bwtAWu5C3ANwBKhzQca5ffFZvUr1828Pi9moi6+VrPHpgvamKLBMn3N7g3ZtI
2M29ZstwLs5mbvJL2o7AxXxFgVaDD1pT5KUC4yKImqdqt3Skdfo+qDMCdp0B5kM6x3dMJxCZWnWa
ztIwEkVhE7m5pWkoQqQTjfH/Pp+1P3zjQRXDBMk88V2V50LRfeDtr9SzukWQiNiJTmhF0jEcoMVU
vs/o0rLOER1vIUfZ7pyaUr4x0lL3DTGy99hJT9MYrwJoXx60IBNoJ7iBnfWv0NaTBDSLlKvL/xAp
SFE5fa5wTWlrHm+VxHoA0TgznLq2jUWZInJkfJY83kxVso6rjiz77MSildFKZ63is9pWS9ZqJ0ci
fFMKuBf4AFMrxJ0e6j56+Gl2QymzkvZRo6aSQKhIY90ZfVSFp9ssaVFr6Q6FmgnLcaGLOUmXGab6
S3ZbjhhU7nJ8AlvjgORNjTSQdDPCHCAjxqjIFlZO5TysPP1VOEvDJZW62LUbK2y2cB38iXXCFh/u
z2friAQ/UeXttF/AxQ+M0gMLZuuYxZLBwM1NvKCSvGfkUdMf/Z6Y7EQuOqaNRIRETqfhcRwV4Irj
JbWfbOynNY5aCKA3zjAlx7OyvKNyGmF6zL35m1lEdueNWmrg++k2Z7L6BHr226B9U563Md8P4P7Q
pT5e5pY2MvnByBL9V9X+oJPDnW5lMV4whTlszW4d09ChvM0XNa3zaUEPcFWH1k5GqQ0FjRIKYGLp
W2Ut/L71U2bI3ERZUNY0MCTh9v2n4nNAkmrSClkxlbInp95u6jYSwJaM+2tnjibZfC+Qtfk2CdNj
Ev31ZX2LXdrWrV2HI+oloKcEB237HMld0P+F3mphDHquJO/4OMXNilq+r0vyKpG3ACSPWMi6u5NA
kpiMuUBhABcb45AtsQD1h6THCOJ4cfgn2Ee3O/fQrHeju6PbyCuVUv4GDZrWU/uPeOs4HX7RSdWx
aUImiRPKrjlUpQ7F/rgpZGT8EjunbIzkpdv2qyXsOzJJVjCSBZLyQqQRiBVFecUQfhZMj4OFOlqz
z2YFhcVVA2ZryocCYq8BD2ofHt56vZPar3j/csV80uLURXurHaP2tSLO5ra+vURM09W4pzbY5p46
2BNAids1L4uicnF0la0YDb47jxJpeWL9cN+6AQQ0FfyOC6YRHKjefa8usq4iuw38PahxU/36yzb6
b08JxhSfWsbkdKbudED7sN0N8GMuqCAiDzV4fm0bgihCqmeqevgMHc0/3tdkJcdGjxx2MmBTRvQQ
ZFJFbjfTjhGMcQ3WKKGUH/VpF+t7Im0nYNEUNn6KhvjDQCylW4MOHmjiRjlsVOixJL5D+3cItOOh
Ydr6Lf+a5K+GVPyTBFDS4ATQ67qf4LT0yxxD/JlkAMv3IV2c9pDvJ1xvQl/uYriNLnFTyzoYGnvG
gwqzkDumF9JGdXgG2I9oSpl4XHRnz2nNeTfxZHmay7XGEukyPDJDfHGnqikBLAxElFEHpfW1UQcp
YG8EjoaiaXd6mdNRYjcXuIJKPr880A9YX4l8g4D45Qx7QEGNlFIpH6m9fffSvGJgSe9kEOA1+pwK
BeXYLrgrZSX2sqSFU9gN2Rv+0LyUGlE0Z/Sylm+9l18ykq9X0CtNp//HbfXhWMSFLIIY/FcG07/t
oBeJiL1fMyVYMZki6wch5nmt3rQi5CJSIwETjIUp6xqwRSM7HGr/3YjOfwD/5EPT+F8HViOVPpuk
KrGv1qXFo8V1bHhN6VZyZoT6GoSQDnOsWD/vCLIfjUxhvtNO54rlicLJ/5lREXhCqz+vxRku1n4L
AYcgIZDhX7NaftVzn8wPsKvMQGvw7uNBTlV77RQ8zwk1w1a5qGj9hiXZW+YaUPNy4yYcT45Yl5BY
MLkfWefIHOQnwaoPlrE5Xbe+Il3uFz6kgGW1msJh5pdjGJJ8hTkI9SILgUoIDrtE7FczMc2Ky6jn
83JBNlUh/8idZk98CaAgL09aUbuloHpC2Zl88/HR0Dxvyu/vlP5eWz5x/2B+0wkEMkoWn4L0w/Pq
0wb46oAqzioJxNb7t4TJvr69nVGcmDR5693yR1fI1Xk3ekYYm0Fa30jfVmNbyBrCKkgIiJbodUdm
MJ5WHll6GlAIVSTapYXrF17HDu471WWSgLkjJlVbP8gvr89Ia9y1vmL1HSdr3ELnmpu1Ker37dsV
fXjxghI3vnz7tAkP0OSyqBL+k+F3TJGv1A9IkZxPGt/FDwr0Ahs/HfQbqd9MH5JG95tWprvdQCHY
7XrsXZB9RjqOMTMOtpPM6YUcHZgKZDdiK8br/uoJQ2zUT1tDxoRUtpOw9QcdmESs9KxePYOo55Cs
T0W2+fH/2+VfRAbdEH9Ob/eHHf7YvGq2JLzjhRBhPUIYvmzHx1Mfg4zD8mUhPmQocgBmuRGXil6t
jttjS6I1eTxaoNoUS0nblHg01/2p4pwaoE7+f8VqnzDhw67fzaefIB1C8QH7v7Rc6+DJnW7Gjgnb
BB2tOSquz0dD4C6eBCi45Bw65NVarxipdiiLREW2EyV6FtXeQDrmPJZulazQ7MnHmYE3PTP1e4v8
mbAPHHW6P6X5CMUaZ6Dm7msXP0BgThS3AU27N7F6/CJ9fF9epMtny/x3mXEdLw11lBHGbjuyVERU
Axng7rp3kbaKIc5VgQ2bdakujWQin7NxSS5dY7Zlla8dhAFkPegwoB71DgDcPRg2iTIKeViIBchX
ed+5HzSjZVY9jKRYm8xD4lozczb8lF7d+p/gSunV6ENlMNn7yByLGGBF5yMFpxs+c37D9Q/bVTtO
1DYGEO3mylAyArIont2w+LcNboAdLYPjdxOiHj2giaKLBeb1pVBx5o8DDG+LQlJmj/osKh17lNCA
L6dSHiY1fBdTgno1SOhRNDvr/qkgaCHVgdACLm9ae/uNRuyKEwjDLAeCdwVNLEHQHot2wIA1C9JR
uhhbSjgsd5lP8idSTN5E5ZoN/HMN+vnAADU+xT5e6YxNVvLP51LQaNDbmHgfYy1Ai/Buer5QdH+O
TkyHHZHa7tT7fe3CES73q3p/j15aI7sMZXol99WsHV+xbkDsxkqY31czHShGf6VqieSE7tYvZeJb
t3AxOT6Ex+G4AgC9jzkDULeIGDuLZkFSa8e9+F29uujN6P8GP01gIOxSnLc/2U5qUtLW/bw5Yu7j
NvRFBp+i8veeiMcZyGSI3DTWCqwaF4S3Vm30xdQwmYtobPR5GOIKw79O2unBNcvzzQq8x4qx5QyL
g1S2lY30jTulYrXckBIHRisBNtRI9a0StqNz7fjPKqNZBIkJHIGOxRp4lIMd6dahjgDhkDS9B/m0
OqgyYB3MHo5u7CQ7vvfFpik/l1TXEB2cbDe3FBIbLd4PmkHj2gv4U0gmKcmJU12VuedZlcSqZD0p
ZdbKOatV7hr8CqW4PO1iwpB3hgjlqL2lnIxLhmvtnZ0kvZU3t8J2UjN/Kuz1n0sRSrrHWqXjANwu
BJLiwt9GObnL3RopAGnAZOHbj+dLZ4qt5+45cUA7Nhi+0V8UzWqXS7soLyuxcE9/XZgWLqp3/oo2
YkFQe9aFR4EXiuxPw9Nc9GPb8i7x7iNGdn9Adc2s9cYQUN+G6eK+5BqPSaP8jmLVqS06kci1krTu
Mik+/hN8sYUOnlKb+BWhZWzCOf0MWc5sy6I+D5JS3Gb7WCoRZUMBv/XexRi0NmUApi9hM8g6D8oa
OZSjzSoN8ll2wbjSBCNgnkn785Ok2mfFNAD4vzKySmwwiZw7mhC6pUU7J3drCtEh7ghi42Yrj4jx
zTc+DMfC7YI6x/lV8Ya1jPzMlslnNUFmyI8ddg+7ReMNVxQL1xNWzxMMjywVB44bwFablkGljizU
8uNIAV1O5wnASh9Wa3YeWxIXZ2EuVHst5+NTmEwujKnfXYKBPuL9ePd73kwpQQV2hBg5NxxXUb52
nbm7lB3iXQsPmBOI9rweDp+bDE3ysAQT+jVU7HLrly3/p2TTuRrsd+egN/eeKXXZ16AmaqQg+sin
mJ1yVOs30haAN9/Jt/U+1IT70jbp4xBumVmgBl9SDg71NdxSfIL7SCXq0aBZ1K+HGofX98Tjru/w
khKm5caqyZovySEh9aBdaSj8VVZ75c1NUsboET3K3/DNxp9gD4IUxIdVYM91STm4tNjMEcNpxdcH
gRrImbuCaWvrP9mAhJ9DyGdRtT2eV3NsxlOwfSgTWzjKmrchguLoqjPSegjLbzc1YKY8XBiR+WrW
JjNf/6pFgnUphWyqq0gRE0bQ3dAPmCQJWsqQ4wYM/jOXyp0tNfoNU+/21Ts8FqcwjeZZo1GbwzXh
svHRH0v6Tei7l7qtCQ7ZrRHOTpq0DNXJGsOAA+DZSvuMzFTx/kBXAmvo8uQa0a9N6333QzWoC2vw
m9XN1b9RRxPPYuSgIhfEGxO3/2iDUJtZn6b3ZPjEDt/zYEWfYTC8lvAhutK2d6zF4rTAfqPvwdpH
ggFhCL8eIjVep8n6UoXVvsPsgBfYo6PBGN+sQ13z1w4OzGzSRx0tLuGVJL7QbzxkMpVQqlODiFXN
tdP6P0rwnIzyuskNvVixpp2vwH8DMsPeFL1KlOCmoxvtUj6MvxnW/TUrkvhITk4MOCEjpCbtmy9U
wVPueH2LvbJHKP/LtGHd9UHwt5Stfj+DSpXMVIS2GXZo1nBNzeDNcy2dY4c8Tyz36kRosB9ccqmQ
YuW+Uxp8Z09l6b/BI4UEMWDavnaG6oOfbXkmklo8TxHNiEg4tm16dN1jzCK3Mmz6KVJ9SXGStDiR
juI/mnkmtAUm8P5NtMekWDIuELjycskuqkwua+o88VfccK8Ym9BOALICjfCxQ4cDOC4qCaTMyWuu
XYzV2tUMHVTfw+hR1ib0DuGHFG2Vg3EJkIy+YhiXRbuSO8+i6hhru2XWsqnzJtv010KpgPER8LYZ
IC5yEgMR4uIyEpJTpSmRPlTJ9bEKa2JN6rp+XvgtQJlINNgmklbusE4IcL7Tv8Y9o9DrAaGuH7Z5
xnXOx3u4WfcSZl6M3HXk+hdajy/Mp5adPeTzFV0kSmMDEGJOrBLRO3MYdE6EZbjHWcHIMuO2ftAX
mPcmEa+ffs0wtv6UdyvQF1pinRH5/g5exDH6xYlI3C8dytIb+BP4IwrqPlCRiHGdsvaitPdymYAa
KOnVdgOsHQobNwPrZCCqwUIJtVkiOflo1i6CrYnKx5JqWQu6mYA2Kx0Cmb3mXX7qUHnrD8FL7lFR
hE0MWhTr+anFWEmbbS+43XxVW4OLo/8J0Z75eLe7ivOf6A25sG0jaGcW8jkLYvTEblgJ6YfFTnEC
5soriXEn0lb1LUFzqtReXyxdtcM30fNVtUtszsiD9v8h5qBSE1azSZPD/z4AdGEYka4o3X6Ejfmz
m8S4oxnC+p6T7iBZDw5VdVRAezFehbQTNlxsGnAjSOBvZ1QgJvD1TY6VQvvO3CnziQf2RH1PMr1k
QZ6hC19uG4ss4YIbZbU0EwUR7OfsuPmiJHC5+D69jvnFl+c+pOA0VclF7uTQ9nIsUfsSvi5RX4zr
4WE4ryWDArs/GPZqT2JgfCzH6vFnGK+f5eelqs+rb7q/J04xgAEWua576skFLkIPzmQ3vHpzSabW
sDP+g2nmOs3cbj/fU9Cj585GRvPwXnRCyDwWDoDZhFjyteMRmyKnqKYCgtM6xAar1s7pilRscB0+
qHehTij1EBfrpfLo8nw3piQtjz/3ddqqlVDoeEYbc43ttDprM8YIiJRmv4kCB6mkgv6XPocHBSVn
FoST0ZRy7FaqrQOUaksna9pHUjEHDef0pzAmFG8rsaORGeLOSyR/o45t7LMOjfTwHBzIRaDRWlFN
J2ynAcXNJQoEuJxZ0Uefsp8V6npjq+UnM4f4FP/DVR+g0EwZ/dqOoyIaqY+HFY6PaDOwo1HzsyXa
rLMZjJbTGZMHHaHXXII2LFLRaezPisamzxzFWGmB/e7sikiAR4YSzdSS6VYGMUpni7QdmLVmZq59
n0HpLx3ybJKyA+imB2N3fx8rv/uKVo4zu0WCLolww0nfX/PVBW119qKTJLawO7OfFcUacZ2gordL
aPDtV8oWFdfwkoiOxn6mlnASJ45i/V4DToB3sKI8x0U1GJbyuxSpMtuHf6cEbfaavcDy7xmOTCSp
fuSJAVgAk85rnImHEwfOZZIHWavlFZljhJ7U/hAQiyn9VDI1SBV1wifatz5j4FKjdZCnpVojLOZq
wGQRziRWpNtJD1wjKzgkHobCUhqqrgvHaWvb5e365iS0Jkh981x2w9XfINRZg1nfjgsyuADE9rxg
hvcFob8DpTXOPsyemDVodfXx+Vf2t0YslYa5y3dRHaWHE9P5jZBVCvNt2sfifOtbMW8iZ3jk/zb4
6wveD7cE7229XxBT2hJbJb1os1OutEYuU6CEwx3LuO1RTs1ErXkdy6exqVxH6iidHB7i0jvP7ztt
nBUd+bvSPzKg0IMSJxLA7CxPMhjRxfBXlYTl7pLxQXwMXH6j+SICKCmRGnmktDAnFiQoKApEJLB6
xzj0qHBF884kBb/B+SLNWVqxzinScTCJG9xc2nWg8ORHULhAKUmoHxOiacV5UnZ/0dNcrf/u2z42
Rbdwv397AohT3k3uFULouyWniSv1YJBLw21PSnGWV/cN1sqilr0ZJ/H+U91XBMxhxlokqDhEbyTx
AN3PmyZI9h6JxBHqsfGTmK31WBRCUp9Uk6hN3mZpSW1LpF0YrFgzJanurKmtjbOSz3nAqnntVksU
n0r6gv0CsioVYP3u9eXQKJ/T2J4KwKkqzcmY2UnD2BH9s2rsK5xS5FVL4N0uwJHUXlLAHouhuqne
K0ISSMW2PBhxUVv84r7VfOqEf9Xd9im+M+KkkRLQVPrpNpa2Z6rkKINtPQG94m1iQB1EkxQAYEqI
SxEqw8FIqpxaoDHf4yhfKGz6bUOpVrGfQxmH0cTim0bDYkeN0aR0tzSlRy6XZiufLNc8EYGg1be0
3KROnfzNw+t4jn8vOU31UqPur2zXQBDvUk3XKUEPUuYEbDHX0PmJNWJFfHavyWXUP5Kv1P9vyGi9
gEIXrWXp8VLax1VR57vHE9PoydALmSVXiDFKlZSX6YPP5iy8/JG1dIZtmYTy/eAaT0LA6Almjhfz
QVg+Ma8RlOV4ZWZr3LFD+KO2oRpwfuj4twlOgHecKXP2AH4IHaKx5pEZZt/vdSvO4JZ0eK8nEPju
J81IcTED5Ojx3WoWA8vGmTT3SXl1eNzZg8G9WtzYOWZJYdOcnWHC+ObH6EM4db1NWK6VZR9FeWI1
8sMydKvRBBvSk+s7PoBqwfp6dnmFLu2tHvn7kdTrSGDVRUnwr9wTtDv7OJyK90NzwGAjbdIhm9VF
pfhuS9ZfshDXGu/UQKbW7l97lByUPXmNxHJGgEgH/2eSJeuC47x8T8lbobILQpozgATKBslVZOdC
EsRFA4l2Ie8u7SoKgt3JpMN0UeRis1vnERxI1zBg1+55bu5P1nIyG0c710OIQm3vTSspZY48tjhN
0nxAddJkkjMbAQcqgVAqPhUq96j79WBumAY9JnXP2Ez4QUYzhmEhBiq0eRu4UXjhjQLId/PhculY
fds4g5rb6B3Yl5z05mX7keR4rVhYlewQ+7cx5TPJDoE3QyrPQRQmu7H7VJrmcpz/YXFJeI6nPjxK
Axv4O3RA/1g6HVGrLvpIG5s2p9vtVIvND2tflohyxJBIjykHJd+/pVo8IIWb4vN4oDjyCfE0Qctc
3JBJVBI81ey+ed/IhcqN1W0ovexPrnW23DePuojxLRp6OvongWd9fGaUHvYDBhwZu1YMcPWDEP+a
jDDbT/tJxG6PbfPAvFNjQ6De5fOQeI6A+Wp4H2TYKpOAHIDtIIjlU0Kzj93xe6inrHS5tLebMRL5
5cSwPl3G5zB7c8SONM3tixqFoIkjQGWDHy1t8q0Y+wUW8B6jYKpmGwBgYNRIuW++PlDlJzUz9r2S
YmXdD5B6ALXgT0MmMiEkm7ez95Jx+LT4hgP0ZcLJ4ItemBsmlQa+ifI+v9rEXFVQ/ZkdACdLnh2D
qwifx2NejUY4MRxbIu5xYJ57EZRHhdImRQEDAu/yzdaj4zNXxtW/BsrasrEkhOT5YcAA+5aX9eEL
dSIvMB/S4+b+aBvcuxhf+blxGIqayHkpQixymuCGwVgEGlU5nu+FMmAdngkQhZfUJS6yMnO3CgtT
LbOlkItkElbYDvf+oMnXG3Un9Zo0d22282Q2ubibZ0Zw6zkmmOLkuXa+uVoNOaguAXqw+PIRc8E3
Js+PDzvJ05PRbiWE5ttwVYzNH/R+EvGsyFosNvaQM0LmLNYA0W5AkPC7vxHXPRVrme3WPbCfcQpX
BMocnzRJ2ELc4mjUC2/oe3g/Txqs1lk/XuN87fUbXu768LuhB37ClSuZg7uWceKfXPxYPvzvRScD
6QdFeiX8wK7DuYfvSlDPYGmQcaPV1w0gwDaEFgm4t1hJmsPfcHSIeKyk6+dU4ACWmAG/JQ3e+3af
kEPSzYbolBNJ/m1FukYz0BK5dJJDu/HqlZrpp8TJFShPXUD8Kti1W6VYKPZvApMIt72lbnPyv/Cx
BDIBW4ftxjmELN7yABF9AfETMANc/cTs90JAwuCTtJfM1GNz3XZHospGe8a9zFCpJkCejLjSZCNo
BtCc0olahW/wioSgBfoXOIXtAtBHJUm4NoqeremNO/r17lv9/IpD/jyDzd/CJi/aet7GxWyRdlhI
XPst9V6wQHsGuAStgX7kDwmnGRgIkC3Mq4WUbdNzs0tuBNFsNPykaN0hhjYzGSrasfP4VrLh9k9P
ZPBNeWz/v76HnU4nN65RkCTUYEBHEG36aYvpvn5IczvHrkrznyMcqFYDaLQ8QVRgdErUXiRRe3lQ
RnxqAZUgeNssrlnebAW9xfEX2kkOHXfWJ87QAiYPLDBLjGw+j3iZVJyRpNqdJffRY516MGTy4p0/
f0jbw2opWC5VPz8fB0QsALAcZEyY14XeW2r2CNJ89UsZyR8TmpuS/1KUH+iPnCg1FbXpwLygWBJ8
MqrnJZf5q0q5DvNp2Yfgn1uAnEkL0sjdysBSrfc4uGS9wy91lG3CKs/4wExB2n6jOJCKnvPwFeH4
R71IKCibRpAvX8C76JWo5mYlxgXFkgiVEFlOgcKWTYRABrEr3tQEN7MbYZDPGhFyeWb1N+37Row3
nkwbI17IeKsB+R42WHQXQwknvEbCTtV7ffNAJCULfmT+5RTpxFmj9d0oBRzevNqwZDP6S0zLrMaW
TFzKxxlVbi3251z9evN0tGfA0aJgKRoTMSN6SYp64b80CRW4hJF1gO/KebHA8nukvDDrkao9c0wz
GiFqWEjePmLF1isEF1W8Yw5BCwZDvwM4rtpgXvuGAqChlRfFAbJx6v6vmEQ/2LJqxXOQUcAe8c2t
dI1ZuxTru9CSVouuI5oHYtUepYvRMO2r+parHq7Wd9+6/XoMHzVe2XtmemNT1b30JIPYv4DdsygV
x8vTw4QuMCcjdoESVuNRHCc58/jVf7fUc3wlQa/gXclSy2ml9GUucpONRNdnPEwsXZmMkrQnGOaa
nQIu7xYwWIqF7iNWw2Y9e42JUpLHSb6J8VD/pVy+KfqfZrEqFnazGEO9Q9eomm5uHXxgx88QRmA5
9WfJPnK4YyQcmeUdHK53ILO9SCS56/tAN2ZfwnFDCCsVR82SSPhX0SVfhPrA9Z0KrDtr+XMyRMUN
IGFRECq9fRwDzqa/yBVLNJiLSFMtBfY1sVplupkleWap6C2xrtUs8yBWq5O0CG2pDClqPB9ltEYc
j/GiObkxf8H3hoeUSXbJXA1T981tHn6yOW7DJYxaZWSQ4yv7tsHl47NlSqVzA2EQM/AkMZaIPh4O
svdfqxkDGAcMTQC5dgVEzKepzb7T5J1LBBt2ui18LpTpPYRHIBcpAbLINBUprLXPw10nbTOsm5fA
oHnMHR84yBTRuToadOHE/QxK3FTjyvZEbhI4T/4LBeHPcwHqaUuha1/vvGvl5bpKU+o3LS815gAk
jz/kxfvfz6XWtIj9AcW3osnHPpdHGcOAdcnynSTmFCqb/JEAwZcSe/o22aXNjWkvltz+fV1vmvaI
tCy9Twq9lsLwXxvhzusKWnOD6iAlA3ODDyu4LjQ8O39Y4HtPHkgSga950x/n0WYnxm4KbrdmfiqR
TTvfqvkQXbnj5tZ8mzhRAZV2LgM6v2qwtxYHvzUmM4CX1k0bPPfmbP+bxyQSRPa1j1kNyoIT+PyT
YqTTca8VfE1RozIXnypBEmqUWyQHjy0G3XvD6hAHiyHRQOyV8fLri8Eh6WFvv5A3Ze+IDAZt88/U
UoFzf5PtmttoOEvh1awFuugsFSMgm1EaIc38Bqy+hlIwh5MbaszkWpFZmhdHUOouOt7PRrMGP6m1
BAfrC9gFSqQScWv+Mee/L4rVkVuRgTObGWxM3GO7jVjykfjv399yoxHO1E90JJAeb9asqImNdyzg
KVklZIqQ5lB1aeB1W2kEjEPscCvjoMlQwS1cgiytYJBYz7ufqQhh1EYighfE3n5zR2yz+b5udbej
H9MXH800kDNeUPu1W+vOLD0BUh7IWZ9abt3VRObR87ccube7mysdn+yo4rQjo/Ho21NguSIsLMrW
E/0fmQnGdcjZolBkIbAIL8/Y9k7bH4uw3JgvI7vO/sBxmoAd85M0/DvXrwXlmGBJJ4R+1mvcndGu
qH9BZx9H8yDut3N/H0ecki9Tg2n2pzjJUVKxfzyPicy+9+S6cK38MdjwT7g+WoOhZcVK1QkzQVZq
KfD5/4jJncrCnA2/w8Xx6Qp2kfpeFmuFx7FdjKbQ3Qiu9eZDW/sBv6sxqbKJs4PSDbglPmziZXta
KPhz99z7ILQ1bymcBPSDAN2sPgBp4DIF8jSrzO5/fcEbFC9yNZ7PiKYh1Mnb1KuaaMhuQrUsjIfj
2ZweSW6Z/e0st5YOVBYmh3wZwjji+iOWso+/FJUvMBUhMFR2M788EOVAk6x6SQbl5oroYGGCk+F3
rhcdKe4kZ+Q5yiOFHIO6f0psVDgBuNdCeh9jD5VW/Tnt0N4Izvlr5EhFSFyQSASBfhx9R3kFZM4H
Xf2ChE4N9OcwuHqb0cQaV3Qv9KrKzvtGCmWZtYVMye/DMSozfzu7pQ6Cbl9zZtIhALDGWhuOsu8q
PAsgUKBfreq7XFn/5gFQzM4wF4ajQehkfZmRdtps4Muw3Cd3tcnAcq+INiDSaM8UVWzW05slblDK
+q1REI32RSJMAyCzz5YRi0oL1+XpkF0EbKttit5QkZNenQTAckag0LImeGpbLJQhWkwJodZUea9z
I/w/CVnvdXvpwzDdqdebx9w+J5xxSG8BQrJXBw29u5NvYZR8icLUGd82Rd79q1C1KlPwo2tyHNHY
X4HBZj+BalbHqHbpXSg3lIypr7GFlgwpufgRskCxroEs7sI5qQfSm0Xp7Q77DGobcJxdapd/ys+o
THDqbQFhouoYa/zZkfpICSYdljMOdYKPH+im3Ny3es4QCH7JEkwi/0gH0ZzwL+JidLl5v7VqXuVK
Sw63tyfO4wdk99rbXKDNqr3Ths2mbptvwNzTo27TYxOL0w1Fv5M7HCspSlBzDFOWhHXRXV0L4IL6
fpBXT9SetmBqd3avvZhdZfA0XdeLmG++DQkk4qSScY35vwXAkC6OePd0ZHkCV+SfP7vUykHl88dS
ifO2cUjr4cNOVHf+IIKUGThftkXxTIzwKV2g+huKxUsIPgSc19hA6GU7tQNZ8nNLyA6rGdllTku0
J8VbUzaExmIl7KpLAT7jAkKubRTno7pXFWrtRJuCgLpcEc6WgCEN97G6qwYdQqs+YyvUiYrTfKKg
FtvtYagt5vB53rGxdpufppCZFWfhwiZ3COKWclM+vKqhBhLJSgMufE8Cai8xTu/AXbo71yp3eYYc
7HbRqCenVnnrb03XbIHNjia8Ioy1PRxe337A483G0dG37QlCS4Rn8vHxMbUQLwVDYWuXe1frEtpG
jEL+8aSDk4L/fUiGMYDwGxIEZs/m3ciAj9JbFUAOuFfTz/bkxYnacQ9qhXIv6rjq8PhFWsRQ94Ye
7jtc4Ncy81yOXBQyhT/KSUZCNY3XeN6wvhbvtFnL9ojDQQ+rAnWD969i7qd2pT1z2yTI89D0vOS0
WEjpLtAwbLYucGPYuuCzGqwg8yp65bltyRy0WYpPu3Cz6Br2BZokFCD5IzC1Zm8EhX/aECgjHXVr
gxS8hbgHV8MMHpfR02AS74z6aqaMpEJbXMGjC1iB719NDUwfSCPscUmqCgt8F8aLjOJmwpKZ1U1h
V0TvEGOLNwItNPQt37fBYL1bXr8dkryQNU+UNYuu7Kjn27BozQMG89+zoSMYl0uFBtORlEF105Yf
2jtQvLXyhSk/iEF1HPLqJ/XYA89UHiXv9UYdpMcLZnkKOLN71CmE+R5M+s0XhBsewP+YD6qVKJC7
DSmC2EB8/geSstfZF+unoPbCC14JI83gwBFM1EUOYYsPuJZLdGvq3NUN+JY0hcJnULtpv55MoIZv
JAh/8k/Fwr/cdpTBZpuGuy3lDzPNYFZZi8hXXn1Z7CMoRmUENxYzxwrLM2FPxuCIBE6QIqVkVco4
fISqVV/tSAC7okcPfvtdV0uZ87yKvo3FLmbajSlXTw5gNbRRpahAmSGDx66fRw4/D9lDNnN63Gn2
MvhKLdb8BMPYLcaKb13C8qR6sdz8KqKiBgmBxRV4A00BoYX+heTMlPrRBU397l9XIkFxyHiUc2nS
yzDUQT14M+HKJibaiEkVc5tPGOwc80SX9DMwdzNtYgbnUxlNYktSZA88v0OabvmcD6nMtqTRXX5/
7ai6cAmBNel/pUcEFY3McY5TJMdXMHJsMrMpznMO1sEEbpdKRA5PQJk6mGG+YQHMxJjiIXMwxIHw
U56mNv+sKHk4pzVOLQD2hWBBQBPUcw0OSmUysNe0Z4WeRtrwZAMunu3PvzYLAds8TLOjMh2K5r9z
htwfG5kSHo1qsJuRHpzmB4YiSuHC5n2/b9tTDdqa3GsSaNlLLT0UW1fDTW1jMILt+z9xWGt1S/kq
CC0oJwbzx+6SSSVlLnsw1RV1UIT5OCQ0GE9uxgKisX8PltoFIUMbxvPFrPVfvMvoaTfIjt0OPHWK
0TqXOvxisBYPavmIidbCgTYR+RRrCiG51aadbjPaYrfUlmkF5UMTrsZWTCrmwq530k32uUmgBTp4
wS/VN7GFdHpZghlcZkbBMOck+KlEE+dwkjUcUNqJv/C6a0ppeuSu/8QvE211Q4JrdwkvllXTjflz
HJiFcskcRsXbMZ/9CrFBB8py5az3uBWAOqxuChT5OnArHd5OXWsYIVBBo1pePzAlIrSVN4GgDEn2
tu89blxKaRgcAAcCuweLQXDPbS6ELQkH3QXkZTtnYa1j573qSeg/KAS9/b17Zpkf8giP044OSE2p
TGl95sqOs/1pOXHz6O9b9AGu8WMAF+HvCK/NMRqqMeK6GOHvGSOnckPlnGZvVL25oxs2qkcNPTRM
EqUPoTmdPVLfpUwnDsJ8J/l8ZCmIhSYjQn8cagatKkoVNCsgJKaFBDphOtmPXq/YDYX4bGVbmolm
XdGoebEJRKbW5J+W1rrE/J/d5SnVGq5XLuGIsZooF71yFoYcd3jFwWHWChMAp2oSDVq8TyjBWeST
7tZRS93eNHiyezfPrwMSiZbD+Dj1B6m43fPCjPWyPzB7mb+RHI8O5Y/pUmnlDdolMi0a6k1/tfp2
jenMK+VuCVmFBvaNv4ouAH/vZfhrn31jyvLnn3CEdqSUlxvMGFpsjckxUMQxLihnGhcWLAulU2bs
qgjX8XQQUtNW4DZf/EqjVjA0mWcz3TKSNDa4KN869pZnqHZv6dP6iKZRSOlZ7nMIaRM3cqStVHfA
644I+/4RdYiINShaD6mw29fa3fe/FB9OLR7oaFiW8HHpHrcMjVRaN6PDJyV5gAV4GVBBhAlryUWq
XkVnz/epLs/2gFeXsDO8Q9xIeoHyVaAPZ7ycxZnEBXpw0gUkkHrtIZlKCLKPgaSGmfO11gssH/G3
BiXL/ZbvUwr0J8cbE3h1OppSWgKWYVru/0Q83d+X2gDnEJAwj2bAc6/YmsT+8WnoSf1sK51KI0hw
0wzrz54py7ZIpD5kAO8q9N+HN5zauBzf5DXqwb7dJxxPsvxAjkF5SSmU9CZgvOsd+onPL7uwbzeU
JzFq/gGFcGblHDPjmxB8ukHDDJxD9zO8cp0kj9rAGMLxCOeRpY6e29VCCCGPrOgmLFnoqwHfW0bx
gQpvy9frBr3728GdZ7x6qKrtlSKctidXE6YdA93zCVPYPuP5fr92lerRh+/7fnoDY5TImTcNoJ5s
TjPBmQqy8GZPEGMKBnv4KJpZplPW24bRvII3znRiFlDQPk56gRFkpVVm5AdAzJOcso40DxVixma7
EWGSsso3+JPfp+yR+XmT7Hk++TzMUgJQZEGqi3FygY6m6efDUR7dGj6Fbzd9HD8oNaWjiYizXy+w
95sfpo62j3VFz1vkcDc/NPTxS9iWnRpRAVEJFtSer8T0+sXuASyNUqcH27g19vdKKaXSRcd+2Vpj
F5AdTV8AC7Jsv/6VuzFfNj3nYRSmTyAtGSAImScCotDF4pTHYw+Y8MByVlA5innf5+cjZj6LvjuC
ynwcgOtVLS8GEXifDsKT3gjZdWCsNQXvORniF26kR+SmiJ24HkxCAZXhtpTZi8zxz+/2/IrIKr+h
EtCcYuxbGhW6B4ejBsNbrkG4z20e6tgyQdbvjOz+HsfuRDCZikAQR6/m/Wt1yw4sqHec9dtW8vpR
cvWRuwOj/Txu3whLRXCdSuW/ocqDuON/2j8Eo3LNm4F6PHYbj+uBkVpPvsOOzKv66abiIbnGOtrd
uqHriQ21ClSyD5OzPplUsGw/rT/1jOHfXQfkz/8NbJBXdFZ7JBVWqG6tU6NMSgQhVcNovmLKYbV8
idLyU456O/au9knB5l8eDrMlNow7JhDYCOgjvOEzsLLzTsFgdtlDJAfjDHSGYvtGaVeOvlOwLfdl
ib6DhqUdzETQDk0Rn4Wu2MvPVgZVxOj4VSrmXfvLlUVd9o/tyuBe2D7cPi57uJrscSKCw8J1UkaU
lK8PonFJ9TdBKvBC033TxDrlorYZ7NmMB7fNThx1bI6kLRkHPhkNv0AtVDlIeIk2ELwt9bYHUU2u
u1NxSTCE1N6SySYDbJhxZjaGOxRz807cif/RX+xqlLQaPzMFNXes1REtaFnkvUGDkX2dWl4woY2B
ALZVvMehAe1odSgrAVcIjhzNHVq/I+7sOINZwpgojJmRXegaPMiZaNPxmnzzUL3K93MJ1400/xuK
F6p7PFMjXqoDoFnKtm8lyEovJGkEmv0stJDbj5dNPEKc2hxvhhD+kKlY9VcJYRsTKvdXHRmnmgUM
IqLyUrWXjcqZrRUM4iya9K5UGjESyoTDpL2uG53F73o7OoJ8Dbcj4WsqtRO/2gzxvWN2rNU9OZip
K36fzA3kFiwwU8E6NQ+7VvNsJ8SkNXxuwU/jT04kxgXz5fcSWpPExyy8Z8Npx8MERSQIxuxLUd6w
0HDERFc3pJ+Slrd/jiG9WUoW0GTfXa59ndjOtoQXw4AsR+81WAZPquICtd3B9+kJlGZHDfBKkdTc
xG0jyUcHeb5Bp/TqeRZpQwjZ4FnWFGPwYx0Dyw47rZr0Tom5+mdHEp7sMx3cf5wP48ftywIZ0uDZ
bvbHcxddlHP/OolZeErCWP2ZHYdqIvAy9T//QEQ5JCSrlcm3mrORZZyBz4YDN5EQ6l2Z60OKkf28
648K2up9+HgKqXZxA4+d9xv6Rn6UgQyAXKFc7tMBpNE/YkJg9fYcKQIyyWFthqmm5/c+hDaSnkF0
lls+4RTjenHh5soEGb+5FPve2mnGgaxq6/i6j8dxKTFptqLyZ9pITVtgvQn6btXp1IEl+KLfs7d1
Z4YO55pXVnYdeFoANfPETyZBYGLtDaM5Xegh5uruUfP0fwnuPyJgA5+YGDlHCxQn2ftNcRWDyZm9
clG6dZHvI2ToTmhbZLljQTg1L8TlfHPnfGUuVSi4SXny2FBfsH+n1XwlTB/MNGZyPNEdVdhF/GCa
hralvDVcMNx89JdvsRM+R7nSKiRWIUGnz9HUJYGQM1DeYyx+8yHVFQzz23H0wb4HLM60AzJLqiiy
tCiCviPUpkI+pF+zVubCtcp9k1Jyv+Kbd+b+1GCZEbKmu5COyDPrtqD6UNvBFmxXT6emm64U2hMz
F2LPO/6iE8SNjnmjAfVWPfPA66TypSH/zqPPMrJc3VTvkXm4YCHrDrJAtkjMhE9YHTd/dCM3Jeul
FevgLj8nDyht+Wn8jfBALdZuT4OFJ7rFn8MD7/zjOQS8DUUWOZEJD1RJlPav0DEy9xljMEWbieaz
4tQwqaLRRaIXa3BVfJaCtl2BuxRJpNpbFUSgZG1xgvvL/hMeD1snn8Ww5Mh34hK4YHd20Qb9h0YT
0y0dhq2N/knZlO5mhfIcs1fzmcOuWzUTnz8E5G9ouR1S86Yp0IgTjCLXqlYLlYF43Q8wkVhsM0Qe
k1BQyZiPJGBTz1DgWXvp8oUYH+D6D4K4ulvZUKg2veNX6K9aeI/LYvlXwIy63wRiW6CgOjWlKDDr
3sioTQRCKl+VC5oq/fHir7j2NjK/d/n1IZlcRCdE3N77KRUmcxWqLqLKp6Pfh4FpcFHYeDMzeghy
KhLSGbkp10/6g8I6H8VnKu9TU66AYr4J4TV1xzvWo0cDWRLQZI3tyxGX4ZiB7bUhOrhtDMZyKhTA
rl3lnuGJHQjybqFc98YMdGqomgafXOfrtPc/v+xodnAUrSVQmleuZmj69GJUsjTJO5/qNJmIitV+
WWA2t61Qkfuar7MesW0HdlnIFhBVL47lENzu7vpJuJVzGg/oVVPJcBGScOE35pDkMqXMG9arbDTP
WNM8nxeAsqSHE3nqNtCYL0D0dH6N2qkHkMv/1l8lO/8LLPPll1ncHW/UHgeiLUfZNz52abkpzEap
p2Db+UE3xdvKKGAGM/cjoBvjizmOX9dWSuQvpWVD3qzF1YOR39rFKDyA8UDkNjAn/FGdIZUTDO5f
fBA5F2h1U6DXjTYRpW0PkV+MZ461GfwVGWWFTsVMg1ESQk8+2VwTjVLrrufRSVYMoowiQjNKP5wv
z3quDvv8iAbumJbPI1vPjEOE2ozKBNqFnuu6I+4bl/8lC/Ze77zvEZfP+KePcB/Lh+xVbKpMJFWq
0Fvk7XEuZoNV46WaB2IWdHZx1tqlnSx7e/NThQg6X/p9C0VhunASYO1sexNzfaz1rzo2GUdpGE7z
RfBbUvbcsXY5olgNNMTpXg88veZNLr9ityBbvvcThH6tjhBWVdRJuEXhLyimyAQdwpCFZt1TaWEp
MVdCC3pW7C5totIVmQmLHBhJj+KnrQhdjUQAaE/ygBWN5yd1NA8ZiPRYbi9J/mRrSONDyzEscnWH
dTPvSW6oN5fAknPeHlX4hiRpEZd8h0FatHBwD5PHJM2Kkd8moHx+/Kl4xf4Zw4CPdHOoLExsYfBc
OIIj6ERpxej/PAQHbTgwq/2149xzh3UUQjXWFjCaEhr+3taT9scSk299myt5hEOg082kGylx2Ati
XM45KMP6Kxfe9CbrukmvyAtnWT/PDwdEGp8CoCuqf5MCHyNP+1HMw2GLxPMPsZ8kWoOtSoLPCHjI
m+GXj0harSEmTiKN54ySutJSkWiARuqKKPLhsUhjI+cY0CsUsHO1hK1Twvv/Amj4ok6RZ3dYRwxl
o09MPJoKFWSWA2SzMGBk0HCaWFXRwvEVjoegihgnpFwOzw66NSfP+wsiD566Puw3JM3cLJadrGov
EPKmk4/I3fpyAOcERRdVZpcuje1P3jqwoNEjw3a8NdJzEPEaASAJV5vfKWMT7DRaZh8gVvomaR3e
iSHLFigtkBd+9avHyCRteJYsAMc6xSBbIenyZ7Pi5AA9lFud9d95TZWt/LR2m7fPoZSOOAP8wnUl
Yt6Ekgv1xppm5PWsA50JNvUZNc6F72HzMW2fxGvpdzqWZ1pQ8tVcA9xk/teTc+dHW8ZkE1zM9azh
Uljv4HJWGZmWGqz9C4/FGVch+861XZ7Djxx+aiJgtw39Bpw3/WYr15SbbTuEH/F+KIEyeNW67MMK
jHWmRn/tEoceVZbiG9x8h80P00Ty4Auckcet5cfwF8Q7cOlmeSVlYVuTSfsiAUutWJebtuzrIGiu
fAYpyM4eXL9zZWuRHCK5gYGY+6e2Hw39Vem2iIwP4ZD9sjRcFnEpl/UpIPEYhIeC2A60dz66D5Ld
TynOYA70HSF3rtj9ECkoLCGBOlZEEf9iMWC7CfgpbvJqbNx6ZlJz22xR8PKuKqAGOBvVOtzS90nL
lZIweE0twoeGOxNvQvySGjofJFEqcY4u2uawPd1lmqjGKpRGldj0l8DPdKLM7Nbs7X9nTz/d8nir
j6NJalKXTRNjLSJvAK0GlhkeITihCArUGI5314bkVI3hab472lcm9n7iGvBOBEZBjXgw+meAG4DF
IPpaAc8DE0569iFzC8ld0k1MWkwIQJhd21RfCoNAiER+C7fs6RYmSwU/df/XwDSLWbgi2nuxbwpk
xdjZtXifqv4m26pIHAJx2B08mPt0SpcO/XkoV44S0SdCyQhZu6ZYBoReHH7UWdqBO+GZl+iqBTsw
l+SGYdzZGY3PVOIB9dzqE6welHguyUGtsFXgmmwpbEUZLu9d5wkWyBqPSFzFw2Wubmb0Piwz26ZU
OoOfsJ9bq5xbtqXvYaxl24ISYugy/UhxRpKI1IVr1LctQQFHWAi9kNwr5i7nt8n3BlqQ/JZcx+dH
mD7qDD9MW8WjKqf7UnWrK6zp4gStyKaw6QB9RAkxgwx66vienEnUEWHfcDn7iB6PJG3GtilHAy50
LPIqm3+C6NyJtM37+31u4FhZ/3JRYgsjvQ+FdVHrTKidWNF6KMzFnAaI3AHYQjE/LjofhWrBU97f
puCgxLzAuHbK0hd7CNtTQrnw4Xh50cCxiNK6+IpT8rX4ubhGFyHZJONVwzeUI2EMX4HOj8SosC57
+jvAo3DW8dx3i7iivpjarG+f3eEAXjKyEdXrVYeBr+FReMyt/zml+YAPXub0lDuGFvhGC4EXg5i6
Im5+IdCK1M58AWFmiEGFaTjFwjrG6zlJ/7by5WNiVOW603OWONDqT7GjJbwg8hZ2GlKlOD2ZfxRt
hR/yv8aZWViY2xjGGfUQdymuwwLDgMX7lxhbj/G7fN9/h2S2EWgIidNnJcKtgHrSJDDnS9nhdHZv
KPydyXdc5C/ITIhOjvMvxJ7NzuGnhQnuK/xbPULZ+eC4FSYyk0BZxaaFdQk3TOq6K9RO3sTKCkid
KEEb8bV4XKFAyL9lOorZ+O7Wcr1oGKZ4nI5PD9aRVqEeREyr6Liikhr//PShyta9X4HlygLvvasx
jJgplR2nPFXB89TEZi0SWEqAOODALfoPGd2ZIxpIC1YArJJF41xhzOLOT29XqA8feNijvVzufbEJ
NUjdgW2Ijd9FxY3VdEqo5AmQdLYA+9WTlcM4MDuUKFn/Q3R67GagYKMb8fHavDNy7Gkc++qRQcw0
0PIFTs3LFhdi6GSr9zE3vbC9Omb6d0Eq1k3Vr4hKZC2MNPlrODniVDlCg+Ub8ctJZB2ICYeBICdn
ChLpizYw4B6YuaTgHie01g8XzMh3ruPv6PLQDjmOVoYUB3JHp+O6hnwJb5wFT0J7sUD1qLlOWr4e
Ap30sQBTzhmdYaMdn6J7PMMkwd9lXPtLVBx2rNM18VE1jpQ2FKJzVFItwgVi35f+tW9bOENWgA7C
vnF/Z7YQrSD/E0eQV/W8A3pML4kKNDZU52yuo1u4MZShv3ug9T/FGnvVc7qq8hSg+CHM6VqxZtDN
mLp4V4jrdcLAjVLsskYGVL5iN/sNWrzEX99/5RITwWhItU0d3Qbb418h3/+AYW24PCKdYi0P9wA7
b4KnWGDSZ7gghIKaJH7ih7xC3xnt1tjXQ8SvH6Fy34uv7GuVAGligTtd27ewLFuvYkYWUbX71SbS
FW7+4E9jbKjVUUYlL2Om0pzKFlh2SSwpsDSgFGOp/n3Pe+l3bM9Qz5VqkVHMetgIUM2qPieAo+eT
84WryS9NFz9j2T1dJRZn9s62UOBy06P/oSoF0Mn8OnYGtlXFS2N1b14BGHKvDp8Ao6YhgVEJvfPK
OIchwjbYMmXlhM6UxbtIS9QIH4OJBhfig1KeH8vmCR5s58lLIwuVuJYYFCZqZpd+wYsUtmbLAgyF
GgweTFhgjFccRazAx4/kcwVfkk++V/VqLDQ6IS6PppAaQkEZOCz/0Gct4221rd1+4xs970N61ZJC
t+dwnIQK+pxryxTQFRcKg4vtYy6puquIKehKEj8Cn7mjwTYBnbmunR1eiuqG8idMS3xTiyasL3ov
3n3ju3RYI9wobtJ8nhk0f7aoU9UKwZZbNH3gSedmXPN2pzTPhMR/Y5DKbUDNMe5XrTklUYRJgli/
LZLeTC9/BvvWXE38h7lDDL+ij3YL9HZnD5PTjPd6Iev9SnxXgp8WADpZcXTcXbtOl9WcmnLh2Xoo
9JDyJ43pSczBYzjMoTpgU/L4xWx18jGR965lV2FPIswr/opaE6EJr9rBXIzMlrbpKXwfuB2rxEEF
LYH8RniJEDwVVCI9Fvp0Py/7DjQlqDi9l6Pqugj5yffZTTVM254f2pupGE3KaiMRoym489jH/n2+
qKcNMag8v9pviITf6/4HLhZ1YyBALxKH+4Kjl+undGkRT8S8nlEinyFg7AQL7HzGT0M0gygxm8iG
wWhNo6OfDEcfGKC4l+ydH9cB6waYK8Tp14mMN5kcqXkYawRz8u3WB1oEcyu7oO24QtfZfY5Vm/lI
EoQkAaaOPO8tK51MOBHZZlI0ohTCMZr3rxyYqHVQYeWTWbo13Nr8/+FM9B/jaw3vyhNXjelnvmgW
qNT21i650SZiIp0gcExKZ9aF89x7SspqNfldfmVdMyUMs/PyZG30z2DChulA5Smr7mGbhI7u5eeQ
16j940UHmZXGqgCVZAMZitci27gwMU+zUzG5W1L52hrdzOltVL0EO+KI6GBr5cuWtznZswNaZmbB
6iocoakVz+YvtlBkDZAejtcYukP3vddKuvl4iOFKqUsULtvTV+vw1qA3nxew9cjpCPzUllcjV0no
DzRe5tDj2KEMIM4rKXvgvphqwcA3ASoVl/SVrv/gH1qu7uRkwQS4js+yzTOv5thciCMf5C49y9y8
5jzKXlywuNFXo5ToO4dPyYfPA2SNqn54uSBsVhqPuBsanPhoQx32sjiU5W1xoZPj5tzAjS0z2zAO
1qGbmmI5opZY8kN/P21bOKms7lcQq9Y49pnns2QBa3/z6EIbZN8mjJgpkILYD8zMxvuwK74qCaqG
Vf7BpNZ/btRqlkU4qcENY2CcQTR+oSx4ErJp7mON8yameuuPiETC3yu+QuIxsHweIQw2/wzu4Pwx
lWOS0A5l2V8uYfgwajzIThBryHcc76QBFR4T0jevecO9zo66rm7TCN/7DLxjm5TenP5rrr5iXq3Y
1ghZYugH58hUOxBHFrTcs9jOGwx+aDI1V2tx6f1snLT3WwbkHL45DJ18dTopa3KDa58RF6rmToS9
EoZ87aq08jNzWulqbBwzyB9J5cIJYPn3P7FIQb2/0hyHNklPrbcIIzpatp022w2MAKlMYKFnLCcA
pFOUi1X9vvOtvGa9APZkR2SWbuzDc5sUfcSlzurddgT9xTk8dH9/eWZi0QJI/MmMUiKCQqS7LufQ
nmVSoj2jnMA9QP4EPCvkO3RsK+sdf3u/aqw4y9DtBolZRXQO+svpGDwlM+iLG1IQicJy2rEMX8zk
tPbcGuXsV5GaSRAmDNzcUQGYuppmHwIbWNbzdu5veOiipqp+3mJ9AX+fllXgVJ40Dj50oVrqKd30
1hWU/hivUb7twZFbrl73e+LB2o5rAqqzLJGppxwt8RY4F87Eu7siCd6unmUBJrDfW/zWLv4ZhDmd
cd4wfNnMAA0qzfCeW1zLF3mom17bNOOxATCa30GAoSFOYKNlpDpupCPpG8+cwJGBOZR1gO32aCU0
FiaIy1rEPUAz1ntfGO9guqplegbmNQoEZTX7wZIEtWFaI3VikjMoM+d6soIYxTJwMghBEETPOPyk
iHhSpTmL5wPZnroLobgh3VBKaYn/sYwMfnM59DNOjJhC0k5Gql2KjgxugCg8IofqQVkH6Fhhw4qL
gAw2VleddP8LjuFkQcvWrpvfQ/6DGW5QxgQQEeGPIPLQ63y1Ht+9yDyMc5iEDWMM+GZBKWJy1ABI
7Fk2d/9bMiGBa2+4c7V47Ryx+kjhZx3XYCe6Y0mtm0IIEdncJZdfF958bNAODsWotmLqG4WG6sK3
AAPdNO+oCLxQ9UMN4cwpQDv3V0Bw8Q8+VXdPo91YXuMrBge3aiAStkqOFKh8c5qozJEsZAWpgGWu
Cn84NcS9DJyhvAs0V0WeHxucxyGXgFTYYRmjMqBB6ZHqdgxxfZkOGTRw784ZlK2pBlM5+/ftPpJc
mo5AFd2ygvvzPJFwtUTloy6D3nWUmOSKRxRQIJNgCx584O7KDeN43Vd/DkbU8qSWDKsejOzWVpoD
+OTIzxjQwFS9duxPgVZC2GxhZBI3qCut3nH0kfcwU+I5flg63HaGA7DvmsZ1WXZM3+OwLNynnCoK
p84MP2gajBCKmheWE2YiyK+E+TpUksNMh2jqk+9kfnpkgDEFej6C90ppiKccEwKwPN4F64ug6eBH
E9eAhfHqJnA+fx2sInZx5GlV7uBvdA0vm2C0+gDeGFhzR5mzwJnYlRtVSoz9Ag06Oc3s0rExN2qE
zTOve3pH6/2VIQgFldj0GZwnfGQjTSsxYGPVQlE4tAVGooDbN3UhOlvmb+OP7M9lYN8hzeDZTnvS
ADMCMmSseSeD+tjogdT3Qio/Oey/Ss3eH/6VEPiy5ZueE1ngkXobogyGehQoNwZ0wWFQZ8rFTwwD
1noj3t3CTtItwcwe36QtWUiX4fPY6rGzVMLr9lGgXvM1XyTXFJieK3l1NuLsSP1Y0nTxzcZlao/L
Y/BVdvP9mC4aT9Wy3tJOe0fqDT+F+F5Prvj15Di8G1LJQAo+po1XLldvycwk/0HNVvl1bb8TFUw7
FEfwnuBQzx4DOtoY62MwS6KxOAhtGtzc5BbV6n4sdOcspHycjiTmj5DCUhw2wWSbU/RnbdP7+3V4
cTdp76cNV48kRo3cdPqtLHAMSkb2PPb5yABraTX4Ej35XGuR2xJAx+mL9E+yQY1Cdi62/zLKKT2G
GaafNabqn4DZyJy7ur90cEzha6KYOJaAQSiVh1XDzhuearIWxIgxiGHeXimoPSLB/qePJFUz6jzJ
VwcH7ULkzeWxpMkbFrDLdEsCZ0EGLd1sea+EEJVB+ry/8/ARWTqjb3aAVUyZiRrUNQgjkVoaLtRi
m1R7cmrIUEoW5WWNEnIM8qFebriJh52a/y73tmMVHicuflQqWnLhoHqNi8PeNsyFHSEm6jUaMH1I
3UgjBP9CGHHZAd0ZoIGOP+0d7ZTN38sNh5cdG9pLvynqS9pDivnL4JYicv1Lgw3methaF2UAANwn
N8BRO2wK5j12STxSQRKOgQu8iBSOWy90vtiPA0vxTGiBwb9vAGSdxX8x3hlqT+tWupf2RXne/Bb/
oVYBRtiolRSHLd1hff1VGu0YdI0zS0yGOL4ToHutlrL4X5Et+3HZxTBgLYo/G1zgfQxm/CnDBZJI
dvXka4ge2xk1d7p/ZTiqYhQG+LDSJQuVFastsRoMItNCaOK1y0uFfC7IxU4c+Ef1mw/2YRMY3DG2
LiTWmBE3oHMAJ+1tRaZ+EVOifOp+TO6LGWgaAcQbRscbO/hlipJ+fyEf30lhaJS8T9Ybr6/1rZli
mIp2ZLUwlDbRuijd9L8p8ZGGm6S37BLkTKmb5QL+v3CR8c51QjdlY6q86jJ91BVzzu6//CiObJ5K
Yrp8ykYdm6na4AxQRI9Ym1c3nw76t6+ugaebawFxFbA7zCubWvHtUezd23hAg+NgOe3RoGgqf2c4
ReNquQcuWf+vUSbRnisdaaHKNNLzrkyC4t3hPhpw3YRILVuY+m2RzIg9WH7eMQKGIpzaKgSj/BRF
pxLfGVrj7zHDmZRwkEa9IuM5b+qvNzibZv3LuqlRtJkObovnr7nJ4RSWfSdWwLkXMWAjZyq/6Okx
P6YoYva6dW/R7N2liU72RqCLVSLjcWkO5zWJOCK0Zp59DMGAQh4zgrDzKRtD4Zbqgiza96eFrGHG
QY+ZF5nhIPlsJIhuBf0IA4FWr64hDuLts5a7QgXISSyN880aFH1y5YhIDhYx06+i1n05d8Yk5A3J
dYLdqt8YUcb3kz6P+ES5u4WytwQr5NzzSip0OtwN8h9cjvEFQ6W6zKzSZKt7xB0ozj9t0/W2Ei4B
g3RgKAT/87/0pYgXAD1PCpekHXqdJvNHxSeUXFrQ3jCA88h874Tjx/W0OjMTipqscuGlzFLZwV2I
FC1fbNf06z4zJ2xi2CDlYMqHYiyK0xdS/Q49dhYS2bmyLjpMZ69YYmez2F537g4bsT1SavuuT1l6
YySFdxvaxLsBsFbhloZDqhDEYM4B6Ci6SviKKLnaMFVkw4rEco81aasK6lzez1Nl0nT2ryjLPC3I
e9pOutjLLwgoxYN1fI8lXcHDUzvXuaRMmI/CF9nLyoRcE9eL0n9dL2dU3v7CdcqZKxlBKV9BUbd/
HdF2uv190zWpIsRCU3gXy3SJpu+cLoEvpqpcaS3zOMpLhP6qC0+t+53mF4F/NBtGDH0lp563tr6n
VdE1J08Mek/CqE7r5yQAQ37nuOecNa3o3s/AQlBIZ/FxIedm+yC22AxkG22whi6sfXh7AMpMPdWd
aVmKEBRiHewajB5ri/M38+KOzivWcwQftdlCMO0NYbYwj8KV55hGuThQAT4AqBcStS0O2pSWxA2c
rGQ2Q3mJ+0TeH+A6c4FyEXW7aPpT58XwD0oAqGlnlhXgPznCcPiufF10Ujajmw4eK4IM6DayP5Y6
6dylqhh6OT2HjX/SWMWr/GIOk9j2vGH8NSud2uDodiDuh1YUb/4S31hWGQ6LkvSVvXFnQgSg5wr8
BdihsQq6GBAkplgd9Q8kH45tGdUoGuFhX3TCyzh9tUQ+ySr1CIPRB/z91tXoXJ0BEHsJwKlBV9Sh
aomGRBoEW3ROItH3oEdqfBMybVmrctlaOWj2O4zVWgwzayLmtPIXAs6GYbDiOnnfQrgARWUu7RCV
9KA6ePyqTK96vt4IYceTlKvNS8Afe+gHkQvgaM9677GfKCOXYhVs65JfHhK8vbxagxYM2gY75Yup
hHZSE+Ohb/SnqXmbYOmIq5tUevL9WBLgtMS5isHUpEy9QdVQdXo23YxEZoXN3UAkQRW4Jn7YkSOW
felf5u9mkteTAZjKIitqXdPFLubkylSA86RzK26gD81iQoNowxh82omtC4bohgxVYi9Z7/MtYeA9
O9gV6jFTdYPzIKCSC4thI+tzrccCVY1XZ+/hoC152d2hMaMAn8lnSmTP8GjeLTZyl2how5nREF7Q
/WxlGrVhhHhXJ4ibELi+/WhFDbUYHtgnw9lelo8YyJPQ1FmRLS2KrWEv7duaRbrovnOxDJpY/Hkn
5in6K7J7WBZClxweDeiCpNRWD7QQjuYe4do5AOIwQOz5Emg3fOyyvckOfWxLnKCuy2oCBbvmKm7V
c6wRyw5NX9hrX+63l/pDMt9pkwrDPoCikGKWV7oq9uzcqZB9TxeAvdQuh/vPepmu96jEj6rU9xsM
fbXLabVMWiVHZ6iUZ4HAdb2KLFDMXfpyNYDMU0/Y1RIURjnASMMTXAu1sM8n+6S7qhAi4QMaPsgW
6FmnUWzfI1pcRCaue3UL2TkcXbIIPTD+Uvt6bw6ONIr9Ft46WCm2z+wUnt5e7wu24tFrmwyZjc/e
Y2UShrFYbuFq4oEJBuyT8b5QTVLtwrnqnypI2NFhc7aslP418l3ggZZHxMBI7lBrcWB6CVsQOUcl
SYs4jfTxtaBkFJFpej9hOCov6As64LrJ4Fle4S76EJvIbQorUXT0yXacxS8hqSnPcOtOljlHqBJm
ilKgbFAgfjYcwIZcrSDqapPcQD56NxHaHiJ5YeAiuzAlegvs/+2VOxsdB4Qu8A9PfcO2KZWkS5f8
12gNfMZzE2JCqqxvVQEiHgPfPYlvkWOGhR18zkfVxZKuZn4thC+AUfylIfHVOtPSn0ZFfPxMsaRc
TWXP2to34lkwJS1Ie6VY4qHQYPV4ic1aEU3MXqMWFqQk32BpxWe6qF8Zd3860XMXYbGpnReU8dEo
SKcJBjhiddTscYL0qycTLoMX8FNcl417l7T5MMgLsCBpc4DpzHW0LQfV7T1pVy0mQTHePvIA38g6
c74LoTuManDOJ+xUFyWKo+R/8tBPXJccEkY5oPRkxgNDYdrPY+7PQ91PP2IOAkIML5K/sImyA06P
h7S+bstr/axTdWlF8Zp/P4dP+n2b1RUCqlgj0rRbZfs6ZsrvuI0NhApBTmRTxFN7W97PLCMx/UkB
sHnm7CYBSDAqKH0MByNplGcU/po3+jKdMfhIH6BD4f4Q34a2U7BfE1oYDPgK5SzRbD6HpkCa0QKL
WjIjtlH/RwaWpz29wxDkQ4VBXqIrf5yclk0zdIgbk3MhWRJSqhuj9EqIO36WwRld2CcdzDAsqxjj
Swdj8ZJHa1ZN9opZXGgZSfs2WEMqmSE1HrfmMq5GhzvGGh3TJfryLmBq/jOoExmQXOTa6tmVjRHn
KS1oS+L8p8IGIt2/gsJ8135mV+5XbBghGTC4hHy3DVoyKbnBc5rFlH0lseTTl6Po5PJo0XrWBo7D
DQHl+P2NsW/vc1aqUic48NqVh4Wkyqu+vUodBlDFa3nNFWgnbBS46Pg65svDzdY8hDyQOKGf1pHK
LVFoOLYuYsMDh+C4VvN7nGsYl3xUCiEK+AU/mD7CbSeQ4M0EmvNAH1BtJZIwKg5rS1ORrJj2XTJ4
hnv1Xi0wncoQdrGkXgvcKETXdKdhWE56HM7N5a3gY/lXR48PSkdbrYrMFCse2Z0vflPkp06BZizf
2HZFFfVa1QtaMXI9ah0HFMNH8YAmFm2Yz9HtugZfJkYeuNhb7rLcRj0c8kpkK5/0Ry/2pXj8hGri
Kkre68o6/7IFrPSrOxMOQiLlQcGCBe+Ok25m2R/O+yQJn6y0Rw2gRM+fMWw5Io5Dff0+k3jhmS6Z
o9Zettl22Cshz7bqYGmENOpPSeIQ1ANINbcQ62acHsoVBx+Gyn9ILl8WrfQfFKUg+Udgho7zdWgY
V2tIyH09UgS4M+ouBrSwGGr/Ajg5/D7PqQoSpNJKME/2+7naZ7MBHLFeGoMkuV85piHOzFzudbpp
2sOOcD90WfANbPN1s8s/razqcxlSDx1+INtg/8ColnQPi/lxN7qVt0/H08OVnZkxNJwS93Go4dsS
CjpNBw9HTINFiRd6CzmXvlnKAlKp+h0wAdp8eu/srU6ugxNRligxfLIMpOkmwf+0mfoXCk7X78s9
FPGBacKpfBWhbedhXfUI+A8CCgWpEksIIWK2xnm933KXaMiPnZ4saBslUB2g335HYY9yvs1CpYEp
/U/kCzfuwgRjXg8ZRvUx2V9vvG5ZGPn7inMV7t/rFAmVJ6JUJ31wPDvqtCYsq1EgjaqJKtxfReKx
uEQXq9gLekkHjef0RmD3Chwo9gmJ5yv72FrD1Y32EKcb2xIF2I9oXt9twgI9rBpZBvCVkHpmxlpc
Mih7zlvIJ98Np7LA8e033sRSwkeiBDNGQOTlx98SJgYV779/AdxeEzdRTLTlGIxrNmfZvzK9KHM+
/B2hLsl9ql8TMcsZh46s+RJ/DaiHosFJKbi77yqP85yy/u1lacb7so2WfjsvfxhaVz2P3lwsT25c
6WVNEb5FDQBgEpT4xQ09vD19umKO+fyaX82+l1vMTC/Xbd11nGF08sab0DuqiLt8cGecBgVxX4Q4
5KqDq4B/z1FTT2TZdRya/EXkwqMOj0XKQz7jA2qDQiIb4uYHJ1kytUOCUM2mxXeKKyQ5HmjvzjJF
Ryq39a9GJ4cZ/quUfBkucbRsJjZulh7i6yFco4rhPG+1AIN8HYLGdSqxPMYA7W+se1X0gfeFvXHB
OJqtDz8JEmGCyFHAwH1CAzCXUAA9BgwbK2ERzb4seDJbIPkG1YNwAE6QHKqYBsRliPhWyd/LqPnJ
YxvXxi+LLx30Q5S0cjSwXwaazykCfkGhiaVCr/XnJjFcL7qKjbSR4I4Z+v2+O+TP9uz6giZNc8E8
7unxI28GMIr47E31DxamB/eHv2vsTIBrNISOJsXyGTsp14dcw8XuZiBYGPwkQmTIeF11dtOsb+dk
m2e9y49f3Kq6ISIjzw663N9qXUg0TmOc0cy7LwofRVoz5RmJAPZl1thJdJnkWkp1BpVT+MNotBOF
fgamf39u8P+8nrkReYp5qNWcYA/pbi4YlXJPZqG2fTiHKrPY1CGM+gI8MJoJfiMbmG5RDfbE4Gms
rxIDmai2HlsZ9u18jrvhSxW9d9hK7/JoM/z1uV4OrSRBtTwKD5Kz0W56oHrmKS1VbqKsXPAvsFSx
Tze9AIOApPaWQSSigF9W31hvBv/OOawcBJBgtlFLGgwr2zAV9FE/1p4ZQB0qcF9/eXS/VUcVdgsc
E64fKEtf28QJWpoMvGuFhq1I+03jJDCUFYQS70pIZUEgr2iGWeKPCHH7HUeQP0SpV59JsDt1FaOa
vrsvwgGVYWcwESFmyCXluiLstB0GtmiFe2ggH8XKvTzUJPsk7ump0KuF3Q8tZU5qmzV8gtvGwhvE
MJ1M8JArT981oi3bnQ0ak/CNFQgo7G/tI2NTnxLR1cq2jhWik+dJF/iLYTjyB2g23Hx7dYKtPTik
XjWYt0upYdshpYqykoiuJMBzQYt7v9zR/tr0B6KUQThktIbgN7Dq+Ar8e/skLpzp1/k67XqpznNu
9oqFn7MsIgFvcrhFPTrcT6LpDSG46xOg6c8vBOk2Z6b/2BjQLnMVUEvifaU2Y1iTn8XvKIZGVWdH
7H5P+yQTc9a66SNOmAvbQPgSj3tmGeXx6oZZn34iYESyey0/WxWakFUrSM92/s5autJ40d/B/2EC
OTOGzqEi81RC1jzDUib4gS+h0/Ui2+8FqwGaVAu4heuwO1ZBYmntLKK7WTygWmeo0gfNwifB4aX6
WAyHoa8oYtkhaBBkjLVZTu9zK34SPeIK8MNvNN0Llc7PIOSqOnFrCBS8udwwoeXdQZBSzMovRlP3
zsyK/2zlr0ZgArhkD1aGrP8r2Ix/zrPnHleqLfNVi+8uzz3hoYtImXtAewCzBKfe9CaJAaM+yHsj
B1tYw8FDWINeeUeEK/829xkFdM74DUfA+P94Sprmfk/KiDO890FPFCVByFSsbypp4BZgJ2rJWZXq
LZ5TsY6ujp18oSKfqj7JcswHsREulOCATNEVkDj2jWMQGVdj6W/5YbO7pVPgXxc2fS6iNvA1nV1Z
n316oX8GKLJt+r0MabBZa1XOJ1qLQvUO61PfIu4xA1u76NgXtj1Vl9SskEHsXrx/gglDrzBytluA
nIV/KpZqTfDaDExNa9ci8YvsFow1x1xa1XvX5BS6mCGigO3HcFZSy8FHH8q+nEqsSVfzGvN6exSF
R0e+XeeOLMmP77jbJn9Ayz5nJ4G84wr6cu86pVJSD4u0ek3cqtWhuWIuiaXHxvOxkFgBnGDhDsdf
nDfi4nlqpkzIpvdlqmwvGEO+70Muj1dAlEl3idhbT/ib+nFq1AAqm2n0Ja2JUkb5VigD8I4PMRhl
TqYm+G4ei1zV7h7fKw407g4ztaSJm8Wu+Z2/e4luLBwnZK0WNrjdHzY9BK/ng8PkzFSvuZYcRGJo
srVIxHNuqPxDW3uY+YaYapHj7AwCGpUPnJYPCifBu8gvKDfINl5SNbLUGHa5YaV9k0ylARIHOGfz
4SPADv36HoLkvMnmcZaNXeQwFRb22+pUVdfT8nW30n38TJ6LwKdzTNEC1d7CFQg9CPb+4cLAYb7S
G0VImd7I5+WKpfAAdKfvU6QfPPZYjXKuN8R+pYZKma+K0fi16JNVsOkpaCx8c+hP8L08fSkxEJJy
A9PVa/tsEyjkgWHa+jwjLCkrVPYEsGgLVHOJJbCw2fpdvsYMisLOgYeOIFSFR8+kEO5NmWx8E7bL
VFytnSZB4c0UaLHja7AVvcS80ABAk/xaQMePSBHK5By16kcqZXomSPYBd9WLA8CGCDjGMZIQ3Ct5
Z6USzAref9b10kvVEctcu/hTn1mqZoMJipJ6N1LVOxMUaWgE5VWmwSHESJcmDwou1RZGADYRVuEG
MStyh0NAQnwvLGzdO85A3K3MQR5sIoghVihyM+149CLXvKU8E1kDr6xtglBB4UyHQWqW+1XfBqDv
Rmbc4bhZaqkDrUZN9ojYyCcE0uO5QBPplA/3CEayJLjqpN+9FcCSzEWuXBikRya20TCRGlNAwgX9
c9VbWqEbA8NBrZwRY0ySqi2omoQCiJOOEexbGzj19c+1Ym+BQPH7oFS111CDNWqsYUr4SFeVRW8p
RTEK4QEn9JqpHIJ9EiYcVAr1INlvRzKQE5XLRDYqAtjkJAxd3UnP/Rv9zexwC+OK+SA8tkDuLrnR
/CQ0kFBHJljQi3GrBaBFjQLC63AJvg3Jbha81G0tM5eLAfkwsDj/t/pzNajvrVnguZB6qGmH/wjs
jMZ38VfBeuun8cswGxJ8HvKS6ga3CB6cS9WNPZmDyFDW6UEGb/yq51vJtQcti56/jVK+WArCzjcx
nAJpMKIo7zarIpnlYykJUa8rPVYBXWrRtMfs3vfTuQZZufZACX7VJwa4gAtUDfOiIZT7wY6zEmAl
U81itMfnqHdo73LO13cINBIOf1Q7hQqztVwTCqarrtiAAKVwuAw/8nf65xA110jkRznSEl+Bl4v5
BYyeGxBz8fh6wbbTvkm0p122nUhoxxFlwKQtcHkwgkmTU/dRnTYx4e9gx/rVSIeOoO/FjJmIkaRU
YBjAAuJs9iWjjhnzIVdlxDAPIVrMe9t4/ZU+IpN595DGw5Z9v3iciFN5szcY8KNLIyDwIW6SCMxR
zAt4xItV6Qtd/CYvm4CFqgo2kWKA+CVSo15iDc0FBvwU4U3+Us0xb9LwYWhC3U1gcVJnyXhqu+5n
obROy3x6Enj3dFBeUcDISninWJoys0DALuI9cDc7P94+Ud83CTS+lFsAC+z1bVJxFmTbbynvFizm
S1XrHmb8Zf8UsGgWlb59/6Ij5V/pPbJy1KHQCzJheOwIV6TY0LzoCBdqHqnIbBo+g4O2c86Kb9aA
h4TBgqwnraJWb7zv/mPZ0A9tnNfVSoNQhqjgZPLsX2StfRJq8/ndnTvGejtpX9Me2OVOiAgGftxG
cj5kqrS84bG4d8sf60kP+vfhY8jduetC1ugHNLyQE97d33W5wbc1KHeF5cBUgSLwkQ3NlpkBNlPG
275ersXgCO7IRiTmPXbOKoPkGqSiQtSMnQqAL3Els6ClALiRqE++8CCTiUFEDUHDO/jC8HKsJC61
CBHv8W+Gu2ioqjFW7SvJbi8DEsnRyNnnF86EoalDNkA69ChDYvNkbY8oqX5lad2QoE9mfsiOnDBC
8KxGEhYP5nJQWA4LbOsDGIe+oSBd7YiClbsUKoAgbE+rHGrWmp5pAn2Fj/ZPhKxrbWXyIpQFw+Ru
Vax4atoxErepz/29Z8kG5eUTsVacrlpIYq0yPbHIW4/DRl+c50EwOJ7P7EcYbg4kwcNKGEpvNjKI
X9Hf3aKlgg092RgkxZ1YPvVOMN4OwjxdwDdOfwFgnCVTSMKI3h8FoQAbzd7PBuTlU8rPFMyVG3cZ
nv/r6y/acJR0jgcd3Lk5VAwX+0A63wr6NhZmE/UatnfLkKRlSaAz6qz+KNAIaWCegKM5j5tG5r9O
dEIvpnzfns3xT5h2ottfebw0wCEuDnacww2TrAHLg9Yk60+3aoY+OHDim8kpmq9hqR0FXlPZJOql
BVZ5j0mAFG4dxv2M/l89jybifNyyRrYxFRyn2DL0qFy4iC4IlKrt3JoIXgkMtOAgiFlpS+7YU5s5
nAL9VmMhKrEKNrabmUTEqEmjt6MXCBLwiPvanHPrETv5AnO3BrxX1lnCkhcInIA/awaMZkHz09MS
6nKKVh+II0h5HKp9b+OCqaIbIPnB/orxUXxaRcUUnKcucVPO+huSKJhTGS5ONmq9QvhgmwqCbEa+
damof4i/tGw1t5BQngswrpzSkb56okxDEdxE6Az/Eicp38Ow9TtV9PpAVir2uT1ZHb5PXiEStpwc
g3WORry4bjC9HgFmye1oaggATXRaCtSVC9bjj4V2tGN8Kp9iQ8f5+2hwwyYZtuC4k9BBC2dwwrxW
ODHfr+ogF7JqFjbN4TdDiq2XkOVGAlFl9lPU/AUv4naNYqTRRrZCv53a8RQLjvVFsZlJK0TZd/zc
GFbUKr1UThSqRvlv60m+Us7fdzQxC2AGjK1ARzt7sT3AaIxSzMIKcWYeCRWfoq/1mMLGeaJBF6t+
4pwKhLHLGVwXo4gYgUyeD/P6YYiBs0U9z8zu9ammaFM3suDTGm4lkLOdojuKgFIxFvQMuKkkrqrJ
Bds/29SI1xFIhUWvIpnekD1SymFvob9XcwoJQjESbBiJDDCMJzzgsXLdBPJFNrfgNvMWBiB6k9FL
aN3b4UmJvvVPpxaSdg3IymqvCJ6tUMMxSLJcsvQRhMNAscNFHllgLBlfzRoLbIDYriSqDNcSlufS
DLhAWCEP93sj4TW1AaK1z3snlEfKFhmYt1Cj8rZxFEeM5f7ZAR9feFPETm0tk57+YltA2u4ezGjL
naNMwbjcqIA/E9u2ZoyGCvoF/i51Z2p8i1FdeQB5H1YHLdIwGvXywmmddcFtMMVjRP4ecdRSH5Sk
Bo/fJZdyIQ21FByIsQH7SjKYdNarL4whTAdIOM8tgdtclwxAoEAtDWU0z/HqTnFVRZWAuu2GyXgU
3Q/ug83m2WvnzcIDxrzCrNXCSo/WXUEa+n2lHWkVPukjKxL6mP5kFrSr5bU4ht8e+Kjj70G1b8GG
wUjbR9lfzE1nCT3i7c9hgXk68psEESr3+1qhNRgLY7aVvy9Y1dxhXuJtvlW5bGWEoHxSfcoHs99p
fD8AhsGGeADBw+VmaiuWM7CBHT3f/R7ezZn9SnyLJS8Qi+f0WNg51kLLTn1y5OIoikN/ykDn4etc
Hxl6PxBCKJqAjbVRN1+rGFqIwZ+5LAxutnCvoGy2s36odXBFl1YZRX0GsTSQRV4MYHiQBGKNT8EB
tofTqJN0c9wiTnS7UTM3eQB1jX8GBTDnbsFOS2fOgTkRoIv8LAGCVlehErr/yOGi8sEy6b2EiWHi
dOVIlC7Fm3dLvCjrpwPb/GHCA9tW/M4/+YK3uE8jYYVcticgjLQPAovs3k/qeIvwEFtsk171vvBr
IJr2phGk0hiIKg2t6fcBoGtvzSjyAFwLNcsri4wB+nk/Gv2bVgMVWu7g5XvLo7lQBJL1Kv9rQNxB
NCeC5dMIGKOIYfO8M4rEiz8I/0wFjNLASlS1sJbH5qGzyRYMDS8r/PJ2c4dnsK7js0W2Im7hc3GY
6ZsNUqoH3YQ3fsdO/YVgdgkQHfPHLJ0RYN+Nv6t2D7/ao30SogR8oXi5fm8AIK3hPQbJ9K7T63SV
2UNWJGbQxSMLFd/wrmSnT2QHUNeQne/mvXL88VlGGFk87doQtlsenNTUg75Pr6xlLWeggoJwzTl6
xOP6uw1rOK0Ev67fn+zvvKt13P7Ekysh6ACmTlpZThplt9DMmWz8PO5FyU+ng66QwJXfn7wfO4Qz
NcNDsTLaSKpo7UXh3YESFli7L8JETcdQgGdwTeW6iPKV2agkuV5tq4vVlY+GDDBhLvGIQP86lq5u
PIqo1rZOH8xMVvViX+pnsHxGKr558AfHH1qIbaX3CZwCBJT2QVj8q+J502c0nH2rpklw60X1Dv6M
DgbKps4wR7ympum6PoNczx+8q1NdpqeHXoSVqSmtnIRQDrnBSeUCP2iR/gIgvW+OGHJ+9Vf3sfUW
2f83RZZvnG5YGZSQXWg0+WkS2igGkRGOeKtdR2Chl7GrpY2dz1TrMMTo6R4zJgSTotVDI7vM/5Pa
jFfvfouakR1z+XT0bvHZR27xVDmtolUQrRR9t/oAgnrQScEIgv/thbZkSVf3hJW2KCkvvncTueDQ
ebf4X32ba7QI+kn26fw8TQ3bfOG97hX8GzX601R8QFkS7fygwjINRESTGyBLzOBNFAIag7BCzIsY
AjBpXTsQctxzH8pCAdnlgYwnn2f21QaY2ajNsOgBuHpd5pBWAlq4aJpKX4x510IiHtXXKmApQ/XS
YVbRRctWt4Um7/tTUVhXuYXXzhp27bZrlyQDSeH8Pf3dUbnYf1qAPenDJhtb9ivtPqhZho3N5lBZ
C7O9vI/2QW/zEfoqp5oJacUxPDQS9e0P3kbb96zL+QRs/yp8I5A/6dIpz2wABt2hkiIkUy1V9W4s
ujO5PRoxODcHNxHX54et+oYq11N5nv4Mv4HCFjg9BoiNFLgDwAKZRWRV6TCs31fo6Rlg/H+BzHHG
HVUly9sENS1MnVHlius666KWnHuDMzRzeX5wLmCKdXEugreTwE2HOw5mDj+PJcGmuvZ7cavvdxpC
Q4DTp1MiY0aYwGU6CtueB6GX2eI5fB24J080CfN3m52jv2YvJSvTN+0JDYYdjmcpm6VgUZvk8P/q
lXaZueQ7o+r7lT+P1Btq4gKtxlURstJwgLzwXlopu2dDuF/ffWxgQoom7NCjAvQE/yGFCOGTUgf4
fhE1hfEsZsRe4F3C2livsBEQWvQvZWUBDixqD6C5rM9LNB/3Er4l8wOkZfbhk+xHFua9DxpINQdH
RZfR/HVUJoV+7Gt1MSsx5mHTml25DJYPr9/P0PmUY9yN9wLuNQLetNnYttQ1ErqEbXJ3H/ktVwjT
ilOZzlwPHqzDxqIGOutHP+wHORzO4v8CAv8zlJ7/1wa5taW7WuNZLjPsMUvuOUO99NQft6/aCjab
VLbA5YUGaAjEg4L4EpJUA80Q3HuR18iza4NVCCT1vC9c0efOxdeuTYkmDDXq0unesvWUrZnxkizd
mt4Qq3VgrnOc3psd0JnSkwIfO8jvvETRj9pqvDKNHWs9Mj9vSse3pZXMcA3YjGfHmjN2rKgAjuHL
zRznHNRFw7i0yGH0IPZnKPi9LNC2vsfGu799rUN+p1+J0tOBA192F9pHs7H9UgUNqIT2oAna2Ys4
oSE7KcBA+4ta9q+csJgOK2johyugj5CQRaq22xS8YfqCh+K7UiGL00Dydrgx+ZkxAVSvejCtrr/t
94PA6xYmrtsfCwZuKjWLDFVpVkENpsfaSdT1qDAdBVBa3S5Vpjax4S3X9PlZkbJU+1Q2UU88mTRL
Ux2XvF4fm1kylgAJoelaBl9OXiqO8wFruxZtlKB+5jhuFI0ABt9ki21ZlV8Eti3WLwEQ8P54JURt
+xCxfkEtQhGN8/KZWeLGmOghWF4zeSGXPrp5vqxy2jgk3tEwzhC300vMWX4Twi5YgMh1yYmYA3tO
gSCvITd6bgzWRJ4WZDTGxnjBdcyR2p484HuYJW6UsIHsKoWJzGKpVYCIrD1QYMYHmJl9mRL1kJCR
QA/UlBSGSMXPV91CZ9l4jg4AUw7zoXuHeSB4U7RBDad2tKgpBP3+QgQdt+664GLqlZjr9kSqSJUp
JfEUszEtYOS3vZO8O3tXusw4UqLNGoG22e1HHiAS65sx4AB20kNJxNH0oFKAeG8RIoLltayHUkZT
IWIaukec32FX1RCvVxh8pNhZ/HOooL6IQv4ak5X1v2Iep2s3+q6nOjWDVvLKHCoCerv24SrhAnaI
VNHxCvI1XKYzVLdt+h6jSTJssIp0GyBUDEIXQfo0uOBG9MpxOs8Ol05JKASzBI6xtXZis47+/G1J
/o+QYEGNkNKTE0AhFDanokLEX25waywGlnBvmVuIFiedMSgq13Lg89tQ8DkiNacssdPWTqKwM6xN
JlQbM9xyqOdf2rZ6rph8e6xDkxW0BvNfZUVqrOAHyuwuKZmEDNw9hKOLdk1l7m/0rjONBDNF4Ocu
Z+EX/WFyczPHO4tsCLqXbAVwEkEaMthxG8qrGC29VmafI1OYguoZJGRwF7fTAJQCq7daOmdDobRJ
MfXdz7agpMkOXAjwzlPiupftM4qAdLYbvCWIcIy+MsIT1VYTr0Y8+UO3Ox/JsNYJRlfwhBhLJylO
7IQC7liQW6yx3/DdqPEUkGJDRJP4nmIDTnHGKPP5NHmmsCUNkcmnbGC4E2WjHCJ2Z7RTVGCXxqt2
b+L5y4qYGwvDp6KqDmKr5vTkYyQ3KSu8WoGL3E4CsznvFctkKQVIetIONojZ4/uofzNibYmUnEC0
FVTP0k6q93hd5RbMdYN7ZohxLlGNK/NGprnZzBW/B4ekCe6V9rHT1Lhs42ufp84PQqm7z7QS0fe6
bPgYhTPCncsM1GXOxEC+F05V7bPZDMJnyh7IKd8Uq6/ELGMoUnRSMl3sVyudeMhYxLf03oFD+sZL
SvMTRZblxoL/JIf92o8vm//9UoNLsB9HmBc23/dirvd/Kvq0V0kLi0CiPHduSnSEb5u9jjYUz4QA
LNyn7FcM4XqCkBXn0zJ93sm8aXg68VrSwfygyElB+jY9KFB+Fg/UEZC2OWfyfDiqejmVyas0cFSP
K04a+LMM1fntSAd95BlQLmoDXCJpDtKA7ZhUa7tNPS4H/gAgfF3IEYOpgWt+Y9vpZ0lo5ti9u7nc
Sb7pOXlYrmg+Rp6sJpvPe58Rg9TMvi+z/x2EDGDxLvt3Rs6rWc+eb/+mv9d1YK2VtfzmshqPx6hz
mcck7Sq+UWtM37TT6R01KXWr+574Qa+dbm2aHCuYyKT3pPnycVLRaqiF7h7WAQPGxLjenvDBj30E
DAwDONC22XLKwRxnaOvlA4BQpCUT7BeSEvd4JWhYBxzWdBzjEvYdFubOoJbmb6kSXIULJ62REhnc
RQ/nhNf/nr7zpCY95giPifxKGcxOnValoCyzjGqm0G+EDtvSN0Dltdq3PVzllMt5MifP4lfY+5xT
ks5wQQk5/aUK69hFHgP5vPl92xe06fK0zcNfwo4uL6p4n9+YMM1thHKEpLvUgiy8dNTgrXhuYPS/
Gmx3Mjuq/GSwejjwFgJiKxAx/MgcFTHKbayCt9d+qIjWnKn6f1UQW99izK7/tRbBlvP2cW77oDqv
/jp14fdmiOYxOiG1gzIryWbd9Kc52Zs17Aq4Rjz2d8asrj12XdgBWWOIJ/cXAwbTtIyYuFuBNu+0
YLk99/xz3VaruBd/LjhFUcXAjbcOQdIZDC6e1HtFN4gayjt0c2ZRn1kuGaw3Gzs5P088PelXmnK5
MqlRBWS1sa7pLYrwPcqSpOzO7AWDTWSyh1xBvUK3YugEU0Y7/v7p71OVlPuB4861sAxrJuun2S0O
F87G6QlaB7WR4IP9SBTqhFxc9Z1HMkK27jcYOsLmG9CQy/LcemNOcycdINuLrmEgSXa4B5QvQIh7
1axjZ/aDB5LGF2yn2QXj89toFlebLmCkSEoN56KhVaCkZU3Ym9E7imd9aykJVPEqh0Mj14HYetti
k1l30fSD2ra+2nTk5/lw5Mb9YfaVrJn/PiZqkuPNEdRiUs2CJhjP4hr6BcKT7jCbQiZkIH8tNLub
DQaA3KPIoku2OtJOKMb2tAsU0e30rmHyg3WuzZhclSH4Fyj+/QENxcHXQ8T5UfWNyf67hhbFg+fq
rExQLFEAhJoo2iOz53+FBfZkC8RJQaevI8wS75hPH4Ci6wm4Dq/v916sQo3kplbIJMPdPW8dAJFi
UNeKfBvK4eTN2pGpnsOZml5d8RvzLsuKH4kuyPBEEZMnMrPyR3khD8YXDESORbDrthCEx8kWSrQU
URV9NXoKoyzVRPkYTvcokbItQ39Tmkn9xOazJli6D89up0xCyIP5yDIRoNR/Iorr03k9zKWg0Ynq
PUgYDjQhWPy9970RAZ8D3hAMwT7eSnChfa/ebWk58eIrT4TtNhI7j+C6540fYQsgrwyl/4QQ2BEp
U/52t0kRr+Z/XFnkn1zJEtvfSy8Xke2WQsCzwzvjjItgco8vTPlCOmFPD1KA/gsRu0fuyzOEegwt
GLddeN6b2CMYxrYgwNngEyH3+xdMaR5fE8neOmtIFSeHPhlYEwaaFK0POLqnBxW2KDvO/eveCSxx
yQox8SJS89cDgmMYHiNNnuVKobw3S8vVAjGSNI9PGNyDsBXggYfDefx6t6flEJXSayK6D+xtpdF1
E3Kla7gPVy3QK0iDOgaaWZkpznszJMXoKb5N6R5QgkErxEiXM9YH10cnFu+WPxOItWdbzATdmJHn
WbpKa96DV3lP6U3DSW04yaJ4k3TdLOKedmT797FZLkOGASnttW39WWMZaS6vV06msh4klavgp6j8
se0MwrKxhhYCA8dPjgGNOMYAwOba4R2qO4aZ/1yAt6gPgYtvwpRgojDs/zY462RwaiTB7/dwQVHx
TtxvcMNC2PO5G3lKClcLCJ5cXAYWItwR1lNkvgRAQfD2ezdhUru49J3WPNXluUTTnsljXEXSshoP
XijvGbEcUYfgPTrPJeMaoaP94E9Seb6fZED+h1w5AgLO9HTGhfbISrKDmkJ321i0Aioov0Nd4Fq3
DeIcaSKV/m+Y8R3Ik5RpEVzeW+m84BGtdkpya9T6xXHguRSL0P+IO7fUeFh+Jx47zhlacDKCrODL
ew0h6PJ7QI9Y9EFUhtDXMB4gwopNUs0WbtroM9GISxw+cw6fJ46iriTCUYw5rU1sBeIKiR+8wWqN
YLsijDHSWfX6WmJ3Hz0TyFb/xMRn0szwlOMVNn3hH3oTY7WpgrdzFZ+wXutEDiAg1qatrs8m/WL7
6/umFOaUz1ZUSLkGgrRRV1VWVAsGgd7rxjXTpaEjh3QM4+l1i7lV9owsn8h0eqt/bs9UHHmj9DaG
VSuEt8tMmoo110A2/Td/TCvZ7Ov9BhcGQzRpPD+LFlkhjogc3Et1mu0W8U/VbdZo0FSIFlD0szMv
5Vchp/kATAUh25bHtjkhj4RuU+a5eMbC/D/Ad0XsxZeLnXrHlXzyf9ttXa8HhaeZB4h6OXMQn+Ya
0HD7GRuVKutGwRMgK91yX8I9GBtpxT+F1O4abxq3Rc6RIpYCddXiqarjiyF8h9nVgkmWRvE+y07+
BILdY0LraGnCM/PYTQPqv9QyHorSxW65V5DB1w1sm1EXlgxNRpCY/qXru0pfkAYyKObHsvsHgjwo
wb/yZItdtBT76A+rjUXFww6u533tai2iT1r8fCdyhxfqZUaE8x4JSIZ4CUxCNeL+shMX71jFiCQt
zi5O09Ns5Ga2m/IwxqS4rG+VyUkcX3lgFmj0nwEPZg98tgPIqPX3WBUW/tMHGOC+4puJO9PPiT1D
Ug/Qul9/QQS0TkeZPzjtHo6e6NO3KH7YkpLFnFNRunP4JQPY+jLmKLkqT1qX1/39DUNCTSzELE53
FRE1rbh//BofaCbd7wshI459tCI62RlFCn8UhawOntOG9fAKBJ/XvxmGCM6JUCJe3STyUoOTiiR4
vjEhu22LnS76PrmRYphI48aioDC/PtLZ7AklcyjeqpMamkzwY1spjV98+vY6ajSO0/f1fB1QXTqP
oM9DapP5SON52xs6GRHJqRJ1TG2dnCO+V2aMGwxuNh22WX5bxcwcvdReKwVF7WLsbQ1IZaHTbZOE
Bm5aa28WfPiralyBTb9DQG8KbmTXUMvW93QJmR9hkxYOiBg6CODX9N1sWNd+E79Pqu0xrleaNB8f
fFqRU+93uFJFo64wVFNJ26DRfKqtr5vP+hNZd/D57BzKukucHSyymKAugW71trTSyDMuZB2wC5aF
c6efTfN2cyS0O4aYTXqaXPREXE/yEcfTuzAOaiHUWK796VKjIFZDwgiRliYfF99q0M7HjXDJVqrJ
4OjciG+cP5fkQeqVvV4sabYCJuWPPO2bG1CBihEylvKEceltHOJgqcNtaovh7EY1YaMLNuHb7rqH
747i/jsdD7yyEu3D6E4e982GE1/KZf8SPCZ1Ufij8HwtF4MXP1LW15n8HyyUMtEYnG+q9pi57vEy
3YQ34ZfwA8eJDPxth45pry52N/RzgWlnAyLb7suuT8VC7nn9KFcyOippktkd9EzM7t0K2xWD0rBk
mvTZ0M0SMouwwoXPjXBs66SQwgB0ocWvGxVJZgRCn5R2x7XN1xKfMPdBnAitKYoojpOD5qH93dXi
1q0COJ4SkaE8bN3ob91+eFKz/cqUfvBMaGh4GJnMSOWe75BJD5JQ+9s8Ehs8HCjlIGpCSFFiadTu
+hFvWk41mu1ikGSIEJWYezn+IFaj2SKl+R4M8woZEUVzDAXPe1WnUqKzMn4P8n2qaGrJRGGXjgfO
U7KilYkk238fSRZGGcPMst+oHwwTRU5FQ3Zf7tD2VrtqZqYuLT80D04GTVgDVlPArkpdjtbavysk
t4VtD4BQz/GoCWthw48L0qlBFZmkkPRR0th19NUKLwCSqigLu+adRF2X8iStdJxwZqz87VP1vO4H
q/zplrs8t6IH3Ga5FO/QAOmFCzYCDkIWEViAG3ICbvZaocfb/gVX5gTSZDe2qkCkdcG0ycPu9aUI
nQwoEKa8wDcG27YDCdL5LNe2POPtbnXd/ycCoPBdF6EY3OI+ZIl/v4egHcjXFjUjrrp3y+wImseY
BzxeJTg3wks2vz4dSwpgsvldcIJQuFeEXiDUXiPpKBGcau4pBtuQHUB4upGH2H0TZJy0soMWOPB7
kBKMi6uH+qsJwpY7ibK+elufZeT+9Hpf56sKKGtstJwjvTxiGueVhCIQSbInE4sX7/PReoFXSkoB
UkOs5IH0L5WLXwmx1DVCNv6/MCCs70YlsZ4ENuTF3hG0MdIgSIWJYBQgpQpIQ9CYqpyA8XHyVurt
pZjrP1WTeYvY67zC9pohKzV/slYirH6etDit6ldqZNqykUG3jxu5W1sSy2lz3BWIjtjTPGHWRX+I
ZYGcTGpk+hzoERK0xt3nOJIXgsUmfK0jYVhVQUe/QGxWfC6AIovFAPMhSQFQVoOxDZUf1IeWeg5x
2QForR+PoATHLJhRSBAhVdf7rIQVjXWfOxq5w7we6dw28m1lU5VL07nYKJexUfrzRSSbbH3YgPXo
VnwbBIlcFBYCTbS6q4298uKf8ioCWu0DW577YVrcdQE7qu/1mivAe8f+wFuCJEOGDUKBRieqhjR0
A8tGnsUboY37OdI7aZuKxspeEQi8jlGGYyP78yGa0QpJWizANMZhNCtWmBtKdlJccVUFde3X6omv
RILx9nyKlRmOO6x5VWCcpujK7Vf5hdUkqGT5LH/ySpfSITwVRcqIP161EPvDfFoXKT2BjWf+bz47
E2/ot5p2Rtst/MRykN+TAwPv4YDitmkiQ+eCwxsLBcSZe7SzWmxAvKlC5+lMqtj96KiXDICBrX6+
1JACjPQXXOONkZWWDPU/UEbGlRt2m9TyJ4tGLnDHJkOP2SESqzdMvn3YI9t50g65aOjS5Cdyk+Ug
hEqdS/cDgNp2ZGAZHfDaTBhsrwgI359onEqj+xwc/brJf+xKBi9ygwGnbWYh9u1Htlue6Xq1M8nz
V/sTnxs23fEiLpi0AoKcAUaXoHxrMJGGRyxIFyiqOD/xyt3cZ/bFUg/im0WaeffuXJsRkMRNhZ8Z
kAbO6/QtdLRXf/Y/fW3fLzke0wQSwRfpVWBjHB0qgieU4J40p07ZU2ISkPW9wA1jyTvuy0ZNKgOq
nYkGohPOay6zKKfFYL4v3fiLiC6u38djKU0Ygp59j8pVKg7jGRbj9vqH4qIWeNZAH5v4HY4ZsVse
/jGuvte9x5oQuLY4b5L26Ye5tT1pz7M1nNkbBE+wanJse2FtlvIQJ/AVlv75o9FCVo1Gr0qgXA/O
ZBLnQKEZ5YFggQJsfy17obOmZQdEk5bnRKXwLiBKpVjP6KwXrDAe0bZvPXJXpmo04Q83GaJbZA8v
k3Dc3hposz2ZV/dr3AyAMWylFFhUdcOXla2Rhyi0qr+87br0OqI71d6n5N9tgg7DZZ1CclUha6Fi
ldnja/ySCZzO32DCB81V541+qvf3F+R8/1aXTLPSKVI/SH0+68ycUF+J0L+a7CKJE33u/hk4ihJR
tfm3iBAJwmgXltFI7+21TYdtAVFtnKDSQ0JkwAVWPL1UOSRg2ZT2AnRMKUKpps+49EfnFvOqJUt2
1q8eW52bPReu4gKUHF9Y9H7hzGi3AKqS2pnZ/cUsWbYvLElD+e+4/zMqCF0FBU3o+cyJQiPcPVxw
8FKvSXWoym2anUkWoFLsAQ/jRheStFYZgy2g07Wr1igNr7ET8n8bwHFcyvVg+EP9KEWs+sMItMoo
9nPvrTDDbs6UNCE86gZGpd21gFD4tD+FhQThM2YplBRfOFlIGF75eAGFv+h3z/BseYS50o5XHH6t
ikXNv63vmqORzJMI2+ei7JH+34X2tht8fb7yf8jfoQ9IA6+6cBuoyCPrG32f0gc792DT1zzUqDrx
JDErhbfh17LhkACCiO3VpXfmgB6MQU/RqZ+ZyZ7m5/EhzOvlAQxgS8pp5FYOLVDbk2+vCAuJfZzp
J689+em+TUf7VLOxfQCqvt2UmwbkE3E6oqGIdGU0MXySm79se2N/Pg15osDma5R715zcquUrlqBR
lsqiAXm5UCRSkwNo9t5S3zCq4TsKMJhetJjY2eNxuGEeVvFW0d/l81vxn/vC9QAU5p/icYPqNaBp
PbAP7h0JGunmZWzl3jEqa/WHr01SfbBLTedXU670GDibvcqV3g6YOSO4ZT9OeeKugWzJ7Sd/D1Bt
2s+bNr3ESbIDSinvdQe/a2SN7q2q6ILdzOF0FEDtl2DuFpD6lSpW6r26Ob4Nc7k3ICL/0MwttNES
/7nJxi4WEonlC8gcvBahxsgvgTvH9dqzzIsdPsBRCwVa+PW5TCMUCY9YA/Z6wMxEn69d/Uu4PL0D
oxlRI7pWcuiMJnhmJgN4XdXpmOsclX3UDaaY2BJ9eIZYu2+P8yeDtx2v/G+Cn2AvQcLaTk+yBcIg
RWBLFIHL7gceQ1R72RLxIekKnG3w4vKuhViLgEBQ12nNKhvIOcu+O39njepA03TWigdzbaOphVfa
HGIU/XK1JN2/c2zi23aB0BnYCoqWuvL4p6xxMi4YgRj34tyG5LGlx0YUI+aSLnhWLdsgIQxNNn73
OcSMXh/8nnXbAt0aH3q9jiiYR8HilfNB56fGUUWd6ashUjffxVpmUkJDBOZIqJ7e9LYg0o5swGhW
nd2BswjfBujYs4/uSOh6iLEyOsHfmI/rz0IDAzFxUfVp/A1iXa0MYrMe5+FAuTD+94UnLssTSqnw
/iHCePE2zUU1crTip4p4rOJP3PrMadKKdUsqSd4MeLrkhf0AOqbnPxcsMonUdLL+VnrTRpZdScTf
t+/pyAK5bxspgOOOJeyVA+R6RpmO7saslTvJXnVePBGH1iOe8IkXCMOEpkWS2nTd5JLhUQGNSH3f
FNiY06bt1y1Xa4YOP79OQGRfwyXf2ZLQbzK8ADe8HpCVoPjC8ut6LADsA0WOj8bPkflGWgVuTlXH
d0v4979h1NxUkdQ6ExljXrOemnp9bsfvrM3d6F1sF7jZ/xqxH3k4PV8k8ctOev23TkPRtmV0UWay
pR6ip4Ni5lkwD+QOZ4+J5mswOm8ni/jBil+qZHdyBpttnzpw1SdMADJofJZX+aKFF/OjZoh9mr1f
51b2FjbP4d3xMyhEBkc9XNsBsp9UcaxAk060uouMc7heR9xbdisjQ1o/NLtzWnaMz0WqbGH37TOA
PCMMjXaDzj/Vc9EUpcmW53wKNOqsz5/EqwV9iQGsr6NsW7sB2ySxZiWohwDuJpYOqNSlBC9p1hjU
o0GKe5TIp2DGuI2Y6tajwUdgjyMW+JAJrmiDoaOAo9/8PNtT32NlnQCPjFqY6WU/hDAPKnWaGGaE
ITDpxu2vH0YFs2NWADUwvZvmbuFcNB9qGp8BKh+9kIk4hnTS6n58HOVRgU6r+/DbCOzyLX6xtMSm
PTn9wXCuEZZ4dHiyKzZ7Mls6EvrCI6v7pDflLKDdEMCUccm2OMY0YQBqbAC9dHK5J+EW5krLeZ/C
nv4/SjJ78wPO58YolTSeTn/go2aCyVVV6argnxXAVb6gi08I2W6EZuWwcR/R607aTE0HLgxd/iaE
NaMEkOVl45EOlRPVL2eV4GRhErD2gf5Aa5SHbUVU0WDdblV8mwxWpPg97V14bfOxoLZkX9VWVV7s
wjZiRshysxQpxkjbJVVw6bgIfCT/G0KadyruG38KUJrjBBtfiFLHXeTegGchcRNLrBp+egle1bt1
DqugemyjIlTfgAEkOE2wo4emv66Kn5/PlTmfALwjjLCgJT4sxGK22XLNyoT9U2ukC5tiJ+rHoxoA
ikMTZYqmmHCIpza7b6vPubBsjd6e04AfaR/CSZLuhdrezP8n8HqRUOj31spABOpUWaadXpAr6Zms
yHPiWkWLMFZTY35WpzYmABxKbDMWntbPeXS5ilYvYwUuQO7Jx+GZuKV7YgaOr7WmXlbtgC2xnEuL
CBmXB6ZEQ+0vE4FGhU+dJpKOtLmw/PNpgaLqjVNfW4z38bzIdcbinw8bg0XPZ6w3dt5JI2Q+1q05
cyBtd5W3oshX1wJctxuxAcD6LA64TmsoW5GXzz2HxnBDlYw0srtZmyEp7+qQ5y5+3z60ulPpAphL
3qsKoHPzX2mh5GGBEFH8Vs83ysDvxThfiDVY7e3FNr3sIpM5SgPCZ6wkakMa1jqCZ8ox2fXrMKRH
u7OSZlXCuMMfKWiFGuMwb9o3270P8BRk94RXLL0MvrE0erV/5kQ2WeP+F/Pm1E/IaJ1zkMsrQHKN
OMKKlkjen9Q3TOTHBNmuLJ+Xs/qtTDdAeUVgzecbf/Ig/Xeg7xoud6VZ+Dqrr/09uCwuz293e4L3
qoma6Orn7MyWCjTXTcYjJWj362IRQJ0IfF+t+6l/KUREeTjn38Mi8W18T72oGr1VYFrmCUW7F/uG
3DiQNSSOYQcBOPp4r+s8HYEg/YaoKTOXlHGpt54KLYo54zuP7t8g16JZz+w+wFEOA5+xaGYz72Wh
/8RfGOTRjrK2EB0zCAsuGc+VudEFk8l2bvL4iH7BAiUFy/m7Z38ZwAxxMh/mAIj7rGdxUr134K/O
76XoQhalEdA0faCXdI2HZPKvMTye/StmqwLiBYHgoZ19OmBhHX1gR7oJu2B4IbKLsMDLGkuzPcZc
PCce023CT9psj8Y58/56jv9Ho8GLkXsor0YO18JfqyHzcFWi23ySucL6rDph4CzPZABfQmhR8yep
jbRlS5yOKRq+Gmpg+IoObFdwYKLKSoaMW99XmulCOkiyCKCQbBagoOvt/HRfLktpeFK+XKZ9ETlr
jK9MatswAhBziHCNqkDQ4UNbmfDtCQrrqwo4fu8tDtfmo/BtAlBH/LsvPCU/DaxIy79L5ivR1Utm
gAIBiynsDdFF9N6XeU+evPmXn1XqaR1+wH3KVvvT6B1x9d7aYpWKSWy7BDfAN6HEb/GkXfBV88lI
WjOVHU5fxBZQqDZB2OfvtL861Uqq9fFcy7navG3v9VV6nhkVrAWoolVvabIzf63hjm8zaQmGsOn7
w0rbi22LB8CP1Ozd5L3fFuhpnQw7Lhc67z1meifvvN+OVlegujFTFULW9vm5hdHYmIM+qO4uBl8K
ok6epWFW2MD3mIDIhgg0gCQPgPt80paVV4+KeKDIYwqvFsDES3gKAhlrxOimehJW6Abtv7e7GExv
s030/GAu9QOUnhc3vGusUYEli7JZN6cvSOZMnG6gimcZpDoorvwdoC9ybMkF/isX0L4joMpplJCD
+v7/AOiNP1hfCc1uUWGk4czupk/zTW7VKcjZjuPxFBjwx5ajUe5VN8aDZdvwL+O2D1hTRjKZNkUh
QpzQR42aObWu1rWf/wvD5zmazjPh0fStInUtnwu60ws+lG6a9udAEy1GpzMJcxHhGmCOsr6+ieCp
ipeXXl/XPVZ1lqqULdLxeQzBv3MKFJZmK/nsAPZZ0bz6rahQSNmX7YJwZgoYzGFclStrmuQMSUw5
x1vARJ3mwj+SjuOyTblMCB9T4e8DecxgP9Zt77u1Xhn5cUVPca0kDnyXw+BV5yf/WkeFcG57Zz0q
6/pR0/JLxYl4hVGYrVCl/5MdIKWoA1X1aUYvtZX4DKnHTgXn/5SkWyXtwm/h3qDlhguUcqgmVP6m
2u7YXIjOKl3Gcz6PY6TCRD3GFpOGxqG9wvirdpz2xJwsq4Shl81erWnPc3VkeqIGqGLAiMhH27qG
8pP0Wfhc42dr2qGpRZ+VtvBlfEt6zquTPr4kgOC7fQhRDckWXDtCnHrFOhAVZklrAWpTA3VSWTqT
M0pO/HsV4H5rpXf/huS16NICDj0dss5o3UI5wKK7bUjmvIw1XhN2FdI/iGAi9DMzm5Z34WuscIZ7
hezYYEzRmUT1VIDtj5z/ZE6LSktzoXr6mzjc7/Wg7qz/NiL3OurZXbt8bS1BHgJSRYp35l2sOHfi
cvxAt+qQ61WkzPJvETmn5r3YCIO5CuBN0+h2r5ngzaK9dL6eEMjz4qYOmhE060BQH1780ETmlUfv
iTea0on5OCYQQ8aWmb8hvdKWIT9uwJpSVoPKr98eeVKvf3t3GLtlBnn16IkTxKvUwGzyNTkJbbIe
3D4VD3IHAa50ea/Ew/Os+SlO9FwJ/v13vU8u739WJB2Rvq4Q8Hxrc/5smv2Q/NiOx2KpcR/rXvw1
vrFE8jJ67mfYgpTQNXwZXa/5dr7vFfAcv+N0nnEbc2KUq7LsNvw64PmlMECh3XwK69IlqBkK5xyk
gd1DyvQ/M3D8HD+53fDXCRvX6Pwl152+OvZXvHPU7RLl31eoc94cMKznVjHbks4yeYEskDScGXnQ
w/0oNQLwpFh210yZWjPJtM/dz+rYFACMl1K9tfPbZlLuRqKESCTaO+Fs+rpBGSea5q59MIdbH087
Gad5VtuKWItwi5cw6TkyOrl2/4QoT2MaHDkFF45rVO4Sz043aiTnAbAG4t4XNOVUa5pXK7GX2b2A
nUdSRG8aCI5+HbrS1ZDUZpUdmMRaOr5ooH2PdrQVBGWT3Pj3hg2ejAjTUBoQyA/ARpkVPoj3qyYV
67bIx0jN6fa+QOJe2ynDcnd4BtknWoJvjhqiXNTs3wQQTqQJwP/vYGWlx/fEkd1D5asXW6iYt/vs
P1GmyA0P+zFdDiIQF9Jw+XdAOEe6boav+z6XDimCjKlgNAtz5EVj+34IMCbnvaG/oes6kY0q2Fmp
NGGZwKDpGRkjsfJSrKSVHkETTnNdaahrQfeXUs5KPDr7bZ8+H+ozJb0UH9qsqvNA5ZLzftj7Fagd
PZp+gr2wpkrO2MYNkX7ZjkGbCexHMbal7FXKgwQ5uOFda7fqDPPVgwOnpEu+Teii3Ayq4wDk4FtU
85zx8306dKXcXrwWq0o6SZx+t9wqKOKxDytw7g0AwIROXBZfHs2dZDW771lNBvM9+8DkKzYVfSv3
DClkvcH7KLWxd0wdbzFQ6CSAkWCTX9F4j6ycUUfEts10iMKNCu/JCCZIj3CVitCMuwC0aC4lgrTg
tIUu2nnIMwJPUHQBqeKG+XohHC2JkIfGy/ardIOQKS+a/e9k1yLrtdMtZP4Y4gjJHBcnEvQFkIFs
bx2WwDOlw7OQm9HaVs57ipO1fSm5/iiHF6Q6pryQDy/YDqlbSZiBkPzjOeHCtNuisXlEeNIc6WI7
xAEvw74DTQHefTJ1HZlIzEybab+Wv5y9kN0ummyCr9evOI4WKHSFX+BM+4u2RNEeFAxl/Gqx99rq
e7bbH/epymUsY2s2MQ7RbY7eOlgnzKnUGDP7hQS6s42cH9mB8jQtSChwcGTtaohqAmNy9IXrBdmR
rKpa3nagoRRcteYmo1lueJJHMWbeezmRq3wkvaQUL9FDPN+wGf8WvNAGAYDDe5TMK3SaiUym8NmV
wMiVGv04tNMLNZ3xaO9wLZ+aTRk80riJmD929jCaYFfF3idqmB03jcUvvi4+dPukh5p6+eeNQO1r
pYw6pqYSw7wmbPfAQ7bpskmvJ5XezPnJVL9b6yLdnTjVAsoXVnPX9oJdH9B2kaQQvkdSfmnxLY/Y
iwuq140gZHoWLuYnn26u2dZzwjVcKOjBhskjNd9caLKsB1999l3BnhK4JrAApUfuZuj58xwq3i5j
OHgJ5UVFH7/acG0amm2Nx06pTv8gUl+HgS7V6NFsBQVL7IjAu95F7VC4UXUwT5kHgPLytd/NCIfI
nIbQVwhKpBDuPeiF69wAoveY966hwmsBMSv86LKrJaFPZrG4I1K4d1QShlp/9nFsUEfrW78g2g4V
b9Ljo8fy5sfK7iHpe345hyFS/ILqCDks7HqQZYs+sL+7G3LjWFvj6Jcrqc2+jo19UGw0gsvJ3MLC
0x66/5+fx92xVJg8eP16grIgSGbcCaIzWB571PcLVwogubBJ0BaocHFPnTFFmMK+55XyWjXANzBA
t/P6wEeophN/vEA85ZW3SDAG4yWMHQt/fIoEy/oe8CdIseBnwkgNNF3F7qXbqmprcVu3wrwcVpOh
w809ICMNzX7gEghtCTgzDeXyJs8G1iHEoPTF6pEq74N1hnz7NKJ5MsrdpjDXkW/E4SNOauw+57b/
WJPUTOGwy8FRpsBolcnjq/C2z0fQn2g+uIIbtFjfM913QNDHxkoJHpXFpDTKkIeZRq4Tqo0rKPh6
4/NMBUeLdOqozGfyKeW5fGKnJ7D8IPuV3OibsgBx46oT84aE7ERyQmZVwwXEqFHRRDkJFjwaQYnW
vKIOjDgZdXbq/JBVKWyHuyIwUpOC3RDjN2fTKsqYNlmi+d3icJXaMeuYAqGYV0Mr5nE5Eey8fiG5
u0LPgMrSXtADoxjdB0W6O+et8cghSw/FXMMI0WWF0wImvAZgtUhcnsS0XM+exyOy2wXUhjryUWO8
D7Vtj/rN+ANTgVEtWkitdfBNInlgx3xODSPfL/mX8oDzV7cPUfhztHIZXK8Ks7VounugOIUchWuK
JzzKLZgNazH5qvY4jdWDGVrpxiJW2OPV2zVBg9xuO7AUzmp0w/sL2TPhUhS9IpeT8lz7CPYO5VU9
OcZXF3/lHy6q4cwwQHLAktQYon5tQSW5+P/b1HEAmeVunkiOrF3/YgSnbNaq2xGKcSHAErbDEw8k
yHRzHBz0+4/0LkWUDJ/IVAUU3yc8gtpzIYVbgHEGT4h8OhruRxm6PRHBNsUXPDens0HJfVgEzFj8
sbzAJw2B1sHv+u8CJw8Vzw6y4YAAc4XVWdgwxiya/iy/lXOWypMCydOmWX5zGHVU6uIF7boOLOxa
vLAhbULJ4KhDEDJ3mrxgIB/KggS+hC25px5+JZdEcunrq/MMSUIVI1rMv9zxDCeYWAxjJT654u9u
kmQVG83BjCvl4uWsDd/i3OBPP/fKKgMw1Q4naeVyBbdUVQvsocmOtueK6k5sI25MO3tCFcwkn1cx
QDNwvVTOifABQluUpqWahv+t9VzOhHYOWI7jIqdz6cGgWmTWIhUNZlxq4Dl0PJELeuyH324H56x/
iZ3iCwQuYdknFj+dkUn0Cjo7MEQaTBn8pQMj9l89B2ASfVFUQfVZOFfWgfjza3AU6rsxLWl8wfMC
+7B1tf7HvTR5Ej4pwYW6CUbQTBfUwcemMJn+OAmAzuPbJNJJC9iiyEUC42Nxj1y7kMhzRpAWLF5F
rkfzDG2FI4UC3cxJgcOGJVO00XKWDNg/hxjDJcOS8JsAFExm2hf0DlsmBTFL8HofmLwSjUKsOoZY
QHEQ847PYSAjsLUwOwf4RTnZQpPkPnHuaVg/WFdedaqkxS9OFdEds/OL7zMdAxkEVTXSWY7/ajCP
/0g+C+jnYS5wEKFkRh+IqIBWy95qS4qGG+Jyil2jGh7f1ZgxdA/oiPdeSAtYZRZ57CGnF7evAX74
wD0pq99BYQdehxJ8RzSN11m60gzWYg2KPISpBz01+NfS7aa4ZzDzcUavJEAk/rsFOUUrDygjVfk/
XA9MJBEorEQ81wAFt+i5ITMPf0MGzdnna2hSoTmF3yH8UaF4ShitZx+S1lv5WrAQ3fZ3MbdWryds
Rn3pzQeRRGAynNt2r7hWZNJ8uhACwFAvZp48ZhhKTAYIhx/8D7SEfU3AuokKlHdP+e6PB/q+PSkn
UphveoGMsczwzDg2jFnrqLBfj0G2ezqZj7VTXbVuJvf0gbfMYcSOAALsiHZkjccBnyq1IvEFTQiQ
HTfDpy9hzzsCziuBVyz6c/dJVpo6GL4pQT/26OjjEW5qt3sIEIpzvUrlBlN1obFF2+ZuzwJKVfXD
jiXmr+rcqbvNlV92+Sqp8s0goZ70nuKx+YhZqohHpolHuB5lIXOl9pa8Qm1Ta5SSvPPe8pC4okHF
ro/HdHa48w3PoDAMn8nMpA/t/rHq+qMJOUlUlbSWnNSvp6knjjC4z4QbL1axk8y957iw3qMI7kMu
0OdjfFy5i5oslZLlmg9wyzm2C3IDJDZc+7nFkl3HIRN04qUS4EyRlL/v3p4cFRm23d7rcT2aw62L
PzkU+5a/ifUqQj3m50I6qlHhiE9lruv28moLMkfXsWr2632T6EKe/oy/U7WKZYAlidqdY+e8XzRL
v1Yxxmz/eJ/3kn8u2xJ2DDNu+VlmXkMkI0NjdOl3ysGWz31JA6BU0gvZFr/bmVM1z+/S7UYnCRE8
t/hg9QZoKu5YByiNhDf2BQb0rA/JHFjyZiLvPzH1EerBEfiTpxLf89pcEtBzRReRzswMHp9RZ215
vDAFn5kK+aw+gGYVIzNMRgm+7mXpG6cbD0CWAhhYa8yFDik2Xl0Dpt7VKmvzTGLdAxYLdCYknqBs
7PM1QeXBnollmS7H5I/g2DkId+W6tUtUTklEIRb2JNUHV7Fm3ye9zCjpR6wl3Zir6FdgTdtvRIQz
O6ejxzsxxjZ32mF2YrtZ8fkoV1bgbsw1YrgAbUP8jAYBCH81FhKOxb+SNFOOGOvxPne4/GDEkp+T
hiCv0mtQPlsUa/Ehjehx1MZAXHiPusZNMD13pWXE+lUY0DvE3LdLo8ndQyEpILhMtsQxk11pZsGK
3oKlw9YIbgdmXDzo1tojFMU4Knnh3c35Cya7rZeebG4MGcq0v7bQBjxGR69cR5QSovMo+rMhUjns
21AoIysDUG3f2kbGAazSfkIh8sLv3YI/hLyZOFWGzT0Ao2VWrGx467c23cz1mxiGC3oe+B1DcSi9
wbCx3SLxhSdIJUNi06nIF4LwOGhZbF730MYgP8WEgjklkMJT9J7x8zSfSGtkLQe4NueOb+09QCmJ
BImW5HbKyRvvjzsATJrbyPDYorMeW0KiYGPUDKmeqTb4Ch81Dj2oq61Du5vszECwqUTYqeUNotQn
9efTqF9W27FMQk2j3Wr0+maY8+FpVdtgyyv8K1JQzM0mKxnag3sWKdjjDM+vFk2bnq33g1KXDBuX
KKysUKmihW6uzLsuwr0ez4Q1jfRqrgxxHUBUQpjWPxf6c+ORLgb+qCcTEUl4EQHFGMaF1D2lWivB
jxC2Ivgt5ywcgUDLa0DKHeP816rYxyu0ImyWrwoDZNpNVpVnmwYTUqfxBU1Rq77WQ37HN8dvPYIn
mkfQ6USFeX18y7gvKVGfXtIX7Ban/UKjm19MxW1hSj6B8D1JzhvNyWuc1o46LEHFS25Lwc699675
OB/nSNVc68upueBSMan+coFvW7P1131Uc8OXSDOEaxt675tcDQV99dSU4RwFICRnM1Xk1/aYLHtB
b2jaMhTq228mmPKkzVKTBAqcXX+ezXfcDZQv/+70wdSnDubwgsttbJrN5vJHkkQtKF++Dvc6zdr/
cFtQArYs1/LFA/A6wiz71YGSoWjoA65+ExlRRPu/3WyhMq5fQaK7oezk/mDOFANeAvXBBUe30W1R
NaeBISDXlmdVwbhBc3mQDXLba2lPWCvWGfp98oSqewWOxA8W7yr8S0iO5ssoF33+faC84gm01gp3
rYNeLefCjf9on5wSEyhJ/7bTN+7/ozc1S12N9aQgyNdtX9xmN6BHSt2E5iZdPD2YPAUYm6bUP1j6
1OEfA+zVi0XzRJxMEJRc4YYMlNn8eqoU5V0KUyflosvEJQb56Emh6PT/WO7borBlN1XKM/J4XXId
oPYdoAeSk8+XtBIy/cUa+kN+0GPGnlZ3YwE8fMqegKgKCSMgOHeLirvriY/u9v6L3E/tOu2EwrO0
SXAwXFj0F1RKbrmOaiSC0TTRDVTxo+Stk77gRXRaxOhqV808OegqNdOU9uJBl4ev3oLCBfLICVi1
VWMxzmdaT1wgB6NOaU1D4Zsi4KFP2nXAYktLuSGzLPFgWQFY53SZoun4lZPHHDu7/Ecc+mby3bzs
M3hgkipAg5uunZuboWBZpT1fdONI9TPprfaXZhQNLc0S4FReN4tA7+x6EMG8z1Yp1WtIb970YOia
uV0iBPOH1YnLZK2ZMcwhaGiThy+mslo/n54ybEJJVu7ueM/0B1bUkT2A9wW/o95tgdIXgVPv/9SW
w73hXda713hoEtP66fb6WnME4lShUMI7G19j0pCujvo8pTSRWCJkv69qr3M3cm6uWeJd0JN00yR7
EbhdQR7YfErPYLQoU/uHcQLTJYKBwuSa9ZWAkIBtFN//+CNpFpiJK8r5OkBGbsi2JN5rJVftTGYw
LIp8Qv6ZvH6HnWJVFaPIO01OjASEfpstGdJeKlySowrE3rs9t5xJh1WX7vWVHqneZgSBbQ4Z5l8Z
hXCpZ25a6UlZtsX2GTLQ/8lbPiKabvgKuUoSgK2FTtmPLTds47YZuNzDGyMpvGkHeZKAt+d1ByXS
8Exvq++BNdsfSrNI32CP80bwZk7eDibPOsQLAB0tq3/00SswOn7c5rjaWa3WSWQDmSHBqkjRhOj9
wp6AwzajhsP1CfjDN08d8Zo5GQDkBwG2K0nWSRifb/d6oIaVWPTakkuXjLZ4tjYx5NlWlwl4nHnK
cPd45BrDikYB30j7LjYKlT1JHsT1B1ElU4zN8+oTGViOLEexQVti+v4+g32RVk/+jKIo323QcErG
EvcpcZj1f5wqHQvuCtLaPcKZB495mbKUgveRxJ1z/aN4vvkV2CfZoyncf/x+GBtZUM4YOzMPvZxA
q688pL/BDiStxdrhcA+23Pa//YOEtWxVGyXyAPHh/pO31jg0PW0kUbxDBYoajitm+JzrSWEDSMfd
EjZtduFh8S8Tsk8wlsByuJAfss64EQ2hjZNM6idyla3NNfamk59we+6H3wOejAArXXhvOprWNrqJ
OG54V4O8ZfFXpAjcHg2TLAW72OAi5KEvRUwjyGb2ZYw74hUx9dQsuZ55fJFsGvnFTqcCY5kBvCdz
EEX2s09ab1uERuJRw5AULK9mCt/XgCzFSZ7wmxutKvYH6XPVPQrrl594lV6ZdoCNyfuNuqUPyTGN
VxxmJfnPWytOd0hw6ZsI7qifJVALNTyvXSVkojuW/PU1t4ydq+FKxXNWa1PegCIm27p5RpHCUb/V
q3T1bNePKOeOespIQPPLwqcDownGmJDi8B4/7A/bmF2Bh1zdC9VqjUhQeJjARhOgdmCeut8lrm/I
UmnSbRwVx89m5D/A1jUiqzRzFAkc/tpBvnop1ewdVWGoVcuvmPTcdq+85cIR6DfRO8o9/uCcWfe/
/8X+VYxG9bMahSZ/n8HGoXOB2BNM4US4DzgA04CXNn1a0K/VqAE0tQdtgKo0n5RXVemfst4JDNO1
a11WZVOo5UQ6cnfK73YrpELsv6jwP7MIrBswsSqJjZcZps5CRWnO9oZSh9vo2CU2Nv47qyd/pRB8
UcW36QuV7bzCJdAZpxdSLKshfy/noJsvLnGDeakj7/wHfqOn99Jlh4zUHEFHXkyUNyocKeJOPW2G
iOUcVNvWV929yBKN806U5l5JUB2PLsVaRlWBh2TIREoLCLeFRWYt+zXKvDH24GzLRzxjTT+n1Re/
OkxY5G6ZXafGc+PmfWZc0N38LTuaC4s9q2UohLEPbIjTkNJUjwHY9P5eHUVEX0hdsp8Nd3gEtP8X
ylfGMeVTFviRjeQvs16K4gkr1HD7a1vr+Q/h8FDMq1b/6kJ5nWdvIjkNuwt3jby5vMd0Q3IGGMl8
TC3PQMqF4fwDy4125SGYFgMONq28Gvvz3iWRLFkXhCmao8YKMPywb/QtEASQp/eEFLMcOMnu3Emx
JQxw90roAq5iB8T5hyPPh1eyWMIkK4QdORllkvxNKOC9qWryGazRhLzjelZDasI4Bal3uDW00X7B
O8bg3z+5NTf/sfmW1mmRNAzJdwZwmBKsDFWEkN5VtONEKXaTJ9fQk99XNBkpvPzHaHbiPe3Obj0J
K+WPqeHIuR22EIIm1Sb3OGXbqsrHZdLNovHtCXtdlrh9OAkX4971gjUjXHezq97OLiFlQEKUOPXS
QcSn+CdYidMF9ri6GnvzGMIEp0got2hitWsTZzXldgcR1Ya/xUBRFXR/x0kRl+MlGIVTKME1LUjS
nmgyKbEN6pHliLhwxZYBN+yYRpGQrh8yqz9mz6JvTLDE8d72jiSwQM5RwAqzFPpbmRAasY/O2/Qm
2nobpxYTKXrVgS0spEpeiILMClxV+iJV6OXE5md+f/hcQceP3/8nS73oi3gJiSr/DAeW93pca8jl
oUDggf/7zEA2LYQF2UuKXEG19SJXbwADYjke009BOISo3BOF1bSwSWmTdOMjDl2t1scKD8HevHp/
KZWJGMbOkDwC1mffHBnBZ5IKH68fFOrNESvoZXxuoDs2NRRAm0NGdIrrj/i6jHD7QRV4L0mBQyKi
+BMGxDsIbvD5f47fLNnpa5R2j+CVpAg/OCrPEio8B2u84aWowcCHGaWZUjR2djbtPsSD2XhkjAtk
TVo0hL3D3Q0oCrnNKHclBYvyY6CfzW2lOxnI+gXkhra+aw81a7+Yn5wYemlAonsKlhx3KUpUYze9
DHFiZSEagZlIIV6vi24S/g5w7k81NOwH4GvBeUUaloZMqfILYmeXYuS6vniBFQcmtSQ8+bfyeqpd
QqH3W0yrlsPvch9KrJ2tpGHdp8waIXgPzag4Mzez+Zi2wRqnUBK/GDJI2ZhAjFac/2tQFj1Neevl
dLAl2o0kZthQgQ+ThE3QhuO4mc/hTaEXS+hhZffqbriLoDt/fbSNdMzu41xcWtOdgrdQnZ74WPiu
XEEOkb13x0LnRlGorDwiCiySG7oCLnGZ2P0ww0EwaEKDLNKZ9s0OQTnISNAX2cFkPpqw2O8gbF2X
U5iwLJKTPRbmhaOA3rOo3X2bonbDQQ6qDaUlQjdxOHPlbRGKl41VTihdsHpYKja78NxsIeVA8M3/
+N/yeR31BdwZxJZdb7cXJs9Zw4exLXF2v4ONiDWb3AhI5S2fYK9SySAop9+z0DJyfXAjpe8pvWug
wt8rGxYdRGoCcmD9bs+isXDHsFU6VJMtTHut4Eb8ZURDxdVPVzD/x2fiE62CAvforzv8dzcnZ1W/
+Nhm3QDSLePE7O2ie8gnelXCvYRLW+ZNvGixzqOIy2MO71aWxwGqR4TpU7eEy1R0Kz9cC8y7MbJM
4+QtBqKJ2xU3vgY+p0apUIs5lvKC28X5ofaNvWUU+8TwCcbirwBZAtTZEhlgnIlLW3w0Mc89tDyP
VNqTo9LwQ8r8n0mSlr2E2qK4+sBGV203AZZX+IXgzzRPd/bGFm6IVpq8hi20B5STU3H94kyyRY4K
/rTQ7Omb9Q+FazcZZL4lBWW3v/3oXwS4VN83Bwq4eu/ydP11b5aQMCi703ycawR0bgIjrjkl8KeZ
0ZKe2b7GvtHRGKaar5PFAWm1edJTwE7xVBcH7wiHWxpPLYRnZFPQ5g7wrxB7VEg72OJSL25GQ0LC
XhBgas/OKhqs0kiOcGbKEx/f+w1XjYy0eM6+gEiDXZedlo+BcU6z+f/x4o34+alaYaH+X2PfnQx6
9u1uS7j1uiQAh3ThdAq4+eVKTZ+hl4PFJgsjpKn+Zb/LPsFpyBqiq4E55y8keaHEfPn85ODOcGLy
lOswI436TgtXhkjh0NBGw1wWBfgjCm72/p6bUhn8VAC++KmFT3CaQqOgB8K/1PywPAfBKJkqlbRZ
fuUNd1oU9bHrHXVPT6q+Lk4sSIlwHD/uLNI32w/LUOjCQAEQZPLCadxIlbF7dfJ+nnJUfm6gAwPE
MoPoZBn1dfCv/3Oy3HbpZVrVPvj7NviGX+BMzR1r+wH4li4RXXlhxipGstDEk5GE/mq5JlYkq0o3
yfF1icWunxNG6idshAX7/6JwoOuQAba1Byg8O5+PK7CZqWEPunaY/HwOL0nFit5wiW8Gk+LGZszU
ztojA8L7IcjT8h3SBL3ZDmM15giodSNhcOmYLvQnMqbXUoTuasXGh6Ss3NUvRoCuHXCLR5nE5BeS
BJLw5H6joM7Mb0xuBPudm2C4ubO47tdzzokNhQPHQKWlQYew50x+TiEzP3ZD+eoh0ZSEsw+hVjnG
O2Y0ZMqBIkD/qzSjByjhIztqnbaJxitIGJHZc9tUjP6TFY6x0hrQVm+TjXyGTeEpzFluEWd7dvCY
jnDgdsBlYkZBVvpw6tvfpSvZ3f8xhG87Bi/zuk9yF/Fga8FFSbLevpcLtvFnwfOr3zRS+mOQpu1t
8ONl9oaTyLGltI+rbpZyMPAx0DeLZdZvjs6bRlr63ZLrck+brXjgcHJN3aDjzSB+3OSaujVBEQLc
vv70vCqgVkeVevK0jbOrqAIqlP7ISDL5q+x1WGblXY8CXIzxlmb/SD5TD9yGGpaI9u1jyzVW/u9y
djSlJyqqfLyDcavnI9i83DB6y8ISuNNGVZUOTIlW52hJbJ2/8DqH55NWDxsusQAFGi4VPGQDyBPe
Xy8ndfWU3LB2jjh5fYAQ8Vubrr7ow2zo+0RK+Gep4Lg9H6J4oOjFeFDMIc11jdyVx2WdgCIikQ89
FkTE+XTQVeuCiKv4mr50mRBDg+zNOZ3t265VkI5tdVoXjGxrSyeIql2FafzZib0L4yzmscJc/6Ye
wUrqU92t49jlJG66y+BXajTmIQxUXQJMcfmcnMQVyBrYyp7wa7cInzhkzudOrn2b9iVhSmr8Xaph
nwfr5PCgmdFlCzrQ2v9TW7D5rnETr4ygJB27cxFwh+BQ0SgAFeDQBef0hQjN2PaZRna++fA3MV0a
TmuFQPdqoa5Y+Qp9xDhvaXznCdIy39+QBJt6Iioh0ZXJ4sA1lDEFzC5WuYvnqTzFfZHLxPDs50W9
4YEyGA9TRRbm0N4xhtgLkXVXDUK9/wSh5t7/YNzXw+RqWxBU05HFAU6EN8pr68ykjDh/DIzO4D41
SKwosJTIXal//bQqXAizDkoMu3Qwmer9OjGknif00A+eWTNPJw+KxX3hdN+Jtfri9LxbT7LpqNyU
dr2/kJHSjtN0eg+fTwrXbD+hZaD8RHnvuP4wj8gw5NGYK+WvjqpLixfDZG/uVsP7aSVa81gMT/a3
BZZqVw8/wxJZobnJ4fRWSXNWh4sNRV0WeE629fpYD8ofFHBCZ41ImiShQnEnB69K/Z7jovNzk+DF
JWa0xJgR225bll+heoS9MC1EPGC1QqTOekoVtsWUXL8PwBpgJ2T3V6chgtj7N0Y+C8yoeBRYty3+
m6rK+5Z9z4+1zuhd5KKsMyIidzTJ1MrhkioAy/3mjUYdT5kd5Gai7hG9yJmAnvxK4+5y8pzOG1L5
3tsdbE/Iua+L62eNKL9hFz7jgsdD8RaqO/Q4qrCwx5cQ3TyS6KMRpwbzD4T8TFMlZRVu8716XiQ7
733u7akuntjgcgnScjlRYsrbH50vyVpzQlKLNKX4+1CCIpemeAXaf/N5zDYKvDgMeDY37QFuqzJC
hPH/JHCZSEat+1Px42sar7Ve8Dz1euo+YOrCm9vtJyEpvA2aHbImdAPRtbWdyS9wl0rNYvGQGxCs
CjfNkFcpi0y6RSVl/uSvXSN0X8uYbUPfpGWhaVjCC8py07OeQcVG2E1dHLrDfWLBnSI0JRNrfAB/
Nq90pqRuaK+K2WEVtIlBXj7jTWMAeb206xq+QGbfQXbNikPB4pRTzL+7m8oUwC8F8bgggUo3pZBv
Sa7YMbaIHgk+dGsaITZGGlMhR272XePtVKTmb9/lsIdhohRC5b5atr3sPtSJv8qJHq0auNg0oaPv
KZQShlkEM8no+vVapDyDp0G4gPTjugjwfiuuCo9pjXHyb9NXZinHZozxBeL+2f3w94ckaE5WSGF3
EQgq5W7myIlTpVM4l92R+oG5gONvZtnf37QJfpBc5RDRDLZmQmT2wg0gx5g0s4S5DIVXmsASRtVG
Z3nDPzmmMjWMh+zwSyFZDv8g2cBSRWFSyTj4ED/FEfVSKp7OeUMcL5bwFhScgDVY6K9GHHexrGcL
m1kZM6r19vbKSONN0aTVEJQuVmgt35siAKOZRerjW5LJDsPpUVSP4nL3E0CbMf15fZa7SaVqDzSE
Acn4tJCln0WyokyhDjhq4WZLP7CIOo9eXp0fivAvA5LXQez3BT+ThMC6H2aXhCXD9krA+4q9cIL/
9Ewj49uCI35fd5FB9OXwB+GuWTSqjPMmo48z7/EesCvGRMGaVW7issXxbpZH9FWg21Eh7iBYLrEE
8exRe42IYgs9EnH57K4w3N6ek4vsOIxv9DhP7cqSnmNlOdQIzLliG2zuiz8uSjNzxSJsC2GAjkmc
OD5GfkH7+5d3CUWAWzm9qH3z6WfAE4a+x2HiBXGAGIQujkMRroLIut4KCAPqU/2wRVnhwMddDWt/
MUUXXizrYeeer8BcAm1y2kUPEjo06gpi3LSj2aeVkI4zq7tQBfanKhI0K1vYuOeipxI8OLdpvZIf
ojwjQdSnhPwKDzlZqNOY3DJcnS9Fiv07AXvgyQGOaRdg4/aJ8Yxh8hYvDCf11GtRtsgoh+vQmcmf
8oVhk5tATdwwU+3GPBSs6UgFgcFumiHK1jE6jbM668xgAQYgkVYAeVuzytICxqgMEPboAoPeAmxg
i3Rb7ToINp16XFWhFa7aWuJ+W6qm7qPO297G7lNolB1niZhwybqz+YpNA2ufKI7M8gMUFBqOpW/S
INOTJ9eoRv7UblFNTB2IE8RHtOxTJ4DMjADDU1Dh691wzZF2t4QX607+cdsMAUj+4v9LLEfKahEM
DJh+puW2oHQBnBCuHNeRtRazlYLaWdzbwNAd9M/O/PvY/sMK7lLyUwzQrfNlxac8/aHF5aeJlyh4
C1Eqk7mu6nps64osJFWPfhb+dQhLmyCR9FajQahIhYj1pLPkGQO5k9gy1NYEhVorxKXLROcno7OU
Bu7q2M4QlT9ObfLA4NvLJLfpPHwLlkeLIJKeUm13cTiKpgYQCBqG6Wxbg1CwLmthWBvNMi3Uvz7d
hvqCViW9706sryKHJ96nhzgHCRVvvIBP/NAlNmCYDpooNkrmXhw16shXfsAZgqxWK7RUWYzVUli+
Cr2kjnQr1/MGCY1B2SKpVz3pBEzV+yZHcBRGPx319jFM9UUH7dhT2YE+3AFdFUYasLgG8ItOAcI4
LIWdJxqnlEge0jwLf6yxa+bO0zOQLVVRCXjviLa5Aey1gHV+fsL2Fl0GLOlhD9W6dLnKi1vp94Yn
XYnFDThYARSXuu5nssVee16gQ2oMKkToUzPkhaju4pUlKT0IBM8EZrR0d0uH3OIzhtvTBoPYxb/y
VgYJirwXJZAI3mBrQJDE9v0PBeJ+iE9IWzvRNp0CUjodLHQmK5tjE+T17rHA0etU0CAtFUVFnK6m
GQeqNwcz1R76o414a2oLa2aoWJbbagzBhJRKx3WRTUqav9AbPZ3rb1F3bltEQgcl3STfzB9FtLr7
FE4zAdpdZ3lT1rSUliQyG+MEeUvP8rEaAT3JWdYlZxbf14naW60Qcuv8Ykb7mKeplygaubhD/Xgg
pfyqprGfe+jlDRzSbZbAFFkYbJBO2lzILekZSh11/u2IX3YckToxGo2/idXJM8F4y6OFOkSB6Rud
j5CZLmCr3C9cHb7lnuG0oH/JV6T+38ZjgORbuc++AQsXp8D3qY52d67vmapxGmNjx9800JPnqN55
j1vspJwZRLduJrFKp8QMSQ5q6eUbNwkG+SO1+ceE6auP8g5oyYSz9eubP2VW3lqUkSiIuC915vOy
TPX+nwzMLUdP4Xq4MqoKi/9P8gpxwtvMIgaROnMLd8qyb/ToVedPOCC61fPeXgDBPtBrbjG2Jxrh
i/Kg993XeDTcyDkIl4H58VqXEw9q/oO92gcgFSODY6s99rMADE1Yj9K0KjJVwdCAEwTjBhBa2lYC
N5mAhPeIGHPCo5Sq8yAf0F7qryoOapn6x3LqpeTgyiMQoZi6v+Lk2vS3R45wLMGaS6bMipMjoIub
o1BINP0xm3f/PbOcx9eU4P7dG7xdEOVbcvtqNGU6B1CroyqpLQEqZeE89g2bIQV2b7jPSbIacFAY
4MsNhRE97ihkC6WHSPdUBaEfg6e8rQFpULENZHyOa3oJtAy789Jt/YYj7S+by7og9JReBSgvS6Tk
+QS+i/PIC/NfpnOdloEoITquSO7PhoMdwq9lHEBf4YK3U9SxuLDHZPdHusmniGWKvH+9R8ZKumnm
IUHzD7/X9cBsb+VTuebDQZhydvgKKfldkJrDpB30g3Eleau0bNAIirMlQccb1e14YLOkKUJ66I9l
FLvNRLQVXIzNKdSkjc2oGZHdSqmdp2c2fnhaHWj2AiIgHSjJdgOyl637zktDlWM5FNS70wjYkVQv
ckZ2qLPPwL7iODy8y8n78ils/UJ0HP4QOPfJX4kgxfevWa7JN7O5IQ+Atv9kyebgymAh0VbD7PAq
4M7LaHzvdVfU0fwDPJUr/5fKfjO1reWc1bDQuo8fVJgwUOkSvBwLL3wPDdBFYgM1TDV8j6rel5TN
lEOVa2zOeoWUzEVUmtRZEjzFU01xLGSEvbXS/0LGuwfS+jFhP7l53UiUj2exuJyc5dOC5bBfdEiH
UF/5K7GIcS6DlHj2dhKe33g5B3XrPdzNpWZZ7L31x5GY8qKkmsW1F7YLutfJyDFctSCKEWfBYTfm
/paaKUSJZHAQXqnWpC2R0xszLY5BhUgCXICu6hi35p6+OemeTaery5eEijXad2tXXqyaKbu2Tve0
qDBizikIRH5DziRuh+/n5/Sigqr1DNMiLaN0jittGfeJCpIYiDotzTqoMtQzo2VJd+hUfw2P13fE
shQRNtkIeYyGFPK3iy/IWjZ+6JIIuwLSKJKwtaI163qFeU4wCVkJQZSQiIyXNnspJhtrOLbQ1Ubd
e/UWp3jjD92iV4MOnOIipgKT+strER5LunHQLfZ8Ff+OU+ylFmmX4BQooiPcqRHs3VjjVPWmxB+/
LJS0HjiU8HMD+Y8+wszmkIYJEI10KuURiiO3A67r0M2yMrwEHHbN8VbEdahU8DLv7wMRm9kWo8sV
uQewMsYUF4oUFTbcnDqZB3Rvi/ibIQF7vtP55r9R3W9LTDVIcyxt3Mtho8Cqx7P+7NoJ+J+WYYI0
mJFPl0ZYSsApvfdLDLMpogM0fhnwx+tEFx6+XKsyv8ie7RIJ/L0Cvli3x/I+PeeAGuVmW6DRNptQ
9R9/m6+PzdXNc20gFqYgoN5ipF9OTa+HUBvg3yfZlswYHJ/ASTCgV6lpbsHllcXkJdD0o8Knrm0P
M/fVFvT/4GDljpZneSV1ldlRJ1658W4Co8xB9ZgwG3O7J1x6BJLKCzR6XrmH9sNqnWjx93mwnyIA
tV9sI6aEFaymm8/HKXMQSRYAU4m/PJfh3Cn/7W8HlXd05x4CJ5a58f21rvBUBBJwb+j48OkzkAp/
Iu+ozyv56PuIaKKjjah/1GQENlZpMablZD19DURSQcY7wR3F/f3YF5mNcAAEp8HqdukabsEforrw
zkMHN+seJxnIxUhtZXfZ0YWBGho/l8xf4+W7pxExBEuw36eb5orR3LuYerbHug9CAV6LfCqiPYkm
zaFclD/FQimc9Xf4dvDyI0AI+SEr8Y7GwKw2EPseZ4D/R+A1lVHLnXa9r/Zhn4U15mlYxI6p8BEk
aGhJB3r4cYqniBC9gqI0s1c88PfCwz8UnkJUktEZor0VZrhkJcBUCFtbCAf/3u+WDrVLdCK3NKii
C0Rq6746NGAl9ZwmG3e4xrDMFYm4qlglvoZdoNXBivbYivHzYk47z9z26cM4cQx7q09662352WHA
beaxBnyJhjGXtur86/wwRvHBCMfWOZfWgdlz1LnqxN5gm6yyfZQPTYGqZOJi+FMO3YBuj+01mtDK
vJN/dVLpuqfubmH9dbQOSy1Btfir7Wu5xket4Zh0/yVZW0R5L9yvHUCd+8JdYLxTiynX3KgAczpr
wdloOi/vs8sVYVhsxeErmqwp0tsZNxTnFp1MBso2CKv7rQWERz044YyQkhwL50Q3eQOWTFcbxAYG
TIUALNC3s+x6ysnXxuV1s2z/o5VEduKL9xsfvLiYVftEv8SKPz18VOEGIynTb6ePwLB7BccaeaRd
TUvlbEev+DeYZToynF0s6lk6bGKdgdF6HxzOFU9/ir7cOXBv/NHsdcrYR3ZgRoJm7Vc6L2nvCx6E
zcTigXMwXjJOgoN/RmMfdpf/Ev4JUS5oNOpWSVl6lXPOpZ4mbxZqpMC5gsjXkMGY1XvfOns5/hch
SVbQlKVPUhQpLTe2xNymVvMlvwQos5mJSniXD4vFXBYg0Zo7OOwCf6GGLFyR7hU5JjaOU/We5oXB
WSYOxjBKUYMQif9A4RYDyu2lW+WqYlitkSN7V0jJd9FAyUDlHSSsZ8UHHmMKR40sp/bNQOdhhQvI
FsggS8CnWuIDzPG+BAlXHM1JGHo29aMtpocPFIhseLb4EmbW8+ef957DnMVEpQtXGcsBjHD+s9w2
cexiI5jYr81r9PaKl4DkzUv3/xl1VlvqmIYMW5P73bpvz6QXayE2MiPjMOtrKIFTZoiOLKifu9w+
AyUjLPsgN/O/1VmbdDVqSSvs8qjPdBFSjzwXaXfuxEi/aFnXQRkGG7KeyU+VfdmkqzSEFgtWy+8Z
8pbIpeWiYJAQlr8G9qfLHNDew8RGxXOtOgM4R08yFRplBA+/4E881WghMcXtbEEk7hUGkh0sj3/w
7Et5UKsakHxz92eoynj8B0ZdfrEzyhoATz1PGWDb7j/OF1+qVvT8BQ8nFhD1KB1Cck2nLnlgAx8M
mJuQZVJU4bpDr0wmtfqGUH0r/b6VI+ceu9U+CfSLk9R/ziImurFaxJ07uFr0FETRkXsmchn6jj8S
g4LwWX7rN+sjZaR5u+KbYeJcpuFFh21GiooL4Oo17Q0CUSsFuGK7ES2VZWP1bpCYrzl4qSnFtCwG
YpE6XDWxR3aKhDTcru5l4DUfON4Nh7I9GT0nEbJ01MPoQfKUEZVwNOjAg6RcDFb0x/YGJBgIMk6m
AwfhdyJD67bwRl3/1j5KigVHL1AwSXoGJGYdX6nOjMprxG/YN83m3QkMnvRiPxxgEAYkPmIVfB7l
t2LfMoVtuPfDoWxL5G58Zn7PIJ7Sm5GZq0HMCBWrQevXvgFf5LQ0P5hQv7hKlQtu0HZKcxqh6OuR
9Of2GNrIttR4Jmf955C50f+LZJkL3rPDw3wwyNFyqcKBZ0L/UnqjYSz3av8IEnSwULCO4EcZOSf+
VArfZseBNtn7236nSaexkoDk9R4FmBVdqQ9F4GNM/3/UOTqbrX7dAADYy5zOi20mXWZwoTXl2pc7
Sgq9rfKfjyMhiODxfOJVRgmo6Qz6C9d68/gh6sHK+ymc/uVwi2WrE+kqyG8GIdlBiwMSWBHsZiuo
2+KWDXSim0qAnq4cmGIDco2KFz1V8BB9YqqDT8+EEDSE4Y3d9C/CgHC0wiDtaTaLnoLZh7lZ1/dQ
rJoSVe7DK2kCRQfgBDgNxhPDLL0LO0He48xrbkDbvLa8gTHlKTyU8PMCiUpvAnp1t8aEiXhLSoNS
bNrPNuoyYSu70s10yStV943GuhfLz9yAT0prlO1GLgaf19RajZ8ybA0o8R/h80muNcEWlmxKrNZb
O/0a14z+AfwaRFIG4JNSH/kENO2k4eJq1qBIsCqhiYYbv8j7Uv0DqI/Yig2ZwXNc8GHeB+OhMlRo
gchFCqjzfbDwbGc60h/wy7xTf5knDuh4vqAT1KP0sBZlc/mOES7xs4Po8siYybDKcBuEVl/l2MxC
UvIElQC5jm8cprdnpGvZKHZ0ij6vMDv2xNtlWKq7OykUPuPz3o5FCpLY55VogN9YxYH9S2V4R1Rc
fGgwD60haSYeXdgEnqcoyIf+cBVZnv7HXAKJ6kMqIIRLp68Hhb+iczwPrjMIIjOs36qzTKWF91SY
C6t23FixIMdjHsG6Cm80PA69II4Zi+Oo9Cnde1+UiIOSJBh4f8fzZQAO6AlF+AhCPhI3OSegNn+I
VPdAisp+yTDkgFthGJdeOxNkX1BLCXABwo3OxxKnt9lCMZh4KyyS9JL2bdDAOP0fnd2UAYwZcqlt
ddN0xAGz4/CB46E3xL6kDmu8kYWPqqtS4ts4JlXI3qrEv2QmcWPxCEBWzB+lkXm4eGwWY+9XUCxC
V4lAL/3jgwfdeCFQZfTKU8E5kj78XJmuvlZiSb1JmJUFePl+838gt6NUd56bbmSua6UfAgTyn01x
fnIWhIZnSOgl1FZLYZVUZH0mKACtsKGhxCey7BkCoubtFZ046MKa8XVZ6shUZXYztSJ7BCXQ6f3t
KRfSQAxy9xwVNLDVdg29gzcWcONcUV/8Yb1FYFzpncP2Etw75HTHu0qW3MjOjeP6RlMMrDXaRxji
SoArBwXC11Dj38A8r/h8yy+qv6K8b+XhVhJcDVt9evPeT4JbAdT8b22R92zvlWy/MA4muFnq03+Z
X71P/S5yzFHxzrQcwIPnqWBZPMGQRKgVZATmukH59ejTHHvODejx6vCcZYE2AYXTXrJdoZEpTnVb
dpFkrLClMtFKrHJawMrVjeX91OE7HaszWt0eYT4/aoxkHHfZBBDdKCtKevKdC3qFA/82F1GPBmib
1dPLP/3sN/vmK5e2PY8hxoJdrGfBoj7D8nuPb2UbezeUE5YW6UVcWWy8Ye0pQ4sEoE8TJwXLJ6G0
npvWn16x0EkaMe8U5UjSEFRBfe2u9BbCibgoYMmL99SVL84LeQ+G9ScKmPQ8cO1wNkDKEZ4a5gdj
UbanIE4/cvTdqzvtTmvR4VYAARY3YdMtXtB4kdvp5qENF3oBbZBo7FGz+O1Zt6iM9o+LK2qqlgEh
OdLgxfnQntKTKlqRSqZ26iFHTEOLoLROn91V+b55SGY2Ptni3zwYT8V+JyGWDbFWPdgQMP0hvpah
VQxfpoAafS4TyCdVLEZqkM05kRGFzHuy2R77Exilt9DLTGTHISAcmxoxms9ntoXQwKdaIRaZ5vlc
AjUsl0Tz69Mw+wzWJK0/LD2pAHdPEmASB4pgZ1EPKpJY6nv85DOe5vk3gIAxdF7+kaCXjGmdRLl7
8fNKu21QpR1COb7QN05B6Htj3Oh30W+3CC1ZCV3on6Z3RDQLgMluvgXLo0FSpXA8B+fvZfkMY7BC
xNmpsWqHE34B13OKFDIomrNdp19ZLffe74Xr9RUMnpnSWQNklYVH9XbdoioGfVDKFlzUIeJNSbKP
MGODN3lBZxdFeECvJ/jymLdEeIt9lCS5AhLIAWR5RIlcPEwDs5fWEhsx8gq1uuz3i2LMIPWqio7E
XBf76hV65HDEMTd1tPoJPmfsS8pVqZs0qtEQ6oEVN3XciFeZHrQnLXfd0D3L7lUI5bIXnKy9cTie
twR7bn3SEFhIGaHvM9sRQpBPk/t9Cl94fdj03aAGrWIGyg+qRFl80HqeZ2tXRQjxM4zHoV6f3yZt
Wx93nKieqm5GerRvt0BsmHCOhdMXCtuCagM9MbyhHu6xrxuU2Q5r/zk79TQO5KTOFeCDdUt2NDmV
3kXGXOFW91dGkGdL6bp6FXuFNUrTzGEw9tOurUrEKGdkaQV1n7tbFZS90hjdYanXwsdRrQFhE0zr
bqiEGx/2owB/ZeozRWiqggtm/0oMz6mec6GfmKXYjXwD8o9qc2jiOP+e3DGSaFTKCeazJOO0Yc1f
HyBzi1dSyA//1Io1bdaGo8WLVO72JWyB8CxgKHf1aKejXhSFr70zj/MnrT38qA7q19daEZLgn4cA
jgrnriYuvCV4cqiWJoBlglyhkvF0nn3GsdJFKFZLAolptohR8qNLPaoZsMK7/uFgyUxbkYBFRcQO
mpxPVZA4PPPuOeTYl7GhFLtBsJ7imOIf3O9cWpOKuOBx52Kt3lqpz9Kp0dcGA6PDIGG7KV5inkJp
3l7TZWna3t1UFQmZP8DVHXlQSlRMFRH1f8r89csd8xiVDWwcwlAWzn4JK2HcF0ur+tcJahgsyvVY
M8ldFLKjTndcQI2WofNG8f4kidEnh1TsTM/XfNSXAuZc1QSZaLsE3I23guYlbWg4jD1xlFTRnLTV
gPbpvYNeyyVZdbAoeoOzqihbmpTyBOt84ntPJAETcZPxaKA319o3bCCMz3AfyxnlJnHDtyiW2eEH
7vXXhpH0U1AWLELYsdCIn7clueB8HfYf4brzd5KSwWSp24zqRWy7tDgw4YolaPsOSjoBbFnaz+bb
3Vy1Tjm8VXAWdplDKb0K78TIhi8fuh32RejpbOzdYMD7Sms/G+ezRQPN1trV0GfBuYK4nk5BvnNX
xeV5n5QclrsEx/8chVevZoPGEjOUCKFJXdLEEw+Vm5o1tgKXK8mmQxKftShTp/qKXojD6WpmXgl8
rywjceqERU+gjbRw4YT1pxCKY1W7SJaPXZe5M37TRUDkYrh33Fe3TC4NEtO8jgoMu050vQFVPPLy
jn2Puhm2U3z3LqEEyPNoEttpXwlTvZuZHuL/NH17XjTUkFAMi08Mm5SzuRprkrbTQAFGi8hFN2r9
NiDY4UjGXiJQg8QY/jqFYNsnSEpgdjSX7tgfysxecEOwwM3qm+nMSOjQFOO37zBsoj6ZctVulQKB
xnFfeHdPWyd7TfeXpElU5HcGlF/duoYdHoIUEy7fu7wldWG7URPmlfAif4OmVstdrKVXPJQ8Rvpx
zf86Pye8Teu3cQ7nvgeLIUKCkZBvrGURkxrvcxdkj2zJMc+GmHhQy6M0yigkVAolm+7PP+xf3piu
TuJFbEyGcdan2BnRzqFZoSiuP73oa++jNSA4JFmdslTeg7rXpfDHpwV7AP+Aa253nVZvhEz/FSVN
BrqM+Se1DBIPyXgSVxYjwrY3voN9BVCA9tWXvYpMsoeFnnzctCL7d3XYUn7Uj3jVKmHj9IOTrRt8
3GAKWPPOgC8am4S9LVCc0QLl3BTf70XbLJZe6HUVwSw3SmtaFpVw9ppAXqP1yYF9FKeohJSynyv1
/+N3aZ6dzEXwcKi23xpNYj0tMdcH3TwlEuTF+IlkU52RC9HyxE4Pi9XPADiIlZea8MgjWC1uq2Ll
xAxpDYR5w37zHJGeXAXC6H8dlJtGgLlC/asLgs9fto00gXXIzZidOkecCV56LcbOY3LIkED6OvLs
TL40zYgzqjZ3Bo0rj/cQ+S00nFBv9VvE2kOvTe5TwNlZ6Js3ckylsqi+tb0tEIYIhFS1V2lXorZn
HehW6rMY4024gsscld+VP4GnSDO7cQ5EYy6qT5EcZi/tSWRyjeeR1wjOhMz3JedRLZJKvOh16MtN
vk4vTZKFZN9ugu7A9l/UYDnLm65MqKtknDtm8Zv3oK4PQaL21LC+FEjAnikFxvpR2b/WWAogu/eD
9bArbOJGJFI3yvl+HepCiRPbG6efKiUMeHSCcOEK89r81ZvNtPPpklUTCN9DyvUmkFybeKd4EKY6
2ZgfE3BZcNWasD2RKIFdAGib4Pax8B57hM7xr5KbGonTMuHUsSazExH6KHtnQLSctQx8fZ+tNowk
E5lCXhX00xz4Mmfq3iCFLfrlUyNgnOE5D/8TKi3PxZ6iZYtAO3MXspiuA9X+tZGXrK6p13A+V7l1
TcQyAK3rneHTNkZtLyfIv9Gy1QMcybFencNd8j2WfDMEC3MPyvnMftG4HNoy/CasN2cAORYnor64
g7PLktymsqwu4VlkG79ztL/bUoaTFDdPc6f5kAD+UhznDdeCOOgkYzAuXk+5pVxUt63ZhcUnmEjF
cp/SAvyQDuYVIqvbxxkuz/6gy9iZmHvGa3YVgz+TOjig0K6nsPa/Rn/wtQ6WoaWdb8t5HAdAB+Ch
eDWs3FBF98k568MDVlEIXvOWNjRUN/0TCb04TgJb+WlYUfaucXtCIyqj3IlIBg2LcTHc3Je58gKQ
PNxLPvvYaUYXnW+mkbWAhwG7V7MJ0XvWpeuHJwFS1ravLTQopsAwT0fGZWAKoQrYMXPVvP8WuOEQ
iFxWoGnW/XiX4zo7aF4RlDwyajDLr1VhHm0tNH0ehIbBgPHKJ+qx90jpmO92m3Tt2+g7t7pUbTAj
rATHP2ivqdHeRcjrYAsgkDbsD3CbUh1WBZRNWsCU1uCI1++6/BEyMFNN3KYMOnB53iZKmWO76gk4
SwumZgC196t1XL5xaSsxEOmRosWf1TrLrrFJZrW36YeEbAYiO8UxT8sVGJT9YF2HbTenOhJrVsYR
limA6b0JUcvRh1NqiL4amsSR8V4h5HoQDlx65zOwyVdLOvWNGPsu9kH4w9mNn6b0eglRxa5O+eAw
B8jmbATNobqnBD87CC+H4T619WeqfBrE92oMeM4tecuXXAHsqALnNX5doQPNU5K2ncg/Z7MEpl7G
CrJ88nJxlWvKsaJUxTMjDOQWO27j68V02EMCzwGWWqEAt7Bs1KfTxxJdOM9dY8E1S1ocPH/xESln
AiVTz8Uj9zy8OOO1KkOH6Llo9PXyGez5BTw92cDDgsYgUnfLLmJBUY9l2Wm61PPnkUm6fklX6A+4
Vm7J+zPHL7EVmI+8iOXvhjrEurrgALVLTMWi9mZYq9tG/VARLWqRDscwjzkvPq6hh9IAFjTS2gLU
12TUp2OZskORN/zPiQ9+ALj8EfZnzG5NjTfOWqdUAsJeXVemWbla7Efiy7Xyyl0maCqRSfTyjfH9
IEwAHxZVrxF4bCCBr7iKEW9BcN1v4WyPHFXJHaQW3pw4/bMAce0RS/6w0s8S9Khz0+fSeBXmvy1Z
fyDEFoqlcSfTPnwyPpTNGf1RyrBjRgbver7rT+aSRpeokIAHGdHKF3+3Ly1dHAvzHDz7orX0lNrA
hqpDLhKmlzv7fbk/laGjuIT5fpT5t6SjvLADmI4Jz/xbwyv3tFZ0rxUBCBngJydXbmeBrYFpcE+7
nWjSl7uAvSRDvsFGt8Wb1XHdx5CMJ57ulKPmwdA5UOrUycjuHVVwKOcgzn3oZai9z0/YEngg10m0
mmdZ4Euz1oC/+Wr3csQkDDXeg7+CcTk4QmQoqZpfcUy7fl02xqrsQpIzZX8ZndHeBByv86tFzwFO
lU4CSB1VA+XPYidNy8HACXlZ0TkQtel7h80UetM5y9P1gaL9cAsEf/X5KouHei8LQ4s6andGX80/
WkxrHvKzVCLnPTSm978sUEaq8HrzrqmT/JDOK818SQkWK17/IrckNSgCXoGJ7BHz2vQEfZKoYWBU
tKjgBbzI9FnIR9MDhNDNpLXDyjh0H86MFZH7aS7VSGP9GOYR9V3FRsHmqJB061N+pklakf+bX4/3
8v3KUebIrMDThRiq7QDVE5UremU2C96I6oZFpYrMgsmHjtFBoKfv4MefxdTZ7nxBri62r8+WVddB
1E8H7MuVw+4LNZOMDbP/CX6YouzVna6OqaeRLf53WwzDNccNq0a+5HLGqhP1gIJgqu+exmIG9cr0
pHCk/0meC5iZkQVdJ1HANQPGullg8sEyBrPEiT8zJvpWBfdUjKd/GuEO9R1oT2jbkTagVobZ0+Sc
nJh5vrnMvkkwkn1cCLj6LfWiTH+8VwCtPNtSjJir3Pg49ESC3rPECBiTUawrbj0jR/sRAC2N5qcn
KqPT5S20i0lSURznjD1RoxIiJNBZiNWWmjwcxvkaHcfDtKxDPmG2VnhcVEaOzKGpCEl1Me6sC9qg
94mrJrlsxgeo57nZxJzDQRuQjjmSKp19lXWXAC2ooVBZNv7PryLDnLzt/ZtpzT6bqjrsI8ro7/5J
HES82BTGbEExfJheGYNJu48QNJnhUxyr7yuq8udaGZmKlFobotaK1BxqRzvW+7PzNW350BdTfy0f
yW3zku+aFPuTyl+tjqt9SeFBUd4OLT0RiOHVwWRqvdjG2vHcdpPz/tGPTeaSV0o2xYSofF6SXsRr
P1UNmBX7G34isM7O6jfNPF81kJgUkG3zC5zQULnws8JqVMFhbjn4+tM+8dsqN0ttJyJ/Q+IgvBre
Cc5TBQPuljd174JW0InG5AdgQuYellmqdvH95WhO0Mr/BI2HP8hKKEC+7GEf1bXR/LHCZPIczGez
VvkMBSIG8X2iQnzyQeronYV9xAHaq7rrwFlq+7/kIB5GuffL7hlukn83yMHWr0t5RnRh/tkdj5oP
llQzeayVdwc8IEYw56B1ypDoqrXWTAnHtDvfdeS3HXQ4HbErF0DtI1050r/xlGnOltkrklfvZZL7
8g+ScsL21lXkrAI/mhWbavR7PYHMuBgyeLEtjbli4v9A+8g1kGGVBLoxnFod8iymvYSqgPBP9Btk
jM/KWG3b7UZZ04PNL4bS4Gi6jjQNk/ipnA4COtxs7fbZj++Eok6G2msg3W92SVFMao2qlTDyIMSI
S7P2Idvaf9vl394GPWu/nP7XaEkEX0CzqTGzRCXOflnM4bU7K8uNIOnLnMOR1BuV/W5lJGdfrEkN
cPkzO1wMjqzKLI0R9E4ItKLHk316NKBig2QPb9dmw9CXsLrqAW8tjqCe5sZHkoT4Ppt96LDp+8yA
FOX7toQDopPJoTs2l7uI0fYTqMNfwCmo8ghZi0yPeQbiOjJX64+V9hzYmgN1EBOLf0U9POkqz075
xl9daihbRdbY8f3pAxeIGjvFFOQWbWIwPed+NRGq9wRZmpDMHKE6HKwoE26Sz3rc3FiGVk0QplPu
2JtMmWSyymRppUlw5x/xDboFEd6FMpRvKjCl9Utuquyj09IJNQQYz14Q+IhlZHMlsU99dEfmE3Ac
IWObEhGCJbVBnvMjTcpfOMXdnoWxBT76C+acp3x6px/Jq5Fier7o0yzeMkYpL8L2bPS1OSYO0bx6
H9LpeHHMBWiu44heDhpsPO1K0rc8/S7a1n9TgOIisjfkVTGu9VVj/PIW9emJDBPnxoxvYaZuFihg
GiFb9DcTLUYPnQJ8dOZbR0tbqe26JhtNyB/WV4mhEqTfzqsxLQzIZ5upjnLj/CwznT6WUTkPz0av
aIHawtXGHdrUwOlLinMptrSln8ImD80WOpiYY+ZeFG9afburAry7joxLXX+cVN97Xx1Y5XvIpQ97
ziLLUOZ7MXTGFWCDmOofbHMf0mCVj/LyFoRs7cqvVUPAHTooG9R/l8Kb7XsemXNBK0JJJn8LOm4K
6q6ktisQVymfLdo/YjeFoqrGaxwV4n+J7XYrLHaLDAX3NI/mIe5gOSCFE2PdxSdHkUdG+X88+eh6
ihTarG5IHmongHamVkzPBC+YBOrGBMqi06qqmfJQLAkQ9bXdNYZZiQj4++mCYy8fIcFjuByVDtrc
T0Gv9U2eoQSuKmCS7AnulUo9IyqJxh8AdxAspaqMoPZi1lWGqhpj6zoQRkZ6ss9CKnvB6DqodBqQ
STSHp+dmW8jbVtSud/mkSqrPeFeBE7NFGDy2skPJ6ITU9wlCNV9NhoEjwGHWDjgtc6RlYp4Fo9HZ
8f5A+7Ec7l6IZtQX+qYaziaK/68S6xUe2WiQ98YgYFHA0aRbDJoop3V9KsJYWagxqN6SorCmeLKN
z8piIE1y5ACk7TLcyyvy1MZRHL/t0cI8j4sW+Tzh4JhEPNNZkZJH0yilDUqdyB1D1T8eyrj7mFSu
tzYCtOW0Rfi+a9k71UYwZoZFqWrW8yON3PxK/kRKpc4UhtK6LUKeZPstYuzh/lprL+4I45kGKzwL
suuBKWjAzmE0HpykLnNZDRbSAqryfJ6hRPiorasmGHS0rOj3h5nhtqhoyms0wU8+YnTgYbdxD5cW
h+Asxn8h4xPHLpk/RuTYbAciYniu9RBE1Ri8u9LyzSVgKKjtKur65/Hog4FAS866wnksnI7NnPAI
ydBsYEVLaheYFpcjZ2KeV4VBwiqKA74z5rJ42Li7S7kPDvzpRbMdyOincRh6xmbffiWOLVrMOlWi
lxfXiOyEYzTCFAuvZ3JLKQ2Mbmw2kXySl12klovGmW+4ZsjRvJUYziFOME477E4u1DCSuBg7yE0N
GKHfMmnXXe1gttDdJbfp2rUbDV9BA4YHYmFz1snEFdYjJzA9JN2JtPVyYnjJlDD8dg0Url5czt4+
5bZLbLFuLs2T93mC9ajgNd8tipcklUlFzmSvGiiC1N4ra35J1UH4LjS0cvwNxPW5GoLoZ7YuXbFH
oG48zBEDEtjLL7uLOxpvGFG5EZi1ICXSY28p2GaPyKaZCnWFPkUvCwajMogO3TDw35oXfdDMCv4n
r9m6pOXdFy905V1o0UdHpvz2+3manCJmP4FVKpInk7qAY0rZSvVhsHtMZvZLp0SpyrC0BfId9v8u
ndI6wu7+ycgI7NKkrCpb7qeMs9AprXaYe1PKRjjy0ov5JP80N6/KO5k2InnB7ikEg84MHHDP1+SE
/960zcxHYqAut7zOggwAn25J328ZHbBrjNVHJGQTcW++XzmZb5BNRigl9bffbFi7HcXB7Z1Xtnwv
0r3gjcdJjiOulPs7MKq40t2oycOs4CaisrOJrjEMdmLk1Q/ImZBhjJjszs8DxA9emab0c3v6j6/r
Gj9fA2Wnr/zfqye8MU1ruEBWJFg33XIW33t4GaXbUdo8azZJJJacoB3yRdWJnYx88rc61Uf1LxUq
gl9THkQKnpDTizlQA+JBV9GyZOc+us6VW37W9rE6asX/K2K1lcYzu1ClTRBXw/v2uYu4Y20LmIeG
bHFbMq7DJUj9YCRcMwxOoz0GK5QRFiutez6dIX+GQ3mOOCwWXw6ff+Z4cLLHUzLa0PJdqZFxKU0v
TK3SjJAuCa2rrvD6Hwaxg/wZfHSEuXBFY5PNNS7L+Cn5neyp4mRyRe3e85K+kg5DLzKQo++ThXlq
587YDJpbwlvStyzOr5rkbmLoHlhNmHHpnkC1VTLEcXlHkMiheVe1k3bdOSTQ8sFMl+12Tz3Q1N3x
2Rl+PfCmkN5ko3YKtjAv+I+9Yan/bZLi2owIBMBx31br2ddgjk4bFwzHICfy1UjJwRl2ZwZzUFDu
8nua03zrkOqnjXyXNnstkBNz2MV92TAmPCugv5KV85CHJw5aCLw7ZHNUXLHdcxYvYn+oR7HH3acd
L4W0szJULRfaGfuxJSiCgxu5M9jhtMzVQ24FihXS0EFCV/2/R/n1/N0sAuWJn4uxPozZ5EKyu1HM
K4eqIUE+b+Wx7cZ89+qoU1ntz97S0WhvKDzf/vxiLi7nkc6tccdXbbHITtT4PSHpZGdHuL2gcVu9
JyFhuzpqL6LiDwbip07abX83vkHbe71JlHygMrd75gYb5KqbpEQCTjXVDNOOaR8GdnPCjq39Em0N
Rb7CJcJB73pki+gyPAYt0XyjS43swEIsrSjTgIeokGP2VXA6PqGaBL6sxHfobZJ9Yws5XqCMxpCe
fo8yz5vch46kjGT1e/eIv8S6S4IbA4uH3W3odtzVZFIPTEyyKeIyvoH0DFYa7kjWGZsHWityteim
gaOeFh2uEpNUhPctj+6hJUwhFGXHD8JIueqJR+cj5wnJFZn/PSvMz9+uiPqooSYahgCsoyoSF3jg
PklDxVgc/PmtlayQx1ZTOF60cvTa2gLm2cCA+Dcu4+KgKYW3G0N0tDWgRpLMFt6OVuPrfXTNqnlc
q+7X6kZxDyXt6pxQuRPCuyfBm48cPF7vDhPHXif6tUT1SsFhZJjc4+dF124yH97cpQCuqdeDVDlt
ipZc0mFDbuBAnOAZKzOw5JPrx4UPs3eD+32flpyQ6qaqzsi7I1Jy7wNp0Ode9LcCNMnbDFH7HJtS
D6MrdoprBt2guLXYGP4G2Wl2kSQetG/eXAn3MmsgxQ3wusSKSZfFG75EledkqTZc9M+qviCP1ItR
nyddq+Gq5jxbimr/m87TBmtKmkYVkopsWuEdS965c9GZZO64rpLyHCSA3KW5QMwx04JZOOKqISQt
S85nTBaiE1EZwykjemU/DY76BG7apUt/oyb4EOs2U5eP8gP7gesFVlnZ8IrLjikGNj6fIwZEEJVb
TPGLTrzYGGLqh0vfod8W6ajmKAkIFyFJoeaLKwjWKT15fDaxu5/F3BzB+hx6aDvoWCiS6wF6AdX5
LCsWKVgEYu4Hk+Z26pawCYs66gl6ugT8oPRUcMkvl+w3cXuYlh6/n6PXasYW5jr1k8/AVfUM7GgV
qDs/gDBy2HcUFLOAIMcY4CXMIb3DBbaQ0V4WpBnHeJhyB3LRFKUat5xpPjMC/5QRQ484+23FgU7H
kIzcNxxjx3lcAm0jIiOZOqnYs/stwSsD1wlM2Bhk10iOd6N9krXZg9hotB2czpYbWzIxDnI+WaAA
iLS/GoBWaQn6HHehgI0LLnV/V0yPNjjzEgSXaTNLIZskc/KvKdhOBmpkfqx1lAJ7Ej43mmjD7K9g
nComDOk6XiaVKhDw2qI1d8CNRIYRRbLqJWC6ZzGxveiC+K9EqvUxQSeYCJEJMNsv2kTUITN5dwhE
uYGW5UujOX5B57eqZ8vU9sXhF3TrJ5lLZi5+7vVnitU4F1MjAVioaxNBDTPUQBKLoN06lFbjEBFG
PognpMZAqSol9Kgqbe+uV8SghCuMAcAjDu65GBnZcUFGMqhNOlnibSzPRKGtgFMO8S3a0/VTPSKO
ptpHuAz0Hb9Tx4wkQRzA71tCFvVfcc90GkqfM4Kgi/tnzclcaPOMlkpj4j6/m2p39/1CWGbjHZyq
xZ471WGiKt/HyoaFrLJkVQNrzUMTHcGMBqJDk6uziC6lfQ9ChOtsQOUM7AhVJo7amivAaVz5YlQk
I77ir0EvrDK4XJgjCmUS3pbkj1RXnHmU64OPZIyi2W2UpVo6V1kRcdFPz1Mul0KJq34+r/FNIIRi
EOGUPAXVKXBxHEG1hjx6OyvzZkMnNBp+xAgTK3bU8JsNW6mjUQVSA6+lAnQkL7VHaIHKQeBm+dbJ
V9DBQ/SiTv+oOotRTLKyWwuT//tjCXaWiwpHf1ccbZ6apnTRV4H+Q0Ldw7HfO09smdx77d6gMRnY
9aCvam1Tl8nE0lsLkzeQ15Fs+jke/UK8eJqRWW/+D8h6Pvn6ih6SW77gLIyWxNd+YtIPnHZ2XVtb
0bZnCKaUSdeh5CcbNYg2bt1VjQ46o+fTZIY+xN+PzFvR8ZQ2w24p2vGv4zEdG/utIMjvxsh1U/sx
avh468kfpcLjdoI+e7etlBEDJZGHrrqeqDMc05WYTFbZIqOjlNcVYYCP8EgWlIGFJT/btOescKWP
MW6jMR1fhPu9ZC82Th3ulvcfmIf+pFM0Pca90GXoLNcaYibj3aDs3lAzNsFgHQWiss2Swm9hE7VK
L/e8T+6OIjNLQlzrdEGVx6EoyOQLJwDiuTuCKr+FbXbsPPbRYHN7G0fOujLTD0etmHzIo2TAI1gL
LDnGgSyUdvncfU1DyIHghGSU9EjAw3/d0/dg9zS6DAaKH9iSOGQAj9yKbQXyXXeHVmggOj5zK6Xb
WBfmKmVa0YAX0gCFu1UBddybY7bfslrKL6+AGyK0t8ik1jcz6A3jdiT9pcWk9Qg2U+KrbnK1a6xN
pewFoRgTd61it3JYs/52HX8ZjIJKN6ikkXsgLe/+PJKN3nJ2nuvwITA2Uq1Yo19caJJv2s0YYeVd
rJhmsnO1M1is1q7f6VVIVl+sdA9Qpx9pFoSlgqJcxa3+8lJihq2pOnNueXig5FSPIQS3nY3EcKJj
BK9gXx+ESeBRxfO16TsF66cyEGO4jwjnZi9/m7EO2wlLmAge1x7oaCKDsY7eO5XYCxDVuTBm2FwR
9MrCqdgUdoGVg08/SvFpdK5fm/jyRzf2b/I0ROh8nIb1K1qxxfMlBw1k3pkI2Z6/SNnKOBpf2len
8o+Q3xNH5MzZ8Vsj2dU+e23teqi1Y14riffyDJqkNTDpH+MCQeKBCvUMI6lAIybL8HYG7Lrs/QDu
BV/Addt8a/ZLEXDi8VTK4/01P8nGDyWl6wfXwLhBS935W2A/ELH8F/WAxxre65sJCRaqn3w8Kry6
ezarMnw4EuUGPkPzXEDQbWfMjUkzqnopPxlCOlStaurY11ZaMAqg37iAMxR5YDEZxriDRZebQL7p
2OGIHYPSU2M14uNhdrryNMPjG7RT4Eux2EgcCdjM7DDwg5qIFFyKlrIbqGWcbbTBUbs/oZCQJpio
VvqEE6uw1oAOD2m3KuWRlex8IjfoGmim/XkPHjR0A+l5Wa19IfoKySpS0rKlUw/PAXqLXKPZa6IQ
iRApIf/d3+a/RqhV7/i8vCYiPZbYjBPQHYRi7j3pYHEi+FrOLg0E4NhWQSC8/z5lvFYT2auwFhsT
3BM7E4Kg1CaAokxk2sO4scF/JZ1gq2AOcvYixoqXfnKV/OOE2dKPNVi8wfkHFLBTA2J0vreocn9o
WJdE4+ch6sOj1Y6yhzkVaysbb7xA5m8+drAMxUoUHNKm9dqp8hcfG/zraDP/UbEtnPwS/QRUH62+
WW/nhFqe6XAGTjJc5AwXMd7k8rmDSU/v4/hKdjPcdopJTExXsSEmfde9qM7wwouW6ZJzTFhmiEjQ
1e9XmDJDQiEZ3o3rIBV6rdedy6gCjnH+I60f+IxU4aYQ7k4o0vuyevKRv63j5IHeAjRbf8EO6RHR
UxeetgPrLpCbrPTVxrY2MjT4dC9bzzyOOCK4C3ZFML8Jhe2o4UlPptJZdDrbFBlzm4+qmbPl6okG
EGkF6j6j454K6pTq7dU8zNyBL4iW+wN2And15Q6G8/rkleGVv1kpqvk4gvflmGBvoDLdX6XnG+X1
SQ2FSNMYR0vIe5n3PYN8QaELqYp8vKnuXCo5QTH8WJ8gDu2TwAxtZm+U7oNe6oyBvFnEmQj9lEC6
6+94tQEJ0UuEJ8TDtUWWeR1JgmrMWDyL+QaO+vfcGvA8RlldqhBWdVMgekc9xq2s/ix9NjMWe7mI
kQoOBHwSdbpnXfc8ARqVy+a69XjGL6r0A+Xh9uB95XwViyFuJEKx/MWmmR809zgbgAWmPIbfM6lp
kR09vs+S8ei7Dz1djjQNcWoowoef1279jxy4qGYrvSD87ddhoyUQtYpM6XL0tVyuq/YR6WkMEmfI
TKTb91ajypwCN6hUbOcxK+jhAiJTWv2U7Cd4JlQFN1N5n0wSj21ea8vjrWaty19aISWZhBw3Zy91
78nj3XCJkO7LnwA/eYAiv+NWc3ee1wtXQBl1yNVzSYRAXXNyB1kxRu0yl/dgRt8pBAddf+rQlEY8
Ajf24qAEWYcBNoVgYhYmfcGOuvNzDpItiIVNwFAqCXktSGdX/bRLC1/b1kMAogFvSdnaOIIo6jre
5R/MmX3I2oyIf9cwK3frkfZUSyVp9iL0bA8J2wQfvFPvUIFNUVjRz+5D35aa5ZnuB0Ub6tzxhOlg
B+ERU5ofD5AacwyFwjHEuYt2xJDh97aog/VtHOOFR7Rq1KynwIgFo8G8j2NkC5TS9nrTO6FXGH00
pFhmlVNyOe5eLwS9DbF5guwfo3dv6ueEFv2DZdzldVygymlm5uJc4l1Rvs5RYJdkvHbRSC+Avn8S
ohcBu7SBAbuw2wOsDxq3eLquH09AW3NhIqGb2/1ks2jblI4+kqow2wYdZZgqwbzBF3p89FgNp7z1
CsDf1nAvs7zx3HfqLiuJQrTiWSXUPrb7FX6Mx8UVJUM+wk1nD5/wR/kSVTLQYuKP4xtUlaT/51v5
3aCc1YAXnJLwjfXCWI1OVfFrmpcPfIarOfz029OFDz+5VrdJMZv0d5hdL8RqFIqeO1ycerZyTWwd
wmJ+FCUhFCdl87n7SpEWz3r7ml/WD8KYh0zTDkaSeX1hNT9leCDRaBPY3y8HIl8mnpWu5YjQ5cv2
czPbRC9DsUi0noPPjx/I99nf5yQvE8NiELWpUYhe8/kmGTSY12BCLZIdK/CVeE5vKZRIAnHkyobb
xJF+8nY7RR56iyVHES5PwdkreZWlt1lqK4tHBEQonXRCSafiNchiE4Jv9b2EBeGgzHKDcJW5yQkx
7ln3VYYhSl2g8HHeTClzuwksk6AU/HkhoitUWbEBL62XBZQ2DecYAsG7RRMDgTkRUWS4aBd+HbCc
B2irUrcBSMafLtmVYtBm1tKt4qavgUECcpSYHOxSuCZbRRWQThYY6w6fQPw1W9+XPghTSa2rhLfq
fso6TJU8FogGHp0dUBoTGmVRiDgWO04KC9qhRDDSVj03yAgTrWoZaUUvSknUYYfY1wEAFg4aQSRr
usPBv0NqD/TkOoYvOXISroOf8ts66EKC4ABPP6rTRt13HTC/aIiOSMrEv6SgT98SJRusVGqJPxHo
dnQmkAKJmnxSXH+Yav/l31qVJHiDm4H6whNsmCftMWU/4Q+jV4N2I6m3oHRDFBxc0km6DsJAxkeo
DisV1h8xOgrfDXOAvXNuRxM+KC5t2v9mYSobi9Xy9RWPIo2SljYB6IGN/TU1Xmr6E9wSk37CF8JG
iG44J0oPUF2JyruDxWy9V7GoHlxG5/DuCluxdT3yo425ITkQDs23RmHlTRS+f5257VwzU6CGLK2o
JZSGOp6nplGWucDdZJg4E8lYvJSEUK89ah6AsMIZYxOadQtiIqZ74D5oDKSadSJZpZBayEzC1mwt
T4J2FEsN3ohMNIUIpU5gmwdvvnrBoOstw47g/OjscjOXKOi3/dxwPGkJDbhL4ae5MxSUhwseizjN
f37Xy5u2pHaWSYOR1OSm6vbHIbq8D87PfGbZHcSSYjXPm7XlVjU8vgTSxqlL1DuRrE2WyuR+wrJx
hhzR1OPqscrEztRfuz29F9gagr3sSk+p6iMmiHtl/4oRjhqdnBmIpzxix/tNxdyF11neO4alWItD
+A//yYG8QuGJ0Je2M89PVkYJrW+V4n8t6oYALdONH1Sb2zCzoe+NTZ0sIAGH0wUTB68ryU6Axq9M
8KEZCQCcuQkZ5xDfNxiwSZm7t6ZPipcobEFlQWC2wkuPjYs8Xo70bflQAPi6EW0AVw/+BP/khCv3
77zYoAr4ISEKV4HkQGufqlvzS4e8EiYR+BEVHf1tb0lEc/j+eAtvRrbv/s+szYyaP8PvKt8qdgL/
NpNjYiD1Dn2mrwyqdU9Uq8xnZ4apYEdbd3GGrxsAGcqENWSmxOXJsqjv/XMnIhZLlaMZJB5Wcxbl
mRK3qlqFxDmzJQ2RZRFjR5SShPDO0/G/i4kV4NzGVVIIB+Hu2YUjP3vsyrW/BgMf0/S9eDbda56K
5OJ46+cxQSoeuocUUvxnZ54tpWt5Zi8yq56sZ5dNZu4ZHEIprQ/ddyZjQou6Y3MmzhdJuCclzTrH
TMaQZAhpamaPw0uqsUam+zwqzTrdOCwozwkpxxD/FgDloyu8a4RxHUpMEI6CPMy5ovRTg9ASKkrx
K7Iq1/URaaRdzoidFH/eBdgPstDp1GCmUa/wXTyMCg3NMihcvA6zbft82NpBh4Qb96jtZVEnU9b5
9imGQngjVbOMl/yWpp7r8705jW/Ypgzm8EnrMfsBhRtp6XF9XYxYSYMKhieTc3XJodYqs2tytQDl
N3+C6BYs3OO5P3D/Hp1mW6hMraQtBOwza2ThOCG2fwqT27Y1vxXBsT9hpylTQbrQL4fN+e9cCMNw
DJaADybjS1LmKdp3Tl5nKxTJ46OJSdULsaER+0q/kgolE3miYy4Ao++s0MO1YdGTgsBd8XUzne1Q
1z1/loQv4U+vj9jBGf1UMdlURd3yNuyl9g35j44ch/ggEXEejru5RTxMh+JKiO7rfoJ7UQMoMmN4
l0SZ10zNcXei00y7s5fKuDK7JSc1S7UeKU5DauRrvJy9RoZt60cLMaj0Lw/zYQ8cWy7c6qHYlUIn
hfkZ55hyd4lwVe1YlUQL7DZlYmWpfw2cf6yhqG75pDw95CVFv6YtSN4anpvedmbPwR151+Y2HEF8
3QuG0zqrrhZPReZW+v+guVzsKF94PiFLOzXyVfbs1rDNBYkY4oVr3KXueUOC3N9Wv8pVDLrxJuZ3
r2nWo67CxPJ+CiR+vPCut1H0nRsW6QP5fDXGMKBsoNL9XW5dP3Wip/0zA1q2/rYn6CBQjgiOUyah
N0R27fmhjNYKGmlCDVDAuzfkNAtr5YYLho7niDHnn/+St1FbbfUhl2/C3tuVs34xWVpeP00FOvKb
tV4Cojn+V2oGy9BDwMfWRrXktTd2fYlWybRORbFgwsJQSo7Law2qvEyrsyJ8xHBXHQ34Z84vyZRP
PuCUkLqD5fE80dh7UxAde76/RK4VikhmqThTzTr/gfb3YuJECoxJLCbmXv3noVXMbEC3/qYu/y70
WLIrYC3EKozIAjnaTA/iDaWA8FZ4IeSZVRAGZgbCr1Da7s3Ru4uSQBJjnElR3JbdvPvGWyGS13V6
IeanBjZies9TKbf2FP9x1lssn89vrEHQIz5w4qiusbYtzHqNWoOBw41VNccU3pUF8L+Bq4tZPvmb
tblgLXOuCeSa8Qvwyo/cPMm9dss2wiVIurqkUp/7RCxuB5iaQDyq+104LxHPX9Z09mBMuI9wpSVu
XIV4EsK1BNwKtNGEVxL37jAJAhHg7sN7VWesJgDoPDGuHfZDeogSzun0D+/d/AcaC3h94IaSAc7H
crr0VvTEHzGN8Norowb11emf5aMYL3QwT1HDxSZET4mNSCh/2K9+CXtHH64T9HuSjtfhCF7Oc3OW
EOM+VZwtux9F5NMKniKltlieQdElQiHnQXjRi7FHSN8A5nR++yiZC++REpJ5zdqWPMsLyGXtRxO9
pxQss142yK9mHoLOZprhHtqtPYU5QTTx+wJqVOZmKXHgMg3EcexYIcboVyLuDVflgqXvC0Wc1Rm/
hElYs9C8iahaS4nZDrrzKCpiBvPYybxgS0xdEbtD+MV4bWzWzCZKglm4tvgRfhP/UCEzRCyJuVL6
xMggQSLr3KOTVrGYL4fyQIi497nMCXzI21Bd8s5BTVsPTA0C9zO+oBWWE2NAK1lBdje8pkqQunl5
PMiAxC9lueMoUSWAoQBnBjcNNUQ6GXoT3PvFVidR5ZF+zd3IWUYBCeX8O5hlFbwxDTYgUoBt9KfS
DLVMBPjJqNXdPp452qLfbhAO8nLq0h4b3a2kiwOG7ymXQOrP/CNHmXYNHPyw8NNhpoLxNbSZ/szI
MBGWDx1eIg2nwNMh3wnXbRkWzRkDQwt2ocSLqZpO31yR77bcrKIkYij1tChnT7HpjXUqp5ZeGp15
1aSxdMUzxVEA12lT4UuvqSB2C2X3AZF62WJGCAYQmG32TugCcVl0ZFL0w2Hkz3liuWmthT/sME9I
uAzpt4fLA4vzqeZ82giWQ68cG+0yCHGIEcw627Dh59SXr8KSJ6/59JvV9w8JhA20oroqyhpg/Mpa
Y9rYXAqnznna0R1XwJ2iImAtUqSLqXoB/gDoOKI8Zd2vATI3fjbZq8BnMnOpIBH+0YEz49d7Sl/L
EyJGVb0/70yJkurBPYNudCPvWxtvX91TEy/qUEsK6Zt2QyN6Ug7maYuH95ZmQ02BaDNlP68moGGC
rHVyi3LGbUPd1K4WT0R/7CFCA+HncAhN7V6e7J7SS83fFxTCuOeY8Dl8T0j5y6rOTyzYRF2QWyCM
kQWeu8HKzJiujAUln0e/Z4xLhhxaXOR1T6DXU5CsJl+R5hojJzuXLetzc6uka0eA7kHNlRGBOgrj
Gh/RY0k8WILa/XU70d4vylhF+uVe9G25kkRmcADt1o33NogKfIWo9FhFmR+YThpMUjM6ahdVdyPE
JFrCK08knEjFtU1qZ7sXP1PDUNkgow+cpIPv6hKkVVo8klT00CbBoJzS9v0+dIsxjRojOU23xuAB
9JtN8RkH/dVC2iw/HIMqJk+PcYWubmrntCtnTrr5o6wiJzf2xv96m+8dO1ewx61CCzdehJ9VRrvt
lDdYXYgUQcdsjqrzOy1lgTWvo2AEpYTgDl4Zq+H9J+vbS7jzAeENTuRb6TXyjTsJ4VbCM+xfiDQu
gWOVyQYPw95XH+PUVv7O1IegaA2tV3ceLhiMS+CKCGfuooTeOXMFznp+hC/6rzvqMknHejoOzlNA
lFfgEjdmFaYmfIqTbPSPxCgmtfznX3yXRujRwd8RuMCz/gtDNtAP5QP5UjGWY4ziFossNE6r94Ne
9AWwVLIqReEUSDX7wO+WuUcStvVO2bkdJQyoZJECHoH4OoarmZVblbIAeCtDrkvrWmPr6+crEkLX
WfVG+mMyo2P6sebL0w3ttQXCHEgRZ6xVob9OXkKf4LmeZ9SjPafi1UH1BNrIbQcirgi4o4tBWAvz
L8F6KDcNqVJtPKNvCDzUHopwboxMnQaHtXOC8s49xag7bWYYNl/FQserIiilXNf4QcYj56jiDCgd
HQJ13WR+D0I4FXlAZ0HbiG5wK4LsoGS+y5qTdn0YtGYbihkyY0wIWeAwaYQw+puibbplRVIBvniq
NjHP9T1cVciByBlZx1jsH0b10IMNG1+ndiioRxRExe3TpPhCycYEO2swc7IsvtFLHLafV/eqqlIe
/urljgGBXC8o7WLCLb750NMNXqNkAcNCzLoxxIQDMj1GQK0VdWNeMEl38TSbn8TjkSiCGdzpOZRg
tFJDjGORgyeMePtcIziz7rwIR56iFA8U75lOlxGvQR7i8M8djVQ1Iz3oJEnHUqPE/YRVQIpk0Pj7
UQQ8yfSeqUhTmdh8xvXLaMD9+bDTR5RiQ6+6FCKnvGtm8oIZDTIxCop0QlcQcpv/YJwjfOVw7keL
7gpTXtDlRooO+AVyO2TNqeT+ngTarRM0ro42/o1fVIEcNstJ/pw+3S3uJBkv98CDD/VN9hyt2kJX
CeHcZJWYzS9gZOaEUVifz5VExklYGebbLuQcTcvY17r8OeUyY2IdDL23tqAIQMGZGtDGKW6Zj22a
XA4xRPRtv+ngrDb8vxcLU5iT47UYoR7RKaL19uKDk2MeVTpNn1d0XlcsDemNJGUyCms3vu4EKixc
NmHaLozddHviAvSGzvNqJ53k8ljvlf6zROCOGFHI3DR+YzYoM+C/T0W95doyDNpUrwNa8907OL2d
8tKRrXQtejUWpe26QmwfVQrLNhnttT2bi1DEq/DGuBRtYdCDf3E/9sJYDc5PfEYsyCdIOAmt4clk
fIohS66xtXGxByBDTwec62JjclGEz6xGulTkXPWwF+d1RnTPiycf5es50YMWWQMfvMfwCKaPpOxC
U3ObUGBMKHaIDGfjNZEViHXMcZyFUy83WOwfdcX/86NM7Pv9jMAc6LOSrYZheK1W3UcIHVdEc2vq
qmRYke0Y0C1cdfbvZHZ31A7YCiE6zg6hm2m4X+7Lsni8AhODaExq686v1Bdst8lf7YFLIp0d+psM
KABAuG4jjnPoiLAW2dMBDxs1T76S5t6yar6Ecnv4mk6jEvin1chFjQ3gNYaoPSzVItxT2PyV1apx
b2D11Asos+z2QX0wlferKRuXm36z6FzOUYCVJaIVqm03gF0WSrVF2Qk5qcNeGreM2oIMxFH8aDb1
uXuFQVpsFbGnraHtw5M0Qvq+DdQNQD8r/elKiUxQL4KkteuDIGRmrxTruhjIQf8q4ozisHT/eT2D
oFCNEJgaaJY8w3gWs4t+o/LR/1npQXHlET8h70rWJG2CYGAd+ukxr9ezc5HnFJyuPZaFnUSygdmz
e2EG4/76jhRF5lu4LBJAZa/MVArF8Tc64PCXLYoB52h7pMw5bot+kLjYux/kVrWFTAQG9jPR+roK
5XBAaFw1gWOIRkAdToNS0A6p0O+wwYAchJxa4e1qmeBG12Ax4ht4CWAlvSNuUyUk4e9FKrEVHpF3
ZMSmcf6TbwG+R4UUtB9xIGDEIjtiUdLxZ3yrinZX7DbKkcpvosaqH0PsBZxHfJSUAYXawFkCwwLj
dcYllqfszvO1+B7W+33O0ZSdlnPis2SaR4sCNwwo9FAfYqSX67J3gg2F8ihjIriUc0o2jkq0ZUOT
R9aOr8hGhThatzCXSVw6REHOfQ2Aw7ABJo5BMsJoiCiEa0RtaSEq3Gat+2qcMKCdh/VBrcFhOrJz
t8SfCH4CdV1peykD6RvFtLib8co4SccH6K+9jNYHe2+Zk0kIBoWFSNlZ3sIdEPmD0pndXZGaPtij
t+gRPj1jfL0yF0ai7z5qtAbixA3XCpWL27QswURVZ8gEMkSS2+HFXaH5YUqF6w+OREl8BihU7uh6
ocUdnSX0TP48eXZv7CCSl9BzLH3ESRNn4R/AM5VfCZtOkVmQHIo/uQTYUC5E6yf6ArulEYNBAvAA
BEI1QErHZtUuaHV7wkE5S0WpBp/J6LzS2xtVJ/ZTg8pPbE+t8caAs/pKJspXNLqXqa4LSWntRDiA
XAUIrIXQEjqolRBV6CAiqS1tzQLaWBbLLOZNrMT2fSINWV526f4vNqGhfZDAVzICL4X17Lu5V5/J
zIfNHDnxBfFBT05mqN47/cmKYlRGE5PNMu3Zr8ar3Hceugg9CNcX9LgWTxnmBzFqCt5zaN/OFkP3
tffNRCg9LAaTNcph1fHLfw9CfCygTWEc/7RUXdkyxcP7R6kQOY9kkpKSEbMeEj5gR1i5wx4m2YOL
teFEYYhaIZ2NsWiA1xZ3UEoPxP13970EzoXdBJlzuCQYn/y/3OT4IJ3uQ5u5fmOUmRZ72CbU5OVO
Q0ypsX7DJqWf/d82px2mgl0Sj4nvl1rUaKvGQx1FIa7EJLJJKn6CC+rNjm6b3zHwC4askVdRvOIZ
yIG4ygekWNyLjCUoOA+/KaZf5C4ZP9qpkKgAV2hqVAooou67hR6QiBuBJO5ETAi7+kTad98UVM8d
yWRvRSpbasb4vC6Rnnfp5KMLy3co0IcpKICVIK+CIfRFwc5Aaf/83PJHHPwDVgjycNL46jRR0lHC
J51eRuyIyrlYlkTmsUtgdbRLJh1xZ6RJ25Dbrv9+VvVqZHtQa4VSJ01MIJ8w2XV51JLurtPevWFO
We7WI+VciQVopk2T4jt+GgMLpLMTLmkJ3IdImy38ha7fs+jXBnEF3iLHgvYJjTh1ciZeK+bjKONI
C60Q+fMj+k3h5TAQvxf6IFpU9K6T4PTemmY4YSwOtBCXo9AkFPCOkdPciv8MSkqp65FtN1OO9Oft
it9256rLhEMk9/3TjAT5w72oj7NI0tW8UT2S0rbmrOy1bQ6Q+woSqm2stzZHrIBDdNGYsqu7nBg8
VNFCpwo83UYcXws18WLdVJqb253RiHBEdbYwKj5aD/XK0ykRvrGIgvQn3ArY6CewaqMxFxItwpj+
9TszkgxwmRsb8gkfzZMRIMj0HKwaUsDUHK3PoCK6nAWfo+GucfGF1u0UVdVwgEtX23iqAg8k4wEE
rydEiqz2y8PIvk/kp5qbD+ZzcK//L4lyX48j2S5v+ZGFDO348Udtl8SRgloK2rGy8l9Z3e2tg1TY
J8vb26cIfxwPIUotU63zeEmJpiROoNphcCRrCRHzQiUTMMfxS5Xi0hJjnePsgTvEQcx5v+Ff0fd3
cokLP7/8iNCVuGyuzZPuXHOzG+xsItC1yRu4AMUsWRxCOIrsG0eSLB3jbkuWXoEORLZegnQgKtje
2uOfbD65WPxPtAZOndvMMzyPBy8JH5pptqvYMt4QHqc00vRE1dEYY6kMQmTSjyOi3FNddFEouFa5
A34INkh4cbSAqGg3JixHey1HgJwF+a2YMabqM7/GAebsR+Nh8/6M/7caIFBK1bHzOC13/VjJVlJq
vm1fzwiUYnr8Qo7q7gvgmsgvlOO6xBkTINHn6bomdNs3lOUjcG2Rz0hicjMLOqtVyUtuJ4pyR8uH
ZUnFw3t207CSFNEpu2TnMkC5pRPHnnYuyrlrU/PClb8sfJS+bpXRraGTQYdu0zUYwYYyVwXUjt3t
XDF160zkCxES7csCfZ6CcQt6qFNBVXikQGVqawVn78BsC/EU5v9kKbJzoqnATv/ZWGF2S5Oj7y66
s/UWJ0wXPcg9zVavua+bas1qP0FLuCS/8RpEC4gwS4cFRFb/W6atrC/bZADlgrBCcR4g8YMxAFiW
5pBokoMzNjxr5a3+PB4kJnIFmg4tPi7wCBP+K+5ibH0h4YgxlXo81OzMP1Ltqp/Mwihq7uAEjSgm
8s+feM7Gopx8AEHZTtYNZZai2WRBMnIq0gB1s7L4BlZRnYXFR6OdcOiBVg+ojFyd2m04io94htQK
FWu14RvpWy6r8NI9f7g0JAtn7b7dM7pVDTqSMgmxzPx3e4rVZujZdd6Mua5RPqEjF9kd/JyJwe/M
Kwb1w8bOzpmu/MOx3WBY8cmBfvBOTgs/Moz+Eh1+CY88k/aQWlaNp5JPEfgmAAihIrLowC1Tlcd2
BwwUxFwdmDRTnFNpWyPw7I4YLfjegU4KJ1vuX1rjENrj1jRyDbEKIANzvmhWudSWDCNAUSJdiiKa
I2v8c70Td0UtP3hTgVWisR0/oNTienFK9wDQTUUpHayoc+19Dy2kACvtYxKQxr0o5JQ55tRkXpIS
zZkuTvw2vVjwdthMBX98fV0MUKF6xWDHvQOjPGdy8TEkak7XgEH5ID+rgh2K3At8KeaoEKP7AmMu
h3ir9p5eC99bW0e1wmSmRZ9d7smiMGdS4hz+7gyucAjkjuBrAeFfcvVHsGGeoH4Uw6eGdCR9R9BJ
HqmK+viWlWP3UNttpz8Mqu5clVmiqY0f7xFZ6FYZP5+wrHl/EBt/9smJ+5+bKwA8JST2Sg90dSq2
Xg8J9spbFW/hNrqtIm7H4yUXv1GQwWTjbdD33OSJFStVsAVxTA4dDiNyMuRUPqsNe+imivO46AX1
i4wxNKtmhqD7dtxDyCCx5RG+oKtpURddNqksXLqskQJM7rwV5KzsBdStVlPqgCfm5U3xC9Npi9bH
zICocp99gOsRGjDy7H8QsO6rSeNIdqIREhPZIwwNDrF5u+tSKXENnZRRpYJOSShXtVUJVetYp4B3
lLaAP4ztlp768Oy1tE/pReGECZHjm8hiCi0INp4qpXNeeVaHhIM9YEr8WQwnk+kq4fX7yCjIq4zi
di9z0mLaUfvjpXuCmWueQ0JvjvpMtk/SURAeELcOua/pNard6AfBNso4/RB4OQrp7tqbR7u3iScl
nczTNhkN8ichlogj4Y8aTXyXa7YaJqLR11b4AKV19Gh5+7NjedTQ1IiO3ETQtuHcrXuzKRP2UmCH
mdjhqka4dugG98YwAo89dcbnoalWTent9q2vDQyQhdOmNMw+S/vBtwXLYWie5BClz7QqGgYyM6He
HdLm5Mi2NelWmgtYbCMMxDRol2x4D/iKAnB6KF+FwDq8rul5ygIpVSPFa5bNYhSUO8RiG8TDn5Qw
g+UE5sg6LMDX2Z5bZfq9bWpd/iE0pmM8/0KL0rlyIiNu8zswXS9bBSy02piPg9ZyvKbqoujgvveL
t/WporZoruo+ANCIJxqIrXlMqXAD7JKUcI5pNaGAkTs0P7D2aAWFRGvaOV1zCjCiQn5rQ3VbWpcR
o8CeacO5WWmSN45GDSHoHyWH/Bx4HtKEHbKfpoCYKtF5VNV3udFhguxjOlpLgWV0wFH0XdnoXEZh
c4giWUi+ujGo6ytRMqHHUJ4nMo1Ia2Yctre8BZdNj+k177evRUEAMpQ+q2quLFxSThOgjNvY3WSD
BVO5TtQnQmjPobQw0ucJLiteTbwao7sX3b6ZTLXVfzMw4FrPWkyVGTFFbRAH6WGFTvKcfASlJKIE
aafvNKhJJ43EKn4mw16BRS4J6CvBHmEdEDVEQDicHAQp0ys91okA/C3OMmdONMBbEnS4eqp5005K
NHo7WPkaybPPxquASKuo8KL3ZyabMS0no5iCnN1K5LlQ3ET9ZlRaz38IuJwQZVVfvv6nOcr3LNRk
uxtpOxJv6ZsN4suaIOdcSkkEl36p+P+soBBqYnBDMw7AP7e4w8mOQM8UJAWJvuko0RVu36fWTQih
iI5zRSSorEzDm5LKX1E3i1HuCVp1wTVtOT0xMu9Qgn706iBBId7g52A3eR4ah1o09r8KmuOFgQhc
Ezt494GuV2NqnnMNyOWr4qvWTItPB2vSrbQj+FsJ10UBSgg9TVpkHQ4Oj+aHwkFONTtH+HNouK8P
4kCSaLuH719BAxQap3HBvIBxE1CELO2x8S1sB1Ku0EqHMNUz8JdCTg5wn/Rv4GJljd6JO7yFhvMt
j2ZqZdcrxyMM66cGpH04DuvtpS6dmHywtgeX8lQD0PJ53JfHfLdnKRJfbT/lEbD4UwGx0t1PoNFW
lk5d0a/eEJ6RDHqnkSnWia2lb0LVYhe0ttJ98RFsezFyCfQS6fNsxe/5Xd5fxcN83pMcfLB7ILmp
6x8+i+Vfs36Ja0MausOldv1OWUPhkeFIaRaimuvn+hiyi/UWYHoiZkkqBq13t1KJPCMTjnWCrSLW
ozl9PeJQ/7VuiXPxh5sgSYqbGjsWA/mWCaXwCRus3gwCqLRYY6k40Ev3AR6ulArVocrL4in3MCjj
jFCMznk0CAqWcwTgWre9Ftuss2f5afv0WM2ahI0ajrVSCO1EGEpJbBvmdaKvpc/z2MoYrZybTw6O
8DLKI0D/J8mUQlZD5M5lmHZrODqM/adhOiVDTGo/JIHupj+ZXdMKAt5RNAuqiKqQ2MANRvKzl6GH
SqGPNhBm3+zP4KNtZ5vuu/aWgvUaRMBRfW9a/UROe0aGXLCJ9MPdFGJV8cAVJssH7HJvURsM1ihX
za76NFJJku4bpib3SzLq2QA5ZRL/c6I1yJ0AJLhD+88jCzezXxYbQGQPkz34GIzsNl89Xjezl7Bu
qyzxuG4I/sy0CcXWPVA/E4DWKt/xUC6jbwdvNZP0ArD2JufGG35GabqofPkbh91HEefLYP93Txm5
Xl1Bbn+BcRr+PjAQpxltmzyG/I2fN2S/XvMX6EKI5siSSb3f61EtijpZYcoKBmPVi4rQXt5n7ByW
cNkkOVENAsyhyj2/QN9gWntnLN9VMqAGYcjEIqlETZGg1VqR3cECQqpzDeLvTMOVcdHnaQJBjhJR
tmz8tQ2GnT87p+Hlk2tVkRPdyJjKSa+uHteHLaLiVSSwaPLwZipcdX9CvEXtHNzPlEDd5LOkcr5P
x08Lv3wBmqqaYzUWRbXLC+h+tmeGhbnxTpa7bxe9R32fBKrJIYGyBTiXMUyeU0big+238Vrfbxhq
3Lh3tf54T2oErQjZFXkViUGg0D/w8xwMei48B7DuMXC4apmO1Uxxjvk4vvnvjkojkw+a3VQrYQ04
w5mDxHzWdC5sSG9TG4rt+HUDclbGlGzJBPSYD2+WAazBoI0w/Jj5VIbPmLdSQMdI1upgivUe3YJl
DhFzgy+EAz1kCSWVgFw1qmjr/VJ8c5aO/VP0KWqB0KYKks0voBBTZcA8iK7b4CuuE9CCFVWFTwQz
o7rkjEqsRgSNF9mO7o7U9HtJ/lW+GG/mu9TLLgc99GSilrPLBKV7SuZazxWkTQArBCiR7dHzqbyf
gXFGh4R7+Z2+WUK78lHhbzHZdTD21RtBmjET5Dh0R7k2kRusD5ynW52Eqd+iJojKDHZ5qbiVWUms
40e+ag9nvPWhwGefKNSML2iu69f1xZukB4s5X+bkO4fSPD6bC95/22gGgvtGqzrREqmHvwQHYLbf
u0v0hHGOtkaNnX9neCjVuAoZcudiLiqpkLgGzNQ2fIeVxkCs+uyll1GEge+G8HgNqZtSEAeluJs3
Nx2jAo/PiGC8GUQRU+xPeBQwMdQGpuXzAEhpkAT97ERiG7iUOLSV+vbrJSKLTtxFkHhwHw7tzZHK
780NDrX/YNIBMScIFwmYDo7cHea/z8d2mewqDpGzEhF4V8CwRtwAENG5u+/8Wa+amaf8+I9/6hrR
wCopR3nQK2IUYR6HCNW1GTHogZ3EI6xdfwFc26G81A2f7Wp5bt7UA2jMwcUANT8M4KPqsG+ybqN7
c9g1xArhk659tjpvIkWobaL6q18SgU+lyJN8x69FpO8P4ecJHYQdXeRRApVuGMDa3vg6zLlMuNJF
0v6yz/kKmPTTS5K8j3Bta0/11ivSOOk10vH2UBwxu52pJC3fcSjWgRPKYQE6NwKNFiAnI6HeMvq3
1k3LNxWQvaSoTnt3F0HT51PE8dPLPiWF8W+Yctjke4GA+Vjs8w7RECDhvH25vEfv2a/pEyED6Y7S
Oxq6EhE/TodHZpQtXCBXmDXENOfMwXIsRkd5t4G4+Vz5ahpqGLisRRRNqQNTxpsSgHtWau0elmwF
5uLRPgF7l9k7PzuF34yjS5LhT0SDpl6yz5P/G606GMAnzY3xOWhFCx18w7Lp8S/+66iekldQ+InO
13RTjVgrrWv4wdM38PM6xTt5ch0pEun7Tgd/i1nyDMXk0+kLtw/wLbMYWrf4gcTvwIg802CFWVo4
PauKbRDKgz4KDLO+LEoZp48RLgjtdvaFiY+28iVfGVmSocoAHa/4KwPU6edaIrU3AeSioyPilwhz
v/IBVvzow2K5nxxC/jnmTSyT3CN4Xo+4wlDLl3hvUogaLTmXbuPwGoD6ShajFPWe2Z32jCahxvOP
J+iS97RqIaw7gLG8hysTOVgNOyzvOiUWlxUT6upB/LOP/ZNwOxhfOTYcZGpbZ5FWbcoJLRXyABlD
o5/JTklV6YAZHGujzOgIRcOQzSMznzaBgT5sr9NYDsbdbLupCLIMQY51W90zkHZeqb8BDLOtWFIX
qs5ltc0XWhUweicuifeehCQIVZAeFSTY4h0mTHSJC1x6PEsQRR/9Cp5X23IRgEQDTnpfjXJ4qnv7
plYY8+AGOFbSBjWR+SEJuNhPdYyaAlG3FLHwr4KjzSxRKrlm0kDtEBl0uadbmNuEVtIXX4bQssQP
AUqizhmKXq4DAIB1sY+AgSDK0nPomUL5Hy5cHBtl/J3PE1SAdiDKuCmGWZrD748HNUKkHtXaxf0j
N2eXJlXu+6ltViDFEc3CNE+mH+ZCLJckcY5+bZHMlIWjMFB/kVLbdKRkxhQuabaxqMED4ZJmUVhO
Hco3P+obcb5G8c3BcufODV9dVNW6UCl2WF95AWlwNANkvumQN+NyaMmGlkEhYVVavDD2aPS4rESD
f+m3ou7eEfIQG3zzKFajuEWzfXcd++FbE83VsoKk4G01Xbj38eFSnNl5N8T9XPUUedTA2uh2jKFF
cuGRc5donmMr5fDpKwg3xOoTNqNLn4jQgIJy0RiLDybMlDdj3VNCeT5ky4H6R1/L9wsOphuwVpcK
ImjP7x1jav+l07trmccvVOkVEAmf2+mezFM1WfeWeCoyPmfjEEwe+pKfA7SO9OwESR/PFZUlFMn1
78Aou2OFPrXF/1x7sHynJMZLWlrBLIHf6CiOkOTWd48w/CZr8W/rSTYmy1ugLWOmyqFGlA6ElqkN
pX/xI13TnzX18zXmi4JAV6GY7Er7er3ggDyANzRjxA6nr0vbP8Q80gf2C4+amEnfEa5yDyxwWP/5
tYKrMNR8MokKvnAnbcg7TNmtQe0WzOSAo9VLWJZmlkANjgXi/rywqREFff0BNkVT8VMsN6HRJBbl
5Zn8HWzeDSJ6uYnnx5G62oogcldrDAiIyesdYT5VccJsEiHlbjp5urkgNjEbXzg9/fqEw0PN9bnY
CFuWl6nrUGZ5bYaxBLDP0vhiKH/f7T9xUAjWNiQdEuPmymRgasrFjt7Xal8Qs0pubZwQkYeqKqEx
dPL+dTy+NwWNpGeqGKg9ls9eHzSEB34qf/70NMenRmuKcHYWhDjzT8dnwCBZ/szlwXss+soRpbNx
DBbmXisVN1RrhlXVXDyYFN02xsgKa+abYkhaG6pZ0eVLwh1/G0Zh68BtDQZPd5Owu7BZTBdKlYoS
sR1ZPUiBDA/44dbxHVrkGmBiIdXWqm15r8PN3PBwZ6yvbKLpwrxn6V/6OI7coe+MpsgUA/qP8Az+
9MahAhieEuXzNeL3wXJGdzFCezAWkchMc4rRjluecJ9Wm10+/lxM0xwL4ATVodD09wGK7YyT7Q64
f9fLandFUQeSbuloLo6KNd29a2CjgirrsXZvH33ZC67W0krQcjX1YDSZzQtLJZsc4DNFztHvvaJ3
aXa3Q8ci5PAE54ASyKrUlnF2brlYweeQspDu8lTbz8QSW01Hk8BssRld84PAjY3jxRercfWh73nD
EmU2lVdN5Vchoxu1/cbQqKBSDmf9prSJPfmJxmVc12rRn2+jQwrXpCy8hQpps5CPO00qVg9h7e4Q
5uaeThFB5QIbKl52UdQKBO9Zc9NYUXJvz6Bm8glVtFfxbvQOo3cnr+vVsMMYALrkJOjeNG3CUQNG
SFbbOHj4QXuucKa32D7mHETa3X7wHdMxQPbaLQfeaLqtTVGOe5G4FQg2RoyMm0AtFvjm4NyJq1zE
SRYVg1+CLArGb5KbK+dLo3Axgb9KGOhazpKXuev4FJ67P+TEEijWw6EfoJQtEMBd0hRKERay43MY
SO4g+14Uk40FaLkgCcCFiGi+3reMfQD564YbSgYUNHS7gKDyHEJ5KzfOIiqDTzgGLc2XN+hT8I0s
DeB+xlRLjac3Ovw3zygIPBy48eKUo/29MXiv50VPr5YZ3yvAWysHbBjKl8YTbtbm6Zi7FdxMEAC1
PfVX5dPfFjBiC254/uX7rnpXmbvwVjjMlyGvqC9OpghCKBFDLQOqGhZXTILi+sqOdEb4H4dmElkX
FVKZhP/eQkoyyLJkmpkcgyCVGDUTrpuWRZP16rb791WoZlx0bIMhxHi9dy4eWY2pq6Tbr8I1sCE8
CONNKcvAYCbPjaJZM/Ya0JHDCrNBARvruI/Hcw31L5fjSatXvVBX/G0xoHsz1q3pGWdFFfHxWULq
zwUqCuLLKvKUD+O/g1Ab9/5HY61/9fthNwlfWCbdg4e+Rci1yqmG71Wvomy4jZG59Q22n+lLHxUQ
JLkeRI8jfiNURpmg1axf8uwN0/yn3wfNm9alAZZistpqKDKcmPYNtPLdu3+nX2tbjqBBNKpNJ8e6
I+XRTtMDjo8H5OKOe9c1qPWVXyPq3MRjq59YAyaNdqXCANOzeZC38T9YE4gkSPF8u+EgNnPKBVrk
iDqRvLMiO6j9iwt6xALqfQlrFIKdhbPCZxrgOkXD/btZivGq/XSeVrSZndfjyEUA/6gEfi//9dQW
4uKIBgbM0wNFt+4nD+2RxDGJL67OEfHj2kdWKFGmoxoiG3+5Kq/FrAtAQAlpGh66Vk+CH4LXW/SY
0cZ3WedkCHAdSasAPse+QcX6ZjNKRZrt3Nqr/uv2BKvwFgu0kVBzV5BK9/j57XIadSU26Osz3sX0
7vNeWvfiABOxATgywrX2ZMBsAX8ujo1wrQ8QQC4TgiDWkUMJNLXpgKTXm5ckhx4fioFHNQLbEYBV
zHBTekBc6Ia+lr14aMAqWk3wIkOpzjjKZ7quyAKqb+v5n8zdxtnbF4jMTFxRO4yMBhHgQUCEByqP
koxI8vfGFIb+jX5zDZCOb6nJAmYOsGRiGgQHAgVUlv121vz30e7uK6kPNI3Ohz1Qh1ahVI9il+80
N1D1aglMppwFk4y4nnnyrvCqMH2V9P4xQYOkJEW5P6r6NHvsybFf9tBW1nel1Mqo0xFdi5W4e1Xz
qX2OGUxz724LZQ4f9gVRJnAt/QVJs5dwhz4XMUlUK6woHVmfUZqz/H26cMkdiSUXSE/tu6kDHD0x
33yl1FfgQqhBowgDZaglkn0ltT0Wg3lJ0l+qyh07T6992RHB9jmPPnscsn5998h0bbvuy1mDT8Uu
DiFRCAonoSf6pVIc4dcri8FbYW9zTwwgw+5q5eXi4uOR0A24Hm9ymqYZHQbOP9/sSpdP6TJI4uEt
HCZF7EBeJmZNELycjl0iMQNqvLZj8uOOtvpxcYa8E3svPf7fZ8iYvTR8GxIoO5JpZzRyIj/FpBOB
KMLQbS4o7ecYGsHP0PjMpMdlkhTz8FLxNli/DakOMUVJS0BMxvLWin6oGt0TwZdOt+SBSyl7Hsgf
k3gMzZ0zSXZaFce3h51kRa6CK5IxPz4/vgb079Wk01SJ8eMz16Yle1V1UoxEFvlsLE8PIy8MkBO3
R9KJtEDv2520if0mlqak5iLjtWDt4Og4IO/wBIccv9iykQTXV2XqiAo082OaWeBYChQq5fHrc10+
KXF5NEUPA5O/sAq3QAolI6IQ7IFtIZ/1fkdT/7w6JZpn281C70mnz/BTa1A7yw5M8gYtunT2/HFI
GYN/QBONxGfd5Qf+fTy/bsyyvDCri8H9DJuhYsD0IrUizC7CZ8e+PbBvSbnEdkmG//SewzQ3wp5Z
8p8q2GJvqcgNKIH0RJscfLgYiX/hafzA1Nf6ARAfVJSgdR0e82QHrP57ZemCmUM05to5IFl3XMwE
eDEvohn96FkL4LvwFgUbJRiv5f3G/XWXCM+jP7UW4BrvGQ2FPCzvNW1OhZo60NqbvbI/NWb1A7ng
36eG6fVYGo9AnBzrJT9c6yE5Le+H6Iftwu5Wg+yW+ohoQucGH8Ll5UBer+N6mxo91OwNQ+OTz/Ey
w7vuBrRCq6DtcQc1VRoabtAfhPJq7GyET5xIS3OtUTBtSpGv6KrnI6lYufBDdo+TZnrJuMj1Chyd
kWABqL/F7c+0832wC4Nrix2/hIGM2dQfYe+yi8CluOgdX8faVoz6QlQ6asZnTqiLhG/dcQv6sfoP
DkT+rEPlidkmy7hpqCWeOnnUQhqXcaAmKrkuDpX6+UynGnz+eu50Nymla/G0wfVn0qlWDc9z6dwa
pWop8Yl1qHQDiJ/7fouyEQySmob2TUKtASurQAKKvvvGsF+buBXhVCJP8tyLIlgjb0VcOBvhTfIw
X7ZLGiI/86TnpRD1D/rFZSOVleyqGw0Cf5RM4u+n+O7SQhbzbtZtGmbYzE1S59LcuK8ZCQKYeh0L
LVBe2MO21sgvSH1XEj9/8Di/sZSvOyefPm7mLnAsYnlRwXnprPEngSDdZoUCwZ28UhXvwPdPjWzx
6sM5RBlxP9CMjY3fyE2QGZMbXKEPr3+/IoC8S6LhbSJs8JATWXzYwAaQEpPPO7U/UUkOaCbfALl4
YVuzuhwdsjxEdX1K+Z7y1ES9I1iVq72g5CGs1+1xxwkcmwC7dDonfQFfsL3jkomNKrCnw07DCuP0
SeywGZT0qsYeZYr5RPlKysqGh27FMDl30SbYExf8LrDwtLDv/jjOUVamk1bWgXmcUWbEHOtuSouw
iC2WMw42AbTla4jZclkA4hohtuwMxJyC2jADvHA2ahf1tkTSfeTsA7eQC8UO6+nfnsjxVAyVON9c
cnusd4tu+qCtyNXcEFA/Qm3uaQhK1mpGwd7ik5I47N2UEKLBn6T7KCz7rQPHaT7CIk+yrsA7p3HS
LezGXLhEbK3KsEYy3iTwnNojA5i4azZZG6KLR7fpAZiHpXmCjRQy6cgWkvQWV6NssSm0DTHS+JFk
GUSZiF4Ci7cxRhVenVvj2OENlFjHFa15qRBemEg8tkCQJhAT68wZi60/6+hnINttWJLXRzUetsZQ
R4pp0295EnO3E1TJ8EkO+2nWbQris7ROvYLkfVJD+eJIyDgWsnl4OjWx16Tq0jYWZKMQVy6GeCzz
HyQqSKPQwnRs0Zif7kwKtzObahuJp73wzEkyQF8y8I8ZOi0JOY5qFFrAc0MUrzXz0zeTjHwfJzxu
vw7yRuVa8sCOUtcNh6RJEeE2gYYRuEls7HEHaraM21gulyMnE3dhjs0vL0+RD25IkogdomeRi+tb
lp8uTukpnDMjMXkhmIJ79k7J8Mcx5EME26fcri69jq5ZQoWk0RHLq/y1CM6IuD3CtQnljAzx4Wz5
k3ms0oxl09zbjGaeHmlf3fRyHuw67grsBppsZe3hHr4hv2vWGSxqslu+w1JpSKvK1Mm4RKBWE9Eh
b8Oklf2mFK5sr1TfbwW7wXRAlvEnUcCiTUQcJLoq6OHgs690vx9KX9Nq0VffDaT99AzrSHsx+45G
xaKmdiB7UFI9T9T4HtCoi9gPlgMOvkAKjMcYwVk67dpfRL4REj1C63Q5eYKEhY+PZRIvg2K2JSrc
0a5HW2gL1LNOaLRidjwiReQn+WPO4kfAtikjUcSvUBT7sEIA0yjQ/ijoOEZdKJnP3oli+G+IP32K
MUjHAftgojCayJvfgTnqChfWNQIPwQMpOsy7TVHnPW3X7KuY4BpwTgN2fODfTNjNZg5g7Pyq0g47
RdoE0gY4/vQ0+2t7EYhL4yhdnrFEoKh2py9ANkQPL/+9M2jb0SSwZUe/rfRKQPpQ9QE6QrmnrKK8
Skr+gY7bjfmEXcndkntMTC69MtW6SiWBzqU8w7jkWKty6hMBEcL3opAzn1sd0YZ0fqLla14BTKPI
VDTgp3usTzX1IP66UCfUWH7lUEyN2V0GbCJ0Qfn/o5mfyWd02ARTrfSYN5D3asWLa+zSRVzkArIm
21Pj4eLH0Gf4Nf0lcL7m1xVDZd4FsXFVaNKcoqCB9eXYXO/HoTGNoV7KOr6AeNwT8GBH40zF7Wl4
/qKyXRB6lSEfm6DEWLKnAvB9I+Jurz5wcosvq4vCCHBMQFB5FPe6xoxSA43+98RmlRs2T267eZnr
AmUZumgFMlc7Y3cTeqb8+zvmP6rtTFMkVpLCPK9MefHowLccWVXFTO/75E3Lq3H8VSQeT7NJ+8GE
39lQIa912vp+WhSepDdK6FsVVrBB3Os9JzkonFIKvG9sjPOPn1s65SSqg8mFO62baL4ubVCclYwq
FFZc97NZ6PK4pp8p5W698xyLQ+6iPKnPGbS28ZlwjXxD87Ae6iSMBJa14CkKLhAnoMVG6HZ8Wu9x
FaUbTklujR1mHagdxokafq42U4gJpJDNR4xPX0/VAoiFsUbo2kSLsTwXgpD8+X9rk99NwXsAF73C
1XOebsOiBxg+CbcBf+FSdPhZum3i6VnoyKJjbVh3yrzgXSqDkK5r5lE0PqOGOKMPpOJ9wdyeJP9q
6vmGjWthPMxynwv9Xc9PDzO990mb/b2uge8S3rzc8WdAlm4tJmn5/pMbarR+fm9Iil4OZ9qj4t0u
IQU/FRBBYeJfCWjvtcE6y3siT4JGiuyI81Q+k+LCBvwG780LwYKuJoX8hseRvJL3oIXwt+gPVyDi
zQch33lOJlbuAFNiHDQYeUQ1A/F3pInCgvOdwL03A/CNZ48sWPxYmXghM8jRYpPPV8/lkJ28BIl2
TzuHnv54GwLjB+RVWMX/1LyNqpVkx/HMEhlCEgb7AcTSjO0VjOqO+Km8VON/0IXOfFQLJSOgu5wy
cGHtNWfM/LJs8BVysW4KdweTS68Tei6Sk0LbeEXIrAeU1MF11RNfT6fZwneMJpnAepeatJusjJqK
T2rRVsFTCcUoPNYjB9IWPELG40o4K4EiOszmZNBK2Mrv+mcLwoG+uwKVQfc9wwd6THL+3+V4VQCc
vRnQU/xBb4oKUYK50ShHAobVFyBgEZZAt91NcJ7m6gI0pu8Ex24+kI7Sj6cE+JZy5hw3iZ6ys//O
pAJUpJ+Bn/f1p+H6P5fycKKT2qBC/Cn8UJMB6vIJkBTYfvGtf2RfMm0zN2KVIxxtD490dpKsvdxn
vXfqjHuBqTeHiKpmviEwk1LRYeK9ZpmVz1Nr710irvlwhNLtBHuGPps0+K5z3Rw8HVAN7ZbIiVa5
TS8Nb5W18yzduO8rqaUsroA3Yd52bnBBHa2qkjHJWxW8CPZIOQYJp1s72ClkwbuSRp8NUs7vOJtz
gR63JKxsC889mGxL+CrkLWgnHIxawJPu1ulYexJ35KriWn2l9i7fJkLU6bELjhUgjnDZDBLjJ54g
H/Q1Gkkfd/lP2PS8WVjmpA/FsbjqIMFfZZk7RXvkq+2E6XTWCIr8QtqiwYVTIZ2eSrUHiL5MssgY
QxZmjdzgnagEm5lC/5RZYKH1M+445Xx4ZyagRObNv0w5eItPz+Lhkz0DJvOjgpr4RcqvVnt6F6aG
JlvTzlzmy+rcczrfVHTKWn90+bQdu7cgy3FKzWHsMLMMHiqmgWt0bCMsgnptG3Wq9V5vUW5zLIRq
ugSujoQFHrYkkEar1dNVvrzUlDBcid8zs+EuXIEP71RvkdaZ6Nq1hRYsvNXWkkqztmQAwG5WA4RS
x7A9QLq0jKR8Rw+2PKcVtiSAJz58tYCIa5uB+O+kV12SwHGI/mzH2Q02xKbEVu4tqG+Zq1+SbqXW
PiS3ffsMPkwXKV7Q4AfazgmxjHzM+eumQ9H9+Z2Lh24Y4PVn5+haQmTdhPGpg81mXzSxCR5XaLJw
Ld5QKYO8sBZbeiRyG3y1qoeoLFLN14cQMefUP1yi3VTxa5JhOAviUZxgmjMJtSwOlljf3iy1HH/h
ot6NG+ipj0dLudPRiGfbOzE2mExlHCnVZKv2z+BALJLA7RPVtx/Cu1/n+9dgd0Do3VG6E09bwAu6
lMNip3CPbJlQ7hx4xEAWqeNAZBSNvUxTCUYJ3mawJ709M6HHZ+HQ6TwQEOlVIqdArRHEE6T9kffD
4nBwGPxwj7xXZ9ZEbKbCgtdUHCn4ZI2m8yQjn4zc+M/UNMbtYfht1OX3eeqaBxnqllAzLYYzVi3U
7lYIl/HMidsCfpY1Czm0FUvAHnHYFmgb70OqJt62KAYshL/2guY650B1S/bJyue2dLDQn+X4K+98
G9Xm4bdVYqVq0848xBv+Mgg13+SssB7dIzqr5zggKlFnPEg9drGbcxpfCqIbkvx7ADP6n5ZX/5b4
+BbHetwStiDIlaIZqre5d5YcH0Es3YcdJkAJ6lN4DjpMsYqGbIBX4aaoGrs/2yXkqd8/uQZ+KS3l
aKij/5HSubdLJBxGiKkl9aHeaoO6+TaJWqrIINNxk2M3PPZVj/1qpLe18VKJuyEtAyV67nEVqU5X
tJk9z5Z9ovZa/mCk5ctFEJyYgJ6bg9lprr2fzqoK18Ol0iibITT1p5BKhexa5WKIUlf++QGrdBu+
DKYhUdiBvhXcSR5ifXJYYKHU0bFVkH/KQLxEHr1xcCUIrqoxTpVYNgWY9c1PA9D/6iZR05qXI2op
YHjWVTw2Bjyk/d/jOQHnTOB8SHEgKypv8VxPDejJDj20quggcdNVpHPoVKyCnBRFBG/7q0ep2gHS
HsANt6cBoQKuEKcSGe/0Kmi+tBQBMrcu7a6bt4UsX01jyhKe/w2cVPwMEtwI7S/giue7K5ZuEX5E
3F0m8XgnCdLSB5VAancpOcbLAitrh/XM40v2LLM4XTNgPVrPHoSTxliMXTDH5WdU8fOkdci10igw
/6j64HA+RpqfxA/SOvP0+fXEJzglbWAlG+slY5CNVfKtYEtpwAZ41jOiSfx4IgEX+45ILLLNMHJ8
/qsnAHSCS5eXlSRfokSndS4qGoNvzcymTcTpa/qEHhNMOhojHhGcRg/oXuTRgqCvFN7PDlbljRAg
ghmUdqmHenS2ToP3JgAINds9VsDrNIdLXiUpKc+VWhYIg1RRED4NmIQ+Lekghd102uxyHni2Vqgw
jSDYUxYL6PYrF4ZQ7sHd1UDl4UiZf8wOoARE+AHmB5+CfF0rVZDhID/hbSPthdXBnlAWcyRnkqGL
Sa6yqKLxanlT2CURfv/P3s6g3v4+3RivF1xuWJQ5N+e/VnnvgMzZhnSJx7zw4KwS3uQzm9calEA9
awQUCirpFDc+mZD2w086OfdBdbVnhai1B93w6u4vMrUjqvnNckezt5EG52+agVptdp9oiK9H5gkg
xJ2G8g/PfRtbxzCraSsRj6xohuOBmvfGcdJxJLXUtJSU/nJiuoqanJefbN4k0TNmsLW2Z4+QYVJw
KDaJRbdDk44GJ34zSxCRunKCMz7zW/G23RqDryHEN3ggQKS1iJea9vF/QKQV3QJr60ELex7zkP8P
x27QmeHpv6lzVuN6OfptD1P6uMACrqvIjCgNUNP2cMJR3ukQGGhQ1wj51/0oPgpR0gourN0JqP1c
cx32CEqBKdNKqmyTp1HRVmofad0ebYvIvt91PVOeBA/39ICmIwUHsRLlV+iWzCd8ZKZEokuP+4UL
+fnZ9uH9E0CKdrXgJ0jrfVYyX82uDeH8wEoPbd8IO5gCjJ8N50oWbsxefcf5gdVYZBUFOKVsERpK
8IrdlqFtxmeO6J0oGK+z0j/VpGqzTbsoRbsWHAjW8Z//P1LtoCqqcbxUaUwCT8zhHgGmKTi1LdkX
JR4G7e93Sm1zFkTkKRjSL0HX2PJIwvTM+0U4V2qaK9u2XloC0lTXxqSG66JlaTbnb+2vKYlvUymY
FOc3XjX/vOQCYQmuskhMt77KCwvwIJNgNwUWVjk4BwA6cD1g8sXUyAkCMM9QLIFrKqrJiTWWFKaJ
4KHmLdsV3KovpJ+AD1WjZC1vTEAi2ROjQIUOhiHHK3RTlApJ1I+uoHbYshlXzDRzHcjprfwZkcko
WGxNJ+BT4IIg3+uDDlcybr4z5KYIs69yqU4xgKnDitSasUCMw5jPJ61eQktkPXH4GwLVG+mbPo/e
xiT12AWfAR3KrQDuiT8b0vXSHI9sTn9PsjXJy1Iy9xhG2qFtDKlKUb7VPivsNOZCXkFD1AZYLKXX
ASYSfCNLMFPEClGQDVBL/POWg0doEvjWwGkYyI4kC1R7bgomtW2le8CT5KMjFdrcKmDSuh8AWte2
GUGjB0/9w8hk8XjF3i8mNO+L6oDO1WMTBp/Q9mn9ecyi8M/l3TkAZcr3l4NjVpCdbTFeWqnS5Mud
pLAuCR82/iZJuE5GW4AF7VXZZuOwSrTH9fLfLdElEKiauonrS7DoQ0cs+9qAMS6WR4E79NJKnMG0
ZSlHw0hGv+MudIjjwVP4ofI/xWWDlbANwUIC8YUtPZNzo38IiMUVw/1Nt2O7Sn5OF59MsmZBcxxA
Qn5IRlR2GKwzLhIB8kDSZZS7pRNwMai3S1qtRmDHqOonVTIxWaKSGh7XSzzJrjro28rZjWSV+Dfl
fks44VjYYEEsfYMvbppowBPkVFGy5NQrbLnVK1rnM4cFTjfzpbmDXm9q8Z6EyOjEvXNUds0cYM4E
9IOJlhLL6MnGCCqRa2BCpOBz9VjCygsCoexIIXmV/PkaZLfe8Jycqgv7JqVp+wb/QcyJ9gL2LwM7
6S+NPRsn3rj/HuAi/pRSZ2OBOeO+uy4JSa0yJ6z4JpW9amJDR0ClhUQcACTqixNLXqiD+AfPySIC
w8/nd9+W7kYabnyPINI7lNinpzTxkBH0zPppzBzEqBNqCglpKObO9c3mHiomR3DmezZfECkOypff
4EG0t6aaPDVrJv7RdBhOR8A1ZzPJ4E8D5B1LFfFb8n0QiFFe0ww2Kja4WbSnoSTx/F5iYn24AAHC
MKRcIT+WFsZhekNKpf/+c/7gLYxLuG6zqG5eK4ucSD7Kg3rT/IW9yZKlzaPX6LLx9zPbkNqRLNNq
daxEDc72964uwiPLmmSF9tJv1vm0Zdd7VBL8ErPCCObBLTK41kAHiafGf3LwyYTL5UxWQKle4zex
Nz/LaNq69yTpwY/IWeysQPiTEqdcVbEPOkIQMkw2vaYw5Rxlrbglw6qSpJtBeSv3EYrLGoKB6Zbm
QV1dvL2B/oQA8CoEaSLDPQlTXW4dI8bQGwxz5JyryOem0mlUEx3sPF8WaD97xQqymRyrq6lrahUL
rY4O3pj2u8xOiVXUffaRNt78/cxbuYM9ejsAi9Vkbhes+eDveqk4Fh5T1f+Fy4XAegSXz1PUM2nP
aiIgqQ+P6gfz3DNR9jxmRJBXaQBfICC4XmxAiNaWnVk499Ok71uCcJFunuSq2sZ/D66TfXieG/66
A+ZnuNlgJA/PXqkInU8C54CGBvXFSvtSR62mHlbbWC7g1f8c/6mDNcW1745fbyc82RJrEfz602fA
q0XNGT2Qb6Hge5ewBzvgSOpYuu/zmLHEkdkZnR5aVEtXunZwGqMS12BvxqhP7KthRRS8EJ1F6qf2
QAOHs4ysLU3EozF4q9wvCzPE8qcgJzhco2+JnXvKG6TovPuVJPgZunnNpJgnPQ/mKc4R2fS0pRT2
nCeOgGzmgDxR4YXtqOo8LmIORiqkgCsFlc9gUow5GqEt5os8R21agVHDJiHowLFfm/WZQF7evSsp
W8im9gHTN9+w2qbqi7MxKEniA4x5txF7cLmq4QP2an8gnuqshbJwi4OztTKu1HHJIwsU4B8D/Ji3
sw5LYdOOHsXa1xTlwYdmpLfpvq/nCaLfGzXrlZpVC4XO7nUxdaFV1boxJUK0MNDbvcLGvL10ctSB
/F93a0BrnbzOeQB4PPAa2/o65L5rzBhTrVZavPVrRFFhPuobjO2T+gr/r2WyWfRhaCOvSifzVGI5
CZHHzpVFckaXKwcwrKyTDiJjA+EUIXKf4odXhJQU5okGWXMP5OjlPtkHtPY1FjOGz58/GcCk5D8F
7jR7g4MoGEBV/AiwgoxufQ0F8ab9S1LVMShn+NhV08y7D32sosn2wcBVJ6KWwbLzxlWi0fpxRbU1
3ZiuoaM9Cfjo3AOTcbKiJjZ6DCyhSxe/sIr5lyFCmrVV3Ghy5/smyriAEXieciUwBrJc1YhmL4xY
ObOenIofvw7yg1Z/JDf7bfuHSfzxSRN9MXcdeSZY+442NnhBeeCXw9AXeq69YJurGUfqzhnWD/cQ
+cT5kq/A5F8TWs/HSX0pfF+MB0VKpPc5v6uvV9PxD1gHvDb0FfZrXIrIiMon/6GQ4QZmfHF6TIik
lLa91xmWNd99khQKmJ49Z0Fs+sfJFhCqvJt7E8G/XwMBpzCCVQTZAnIi0jyCmLxyC5yJ6B/Tsi0A
RG5hrdyZsEdjY+jcixtr2vrmKfxYTZzLMks+cmrS3HrX3oSePcmdYBRSMopvPjl4Qew4hreuHYNA
kM/vtf/+NPMrOzdax3iXZlO4wmeS7hbdXg5HN0Z3jZXJoP0mEllTkQIWVD1oZbkNGOEnTyR9hMeQ
iw/H/15Rn7wLrTYywPlMi/xzdtIT5xGnjp8GYc+PMX2JCHwib05WnmUxRAwKWp3rSLh5PnMvN6CW
b1XY6eE6xZWtWhqO3tW2mM5VEWRYCtqXWs3bl0r7BIZDs4DPyslBFmRw8zcSUriN6fX7C2QcXZDT
qCy6F1NgVJzWcisnLxb9xQA5wz47XJDnIFd4xBwRu2Y0DckdfIbnv15OH9uCbQEif/SYleLy/Qjm
q24LvVJqtpIZbOZBKyO4RK8H0kFDOz4Q2o/5kfBEcYnocOIEO59XdoOxdJWIHi0NYzVMLw82TiaP
dPZtKescBDIjbOCOjM34T0vr3ophiPfsHsXF6jeT9K71ZLxZltEI2BS5SYNmfKqzXh9oMVyJRxob
U3NH+n9Ex21lTqjusRWemARcTALERPoQwJN/NU1D9YZCWxzkCE58OH/6scvARNtxQ5BGNJ1BOkPn
TEj612AzQayZd9wC7kZy0E+6vVC0xoiohs2CWc2m5t2dTBVx3h6wUnleV0oop+IdFSSCyYoJPmQs
Nfnf07kdUgy3wYymDrydARqC2h7WrdPyEGIENj2NbExPBjR74FBhdufIkc2BUbctR1KARabhIeEF
KpDe0tXPkbolTf0FP/NIUeCumAdjQ/mDwqd+imBxokSe5VmlZN2bOuQ7xf2NjHccazJm6/btIROu
rs5S2pjnkxDQELyBt6Lo49uWgEwuy6QYPV6uX8VnfUF9DoZZtzhr5YBZxNZp6Sk4Xs8C5wO6U77o
+8lmlPxSziTvr4y3/BHVVQ/9Mnotpyhpt2JYglwmytctHArhVL40zvcoH7YERVeaELr4BSl0WPI5
OGI01PxdBDfX989m5u9ZGjoT0vBCyd7qv3thmm99X61ABk8k72RqnXEM5s6mL1C3F1ivm0cJWzeY
rQ1okc5Wx4yeqZZitIKoyhku3lj+CGZoKnujTkcBLHGZ6CNa9eA3/JPp0rEH8LZl/rPjp7ZaZ16t
1OXRjdLJJQiMDOsHMSWmTXeKmRPqVAWNH2nUke8GwSvHo9xqJW6Nn3u+3TruHXE7JVSVnkrKae5B
uQxhPYAmpDlrkIlg/HjLhnUc/tUJw96td0WVkteLC3E2hlYNpyYehH5MYlAH/ERyyp+vypfi5AbD
qiuvneruA+7jW1dE/HBCcymLxuNEEUyXgHZ8uX5BWQuzMJcgh2j4nh4i5NsrpaJEtD9AxqndQ/AA
PGs/DH72ch5lZYx2FfNEl3meodBnPY/36ItYlxQ3KD+oD9u/ZSsfdy1kMZkWmibNArhMDFOuZ/hn
8knyH+PgDCIgFpTtuc7pSm5bDHkIgWmwmU9CdMuBDKWnvi2DhKTKkYCLa76HCc4ILAV7qh3Ffmqq
02iv00+HtXSzorgrDX8upiBhQJucFr9RDikW8vXY7a5VDFJw7K9JLv6bfpR/CKnTBin2UF6y3OfB
K0B5GtxA1n93+BcAeyOmoXPqvFcDeuT2Toqa6t1CacCLp3nFSC+xJo8GTRB3sCU9B6PZWkQADjCn
1DO5sGVnc4PLgq+v1LkJk7VvxeTIZOXmKessXMhpJi9QlNC5JAg0zJSYsclL2cSmspCpbAJ63pwW
OBQFx1kYu03rJeg5IrDCSrwFkNp0AliTHheL9q6z7nLCrmv0AG9pVRQDYyYYvf//Hy8bv0ZkLAVE
yUkEmmqah4svKxTNAYSJ2JMO7NeFtw7G6Eo/DaQnPZjSFWbHm+ZkhNzSYFnipNNn721oc1klZthU
ghuhZSnF+6/ZQdig4f0dFb5zfcgH5lIZ1wqJjq/kS6W+xBGi1bigIXV+6VWxkWP8YXYaWXyu/HXv
AadW2slSwGIsnamoqt3E+ZZwUdF7QJXN5Q0Q03Q6A/+eIP8sc3wfgGKUWwXM+7PrKOcjIfOFN7a5
hSnP5OZXzpVj0K9mOtkweEIl//MQAn7xjXTItcnbovWThgcIzs4bx+a2Euq07ijxrPj2Vrd5BzYQ
zVyhZHioiLl0W4TK+H0cYRUXdIAEmghbzWE964U6CQXL8SIiClN1paxasz+sgA2t8EIk7EyusIb6
DAr6TTgIKyswRiqG73t62WRBSOhqqCG0pFMP5K+sBH+k+ifF3aXjMVXC0R31VJw1CnmsDhvPKobv
nguhj0LEJPnjNqevt1LrFnXUYV6Xxk5T8dWK7DYAcxUAYKFHtOuSAGTDC1ty7gLd3xv3A3/pUuAv
IFWEstoh54qjunngxZlRz4nXb6W7iaLDYb2DAFAdQXh909awH9y8eDK9YrsKRdncQP0LFu+irAZQ
0x+tVmEWPYqV7LlxXNNPOA+18Nmnfx8LMBqIn1dzjwJquzq3Y6F0QA14/fBP4f83kkHwKrD7EICj
MbezJ0hafaTU/p00k/u7zFf5gVuMfxNH7ixp1U+11gIR6KJqJkO6viA5PZNbAg00/Th/dU/3x5K5
eOCGi48pUvrAoxdSlJd/7DIbvyI4EYrL/3PJ82wsxbM3hEgHRYPUVpU/1ic1d7T4Ta+fPrqNnQhK
werfQQ4uNT1lz9MXG0bADvAiMecU4hT5T1a894YBO1OSahPeu9befzgn+i+EqLOySIwVyOTQlDV6
oITBEcdzmuAyKEnywEf4SpEtuKHWhvcxCHzZOeBaiTbDzOnXFOndaZ/Tre8L9zWCFM/zS6xJDCAE
DMcY/68pDt3e76ZjrOVTzH9O6hI+lrM0EIq+aXz4ep7CRQtT09J1hxasGNlEpEfxQ0w06OCqH2B3
PkLjpoLhinSuTiRpuhLsA5fwCzjDgaHtNRTAZzMmP1qQVv1g/TY01PXaNMTm/HkOiIl7U8EeUiMG
m5PCwJz3giuiVNvrB7IGbjmRfENAH+U5ursQq6dGvkgtcaE2nvfxRlr0x1JcjQS8qsmYllwnbAsw
P90CnCJLSfeP61TKoDJ0ePTjqcasloxJ45k6DkCux2BUL6GnUNW3oZXl1FG8YeJJnqXtKKUbHXzC
0OkCFv5uqliIniIGbWH63ZxYSD2/47TRELTkHG5e8AIfOfjQXx1FyuLvOpq5QmlldJju7WNOs2P3
04gYLIJ+ldQInXwucSGLRc1nM+D6cG/kMm4A3yS7QzP1a4GlErCPf4Z3v2knwx7Fk37lU6Y7j4LS
jse+XgRN2FztwuXEdbBRJ9Ecy/pCddOU6BSfASxBupqwoHttP86TmryKg202i03s3mrjkeDfAf/c
4DIMwTtEocJkL1ra3SoClzQBXogh5qkCHdRvlSf+b+lde9PLFxkCsiOu0Zw4bvIjK1YuiuUUBfVn
lWMO2hdvCNn64vpvDm6W+FrerCHItP580/gFRIhFhoaNYJqKUYqodNnVjGcc+gO2MUzHWv905kkC
iRjRGMO1h1rA/Euig0qtbk5dWO8QIbmUoT+UZCZXR0vgO55ZMUsriPK2bCblbuOvA/Kcw8NcLTn+
L1qqTjxI78sNCw2dhIitcna7r4jmtaDrkNsOlDX9dwLMx3uSkgUSmYCiOcngd9p9+2oGXG6gRUNr
sFcpsQGrVqUhvFPHATsG0GHso/q6ZFGnyMrmFbC6Ywvlz/URuzSy8RZ0A3ihJJCksozBWf2O+J08
FbWTFntPKHTCDkItzj3rgIBmHppNpKCflnEbB1J2lihSxzjCNVsV6C5cpOaBhVxShlZiQgByYg7j
PFJwzrVZPK5UVtZ7TUV0VA5pNjNlhF9KJJgNUKSxrdeA0EiRKJ2m+hus39q9ammFckFK+qOgdRwB
PvNji/xjG34rceMm7RjYf7Vjo65FFx+C9QONLZp83cS2R1j9tmiY4QGqnFASb4HC+u95stYCyqEV
K+4UkwyWK94oDGGIHr49aTeeONqTYF+6d6y1C+nktGJZAwAhcOVSyPThrylOEcF4tHaqowZsIqCf
3r6kWv4KSKJSGhhLNh8EBx4khJjPtHZJrssIC1o9EZ6mgtZcOyhgLd5Z1Md8Fkc26JHKCdsM+NiO
45rG0m3Q/v4iLJaHURZKM21OS2pycPiJZ5AGavzb1R9fr9tukCga0/rDG81/2TmI1QYettcmCVmp
Y0qiwdE7FbkTaam6EreQJCWOi4qBKK3SIOtrO6jbEZV+jfJRS+i7vre2Pf978Q4bw5aHIGbBIrID
ZcALFk6j2Hz6HZ63NfDsVQsyNBM3KsfemYMZ7g7Ivp3zYA2C0txvKBtfQLKnvMcEE65NtWiMStbj
QMJtcTYktJyIo4HcUaNSOHNEKVAxb0qiKCyqVi4S4Aq7PD4R6HszhPhbMDIkm4g7Rtjg/ENSSCR+
0zrmySv9dOWG7pgC3bMJZ/yGnqwBJkS+8u3ArrejEgQQplU32SovKbdZeI0/74Q+O2EO6nUsG+Xp
rzvMSOdq/Vh+elyJWQiEFg8fZgen7ufid5KSNncjBNgrGbmyxQ6Y236WKG2qAvAZnlPuXl+5aXw3
aLhACCVP8M5VMllNVWiD8Om1fo4+1JTKL6wnlFQX1aac1T0NfNcLxighVj3izCNEX0/eFwuT2Sb+
165I0rpaVL4g/3U++p7YKXC0yKIpsE24fAwd71YLB95945deas1mGJS8GJfhpo7ErI04mYKpc+Mc
4j8vTTa3bDv7NoCK866CSUdgWDCAIEFiyR3uOVjPNBoVBhhxDz7TnXbMDmvk7wd3IKTgkyN6ZxHE
NKXTOkrLWq7GAJTyOyQ9V5jKanLrP4cH2+usv7qLJwS1fow1CNnkCelOZqcXmmLWrDG5Dza30NDW
miGxA7CXMtGbsHZ2cX3/H5s+EoJToFFLMpWtR2nDnGDkzkLPWXBgYK0HkFGP0tJulYjBIn62JDR3
evZHybcmZ2KTt7YumIE0/+lnaNjc1wINBVWBF1o9k18uAaUUpOfHnO5oRxOxqtRIT9pXiHmOaWHT
+DaRqc0BdSqXehSRTKl8SYOk6f3MHUAyZaBk6by0iCqnIJSbrZ25sTx6vNF1VVzqgR+4/2EZucTd
oy1C8bgP4BitNYrpLyb+nwqZWY/TG6FQduHz6lTem6Izj3dpPxlTbE5xPvHqvMn74c4i3RoqR/E6
uR3T+oZ+RsCMlqhQDJp0xj+qpn0M/dqvwbMwjaXIwqjAfLEF2jRbwBCFu7QVwbKk326a/m6dpM7e
khK3zWJEX7baV04BPIYwibvAcaQqaBBL0c/CTqqfpjGJWFYP9dARhrlgNyd7/mBxReExLHo0sa99
I7SlxCljD844wiu/RRM7/7jS1fI/R42+wYPZtzMwVmozfrkZMEUR8mjknqcdbVlTM6O6Fyj+ZtHn
fx/+BZxkrPBPfJKagd6q3AjUw+5qePHanl38SVy/j+bQFiDN02+cbaNOfQF6qX5jvLa8TPvOBJVP
SeGYCM9HMYvjyXBf3RFrTOEfjXUeqDfwvtPXq+5ILLf18H9fGfMK+95AbmydWb6oVb22Hzy1AnAL
dfGJ8WNFTCoi7ATZnsxMT/GLkcsGLbqVKSdmPQSV+intxpWyDdq1NBy2PYTa52I4pj1awysiuCWU
L/0UAM8H/nD+G0CbO3Ie2jOW+GUGWDVqW3ouJt9qY1P/MlMro0rBLA+7axYVUZXhsk3i0glObBng
kYkUFQN7LzPdtU/rKG1Z7xfb3FoppNQl/8uLjQAxjHVhw1DOjwlxmMd6GRabbtNH82c/5FnwpLf/
DDhpoi+3Tdu9RzMcW2U/DctoC706rhyn686PapaYE034TAIE3bjxGzQgNbBDs5uHdy69K41cs4pP
ClX+EBklgPyHdfLZypHPw50sxdgIBbHpsS9o8/H2f/GsmVnfY8MVuMZWleRO5KJDb2HL7rNJNC7E
JJOxhOi6JLEVcrowyF58ddrB0w8vVW+KECNRPiug96wj3PFWggSQ3htyXrW7l4Du9kxx8PSOREUl
C2xvU9HLBD+bUoW/dta88dR4bwUWkzMWs8Uv2cnYXG6jl6xISSOyOgjxb2MYqr7yxNoF9UeATyz5
/ESjyidx3hJwjDr43ELBAPgsdJrKB/qVuNorcbfKMrScZpkZFjTZ5+YtQA6G7svaruEUtyvrIgN/
FrDXSGZBdt6Shc3j6ZZ9mxLl4Airqr7QpoqcSzelNtwrlYewmngOF6p3SMmMCTK6XkBc32/vhHWQ
d7wmQVCW+CSLhR2jxoirv8XVty0nUqUHOpCFqB0tOU/pS1yPgtrx/Zs/VYTjDQyYi9TWKN1yJjg4
tZpGOcAq3vuzpZEUZpHTv4pqXHvlYSVpuuDRXg84014e+huESLfZQLffW+gl+keAMe4FCLnbwNPw
4FRVASKXPmerhJ+uYdoUbKxcByMqnRV6PFuJGQzvYtQpsOqFINhttyBeuv6zTP3U6DWX4MeAkBAy
LHYytT7DYLH3sNniOdkutJkPOz99FNgjlb1uVVght9T/XxqeSfZTQa2jR9NygBCcT8HXw6ecAB2i
Gf8TLF7Tx/zenut6veIeiwPNPEaEvQrKXb3M1XDB1SgGj5KIN5Msc0wz9hc6Ij66DY+5mRoHxIC0
rIvwWZBPNyyAVIC90IdrwefzrmRyruvEKmQ97rqP2ywkmfS3yzlsA14Qk1+XO9LDW7r+R7XI0uKe
kxffd3mJIGC/x3X6LEcBTaKZAhkEv5IUsIfSEWH5/IWBKnUvOoDuO2Jcd1VfQD1Zkw37KRetExY5
uo2/JPDQFGm+YfGAvzKUfbzK9oEawZgUqQqXWSHr8d3aaAd/Fwp/RnHj5zYxXjfg8X+y1sLHEvdi
TzVLgszdmC4rn7+OotngQM7EeEavlNCd1vh1G5+RsnAAIzL4pPkLUf89EYMyBBZPn0GYUiNqsQc3
GvzE8kD3fSBC/aljkimCVnj1b6Xq4kyGdZTnJrQOABoDqN861VjETpQJ5UVXrl36T2N5Xwvf5qRO
qUhnm0IgRb3bDlLvw6OkBI4vr7Bse85qgnlcOkKbWpIr/rozQzbe4mKQM+qiCAN+l3gYeRSe7r+R
JFpl1fNFNOxIhxKO6Y4T3NK04OuEVm5hyUVHVEsOwEaAd+Jeq1GxLPvEPlzaY3kBQIfX7+ZGCgv3
lXgYWPJ5cjZm7hWjCNn8pvnyikXy9anYs+wGruEd5K43ytpNejyLjn+9xNn820/7P8zhW9oTcJEv
D6ic7whM7MNe9gTK1EZpoUCUY5m1S23DLkPQtf3i+GmsN0X4oYiea38igynNxtqAigKZXwjX7GUH
XicJhhpGEhhgKzDVBpstWgCRs1yTHOweb1Qpql0EO9K2hJuzsIX0v10uTcZPaNqhHrdUclPUML8E
ewTxEhO+uK+VlXNqQYZLG+HXF8BaUidjYmrAtv5yJ5floP3tqKdbyO9IEb415F2QyXrKXM//DCds
j1/Jfkmgbeyj9Bv2oYk3mvmggSBtEgl9ekslgMT9QQoKjZHSMIAkl2rVlPmZb4zNwDav49JuRKCf
/EoBb3Gq/1DxZD+gqZJ6BP9bglgVGLkWl1EHhkdrX2edSO83TKB9TaAmM1NXFcvS0PSpO3mCskBn
pBQ7hkb6eHlpry3r+Px6s6DyO7McrhGlmzaWLVjqYR8nxt/6Ias8kXVt3cFdASlqkkwQ6jcYtwgT
5IbnUR3tRvgYXbx3Zdq37ArBJZMQboJ5rq+vI+4WBqsrYQkVHKuq3vXce41cDowH370lo1bGRC6i
n+CYoZUr4h+L19ks2rYwclI+EeirQs2SU/XuetlFMabKzfv+17b+i82Ktbgjz8NivQjrl/jEmceg
qpmFA3BoyEVQJ6fknykAYEeix0TOOzEmJLYu/tB0xE/NEiG1IWmAGqeYtDq89peiQcUM94YLy8FX
IHQCVaO9VxpRIItlZuK+F3V3qxV4LjfUCWAAklwNp+WTFOI1Hdj+9zdM2vCm27eas3ksE8l3ouPQ
ojpgxlwo77KmRAM51GWi97/bkLYAQGjSf2h926Effm58BMv9N0FDXY9oA+ATw2sOvT5xiyD99VDZ
LGKESy5xwiXXSu91BHiR1sZIaxrgwIZIn9I6XCWbuF9UZQzDZvgTWp1guObvgdzcVw9DFbXbI0QR
mXh5EGtBSP4mFjByT0wKAexnwvOE7dxcezpsQFoNZvyrKNb712mbwzNmzAbMQzno91WIaS3rdWPA
+UpJSXne1qaG5xilGD2OWKjNq+/0THakBme2YjYN9MSNL2mRdXoA3JGSVmJEoklLjzZwh8WhHq/T
vHFb3GrdKMw3QYe7wC8kY4/9FguA+r7fqo469uuEGhfspLavV+/I4hBicj4UALe6BDUOKksiua9e
38RNWJBXJ1ChhO+/gGVQGDKrb8mqnxSnOUadOgl1KXCoHXhe5orRlrODaHYMX+5jR0J5iysGSQqT
59vrZ9Gf10JXfys5ooSkYRZyk/e7oi8H0N81jd8CQTdnBkgJq+Bo0R2kpZbz0UDbM32r+NnduQpP
m1sIRIxxw5uB7goQKcPBHoxEdUbX/IjUT3xjrahJep++pzy8UsDdQTWXVztqMfzItsHsIR9RE8oi
W5xdLgMZXzA8DtEOueqf51wAzvMP0J7dENP3jSJEpS2OlONQbD4RscHGXu7LSavjwMRdgEF9ADji
MRFrKcweZYPWbvGUZ/mOEFXwJnCW2qGVuiuY0qsr0he4pEsczxTRxYJ8nJIIym3rjo0+/UtNtgC5
gfiPWTAJxAUZ8pL5hT6Ax/EivnZxqNzXr7gMFXEQmpOJSj5lI8uAfZI8MlaowXT9elHEYxtT9v46
iyo03d52e4QvLHYYpoLsR3dfFp7MvKSpMuJvFlsI49awiC0wByDiNnORv/W197AeO3uFYWTsYQ61
aDYzeIKSvN6XrOIdPM0u35SuRokfhOO/YHYeyu5EKrdhpI+brnbdVR/fesLJdcH+y5eV6gI/0WLo
AVoPXR29+1YNhisO2i8dD63z2DW3hzAagO/8ZdfKknENjmao2iu7H/LQj+dwtN+37XKTmmzZoKuK
Rjtr50v9r0B9/sVzSQwMAmU8LT5L6jfP7tekVmKwX4qK5Yzncdg2KGRfuoFol+Koed0aabYsUbYz
EvFxYHVDBE1QcY+5jTVDe2y2Pve03zcJ/q3EmcwW7lyQ4CleG0qPI0fQ6E7zM1E7QpsZTnFMzYDr
5hJiel7sHbmFrHJbsXvjFnY3ncB9nBMTQqOrLG4715MQJCkOw1p0My/O/T3RrxcxP+bDXr3qDeTA
Z41jawnNGXOXC1RYMgDE5nMJSP1tUaiweFpELr4HqiAt44sRT5RddfaHbBnblPg623iSo5txVTIx
enZ7x5boSRnglveKJ1j9Wq6rQoKQ+gJ/0ErCoavRjooaep6HGcE438zwxAGHl2G3darKFJuAcZNp
VxojVrBartzfqyFvNm0qTu0ifw40IT9mVdqzJGUB93L8AVDvDiwlYkShqfeMi5IM0AhJCNi8keDz
RiBF35rg/ZsvEwYupmdWVsWCCPgBnQaRVIdBb8mZMMmGRwAZxv+2MWHr2gUraSbNih66TiB5r///
mUj+0HKwxHH6Y56C5DDH7j3x4NXqfiN5ILQEvEsvt/9yFqqjFUk4DyGy3AhvK6NU+WVZnA5lmw2v
bsquNXSul3zY6WIidhYr8HsYYby+gymfE8rFenWBRlZD+viloJE+D+WwbPD2T4hvwjDKTUNKwN95
7sVW2OweT9fSW77XmCy1Dut/AZ8haXOs49Jy7tpKCffGMJNu476cFSlzcln7yDbKYm22t8KwYYVa
Y8PeKTQPumRcN5hDzyBKFzl7jzncujFXHJgIfVgcAvZ0oaBbNR/Ul+zELvggDL5CrBhokfbZQx7X
k+MYCSpQxrICZKDcO85i5InFChlhmxggW4BaYIMu+Vjj8V0iQPgvk7hc1xoIfyxbLHmaHG7/SJhF
qeeCdqMMyMNBR/CiP/dcJyXWELKZ0OtcoUJrrxOmY9kWE+65qrFRlRa0QUc9NE9SqK+qSuhWc3im
aEm334e5PeHaMI35YazBQnCdWeALtBRD5WgOMeQ2SkhskVy7dntHaify2HR9uOE/N+A8BJqKkJuZ
7izOUkM849y0V7rzdnMxXGQkD4V6XKF4j5wxMxvLLhHv3J4ZcU1V6WULhdSmzj9afPDFX87N2R85
zdxG39plo7fy05LZnvVEa7Ld47zKtPTs617NO3HO5jAMD6mMUusJXCjvPRCEX5IzrTaB14XmFWhp
Gqxh8G14EDpYFRar6cmJiJ8vxWIAclA8NkanoT+lE88rENxXMQqdO3ej3yf71ynbTrZ12YGBSJmL
rPfNXCYeOpRHq5Yxw3iSrDwSWeA5ckTfcwwHDn7RI1ztHfDMG3h8fE2DU3ZmH1L+6gPSPbott9os
MTIDPYiogquUmmUosy3zfx+NA5Jpb0+fGQvlJRegc0fdqnO/juy2m8MTVw7qntYo4qzM9oQw8qKU
/ZD4kkX0Y06ZaU4CUIkB6c+qW26bok6QA0kgjCQ0wxR3ro77n5srQW+4uXVnACu1bJSD8Tb3Q4dR
nmrekfvC0mhjn1y1wdIjdc0SsdcGBxNpjE7wXjjZIc7MfpfKaYzA5ho7qPpbbVvOchCCewPAyZQL
VPFD77A4MTktU3nSBQmGWdf/lrT3PlgKC0thY4YLtU80SAsKGQJndrSpZX1X6iZ11L9c7wOhL0Q5
2QrllTTV0FixhoWZHYW4o7LT1l6ue7NCVKhLhLY/v1lv7SXbHakwSn1G4SwIL3ntoNlxZIHOloYq
UvEcH1P61k3b5HLYsljeu2NcY5PHvPa+iwDfVGzSlLejK+RZVq3Qmyncxl8l4GIoxRPvUzsHKhZd
r549jAbu0KPM/6J3ljselGCQeRpO8bQ92BAF7f6wbxS9grI4krN5N78w/YEzCjFK95hHpAQvFx0Y
5mR4ugdIuwMswclqQzH3iASn+Avq8PyxTs2fcHWwdCDSG89AbvOJ+w5N6tcjFkXfmWbZ1XX5zdWb
ULO2pZwErDNs8HB6x96MkLPysW6EpldIpE97dcgzh7doi9zgdmajH9NhQ01yvI8wGFGnsh6W/N+w
FazwUUOwcuvSLoJzWhA2N52K1sZVzeOau8Xh78opfWRU6Lg2D/J+hUdiajHgoBOH2U/ED7v3Nbm0
1gFBbIgnJssFTaslZIFHowXpzh8YC20aYi5Q6sOXOzQKc5QtJCcgYzCMxM+Imx1ZBbEK1nIHw+sO
4aYTaqdDGXDBne0ubO0jxedpjIQ0Y/oZUfEvdrzeOnyBWJAKDshFARrQ2QP6aWXIKl4xmaaB/11Y
deQUmGluvZ/puZTLllQMCEyeY5YS9EbwWxav4Yp9NeuFd4qfsD8NFQVSYlV8nzcOCORaooabaqim
B7+sKjHEEBxYHLgAYyCgw0pwPVqMoeSx0ak+lmL3K5CaqjjvteDfiKhWUQ4MHYrVdI9lIrJtSxIb
hNFi/RiYVQB9NQbVXbXoQuWuRF8UtFWu94LbPe872mscJCNulFXGCjm2aLgjDl/IZYmMKrV4TKFK
Z3cupz2qIKLE2tlyrOHIrLzsFK9Y+vm8P+xhDbFWO88b9tBTCXv1dDwERaIdFYy5+CoME4rQHvmA
8J/4lMfzrrkCRwayzRhBLVrPqHIxWxSoN4UpE6bKnjNHHyle53AWFiQC43GgQbteMkKAdz5sH409
Rc5js2BEK+YZX43KwHqqj4hBBiSV5hnhBT3QVEo1v7NPxu0GTnzgx07YJ5AmghiEVdd4I2BM5ZVE
E0uKZNM8lh1PoxA9ELQ6lmVFJj7y9S37YmmEIM+ZBgyz0Ml59X/d5+2IJJkNizg+YL3grE1j4lWA
bxntmMxXZSL1aL9sEVvKCUZOHRXycJFKPjD9fNlns1a0vv3CEUIsqOKtGnd0HZ+e5FmngGgrPiD8
xCmpe7+umZV5P1DKSBZaBv27PoiBLA0+gkUB3APQuy/8gHqD5LRBTvFOZuDm8GQ20HFIyw8zNE9b
cXgQ2/cc0T7JwX+ULR56UEvf65TXSY17C2SIJW5CndMKRr54j+c450JJUxSnyc7D+6oYKvxm6J3V
iA2UDtBKuuUQn8UWZNB+fPQTZERKrq9G5MoR82/LXKeILMN33cqlDGMYaKiYkMOTH55P5KUspuP7
sSpeSH0yx+4M6c91VBQjUrp1nvAufzbn7b2CVZZvdmWMvhOBYw4kDsRa2qWR1OjGeewdcvXrzR5T
HpC0qxghUl61OpPZLTNc+cEECvpU2huJyMvNcODfy3UROUZWeYNh3EGKCEmCWYebuzbP5Q9+YURb
o4z86q+1swZ8PlyHE6Np4xIE9QBCwNcJakOekOH3EH+W4qeeFUs41sxEURTT/meuz3UuHWpDHU+L
mwiOsZfI3u9YcZ022sTud4yrEq+h3y/nUsDRFIu592RCTAl2jQwmuseSWRFStD+cHcOaHqoyHWWP
uqTPd4gjjBZlxWEbcSoyOYToVDTA8nDGkxrNICnzxdxteD+mEq/e/5AdaZBoTZU32zKwgwzj5dO7
G/DJzHwK64nK54DprDfpn8QR2JmzibGA53i1tQWH5S0NS59gao+5j6LvHga5wFsnckHvy3s1Izza
b36bjTJzLw0s8bt1W/h52R4T5K/mqcdrXsgZ1kVdzdQUwQ2MQ6TwgIpg4T5BZyPdYP4ZfD0tAqwJ
8nkbSpgN4WJDguDHpgYBWK8VNem/AVnrJP9Yrrgdm4uPjCcOdtchr3IVUhK1CqN0Uy17Zf1RrOkQ
P1bdBW4+pOP3bDYdWHnjyHv791XaH8QLr+M15CVm9DJbzapFSrOEP/zBM0FZNNrDNCZ9ITELnZbR
yyiAudTjz/XqBPl+VMimmjEW/ZwePxgAlDy+yVP6Pe3fkT9cbLGv/EMGSLJbfs2O6ISEjBCawOW+
AEqEr7lLfX1QBAu8cdBLcr7dfBD8A8am5tIBi62K0ESukkeS6hDKtzU41fcrZvauBx0ydFZXKm8o
vPdjyoDJzltBdrHabz3XmVVsRYAdrASNouPOo2LN5dkJcwb+UsE0DLjUUO570bnwcKB/dWryppmj
o+WMsAJ0JEOhA/f5OQAxRgX9uLid5+UNrQ/uFKvHPvQyNRMn2oIgWteBO6AGHU8Q2BP2m/fdEEeC
WGh3O45rRASMFnOSlQuPQirL8DYFRsVrz/pVqkqejMFvc83iDotff06RWaCJH8vRqkhGX1hF7ar9
TFgMQ6hpSlwVszXXMhuGFpHpMY16ec1CJqw5+dp9+Lw66NGiIpycUVAuGafpFvtWW8WZIwQjX7Nt
xW+P4wekkg7NGnMiWuOJE9pB3C4p9VQgpEKUghdMcjbLC0FrmxXz02AvxFX1rKFeOjXKEHw6rdi4
nGnfOJLksCVAhRCO66pnmi12ii9W+Kbox0eJ4bS221Se1B46ixGhDQCVQ2qV9rJjxjjKVF53rlg5
N57t46M7jQob7h/6AybIX4lC54PVm5V9XR+wZbV8QcLKsuPymAVeSGmz8M8X95x7zYqCwNnV0F4s
coxkt3Vct8CGN/CvSsDQpCR0FNQi73Iz1MEURcb/RHmFjOjxmArDvKDEP91ZhBgfAvXqGV3OWyuB
Qemv0d1FQDs9hF+Qa0U510QZ7be6/i0Lahsbu7phFxvULOTOHCAPYprjCFmrRMHANGQbG3NIGfnP
gH9AkRA2LYQIMKVPBqGkPVXi0n1ba3u82Z9TMY/BJTu5W0reVkNAeGKpPl1hIER9fK7iSgRQlF9J
3W9mNM5CORIq8dXQe9gKzX5PmZSrdI43avDLEbNN6pe05vOjlw8xxrkJ22Q6BHhESMKIlNfXXgpg
A1cFsFyfH/gi9OH6KjSKmJCetYmWbTTXsrNh4mt+kihfzT91swwg6XA8Qsiogiec5pGCuquziAue
klx1n3jWC0GBYgqJ6NkVzihVCaFvsl5EltK/mkqDPAHCAYj3DkE7JfwySUb5MplFHs/2cHcE/x8O
G5fkFY1UqkrAAjC4jDf7KzLu9IEPpfEA07/ftwlfUjJenecrX7nC5g/P6FAIEiETcCDqOFg9G4Mb
d1sHJKQkjjYVdeweRzlOK1Qc5yU4Z1ndIHkCx0Lb7c0TRmx5n3c6KLlwyjIOvfvlUk5gAgpZk67e
v3FtxsUp/5EVG4X996jVpnKZacRckb51Ery8QVzZAQAv9T4FQ0O8/isfkEVyr8fdNl+l6di+kMeZ
i6fFnd9Cc0SrlFLPpWIK839jMkJvoDR/4DeM7qr5kDW4BS5Zogt0eB+22b0mp5oU7w/vmobkeXCP
HfsOXjbTzm+Ys9gL1fIA7cATm/J9hGJds00Bwi9+eezIgxTJohyDSOYA7v/O1w5+WRyk/pfrIME8
r5ITvXkF32cdElVC5pAEW5j9TBJqYMHrSShQ5EqdqwTWE6s1zOAYMVG9BnUmO57Yebxl9+UfCLde
s1Geb9g+5mJuL4RnN+pUtyGGcfw2aPLnThLuubqpTI36la6PA1P1EYFHgt9NUGUMdiOvwsPFcy21
ba3qMBLQxDA2y1aCy7qFbbYAIuRE0krdadoY3nffoQbXC3B3xKIsG8fDYy4d/WArbWQ2MqlYfTN8
Kf3mN2y1cKxc/AVO7dRSSOmAFdg9FIJkMa/RRoQDcKHBjXI+wcimMWaalXqGNMKNcJG/IA/ixAyf
Strjc35lvICXaarN9jDd1IehE3VGhnz+nt2E+LbimdNM7vskuike42KjFZqsq3riZIvVfyCIFIkO
BWnCWvPT4wfJi9SHi+14Egc6ckR8hnnMiKRRc9oTQ1G8qhq85K9LpJugzJSB8r2bQsgn2fpB0JXt
ZkenEWeME1GDMVhOT7TfbaGpm7cgS9yXOtyAjOSfZJpRGpcjsijfpxDQdsiINB6fwja6jC+m47z0
71jxj2hzi7OhgTqbVVt9wxUU/l+X7Se4zp96LnBuZuw7fSq7dllbFgA9G4L61wmQv/qV/6iLgYmb
ix4SzsvUGP3ek49SMsTaIxVGiYITVMepChMHbgwy+hsWbktCf9PXtJ6jrVChPGjHVVsAfLgOpVDR
mvPkXtDy54XfDtq2GUF4KRbOTXcbHUGj3wQg1fHdMY3kYzV/n2moUihIK0HEBlvKIMGywUXeQrCL
1HjFvAfzVt8I83s2J4CZaa7f/s0hVtVK1Z3YlVrzO5/ZvTS59mnAk8O/rWdN19oJl5GzBA1CybiT
MK8IsKp8tOZ6XanlWty9jwf/I9o7UNVIZybBmJEtMb/f0mEauVj1MS0LI62K3X2cDw8CkZ1ydNKh
CALd0Zqk5TJRIj6Fhy8lzR5qeXXnepcRmzQcjAinoRGBZwN+2F4VChJyXHV5xHpG1t6mDf2w8S6j
Edftw01ba/LOZtAaWubEfgLLivpzc1Qyo2Tkb4Umior5kgCE1Gs1IR2NsgcFgOE31kvYf4vb7qP+
3wEvdJ0lIEtO6qm7bR11nW0/cM7tG/J2Opk1o4tr6UY8dZOZI6ff7u3TnWY69/NH0AqRP3DrTTBz
ePSppHjFCO5c7fcFhemNtPf/pVzhtu/6sUoM9UgMaZ9PGNxZXqDXGFDConFsUQ55XGtAcGzDKx/t
egSkoCjJ7b0iiMA44J1Fv9og215yFZWcmQspPSfiGeD2w1vwn4YlyGOu/b51jUgnCetzuiyA/wlF
8bQ1/p34NLIQvGNl3DQz6MFa9cKEKiCjgSmK4rdOiHHI6rWTCliwxjSmykge8FCn+Qt50UWAFJzy
mpqq+RtCDUyToc29tFfaIIW5rUdPC59JYNQY5KZJLn9lSV3RFuP5ekVctHPNCmbwFh9vqmL5MrMS
CylMxrcBF+YBbLRmEJm+GV96dIXFzUIR8pUg5DFhu+Rd0I/8vdy2yo0oqStCAb+VFy2jWHykO+3V
Z0Dxs+aAEl8P6pcpiL4huGu4q/OFpr5njN0eFDatsscViOMQf4JTT2G6zmrQIUVhuKLfdkgz64ne
ujq4+M5yKns//AODGZ5Q5wSUh5mhpMNDdBur+8QNPuOGEpSTfpA+dkAtUlu1gTIyeXGEd/rP7YrJ
KlUatY3j+N/Q6ppwQmTVTULxa2Oklo7CxSimrJ0BKiBtZimGY5EXLoibPV2OfoDO3Q2g8lMC2TxM
KBSREkMRhldBw+dtcOsB8aL6kvoLnmmvMKWCemO4W3coKc/jFnKnDoKamMWMzTYS5QujS/LyPi/q
QrXLAPhJPUhNAsI2MrKn8+5aRr91E91N0ZAONJywmBBt3pXnvC0IVoaF7XKvgCJeOyt0cShObSqZ
ff64y2jz7g052zNkehTdEWgYN8BMad2TS7Qgio1QrV+/WFm3g1a5rvx76GQsr68wyrFGWhSKCUzZ
RXBR1RQg1emdH9sWrRGSrct2fZ9PBHXys8tsPqBVTMagy2Kq8V3qxiQo8C0gX7nP9MAwu14J2an5
NZlY1ts+t6oz/aJOWg+JRc9lF6F2Cp5e3pCmM2eF+8cTHyTY3hc4V1UWtLu7DTBN+RYI9k+UMwNb
I1iEfSTt9OwENwp3k0PzAJdFMrx3u3wMgD6fIlIPKDJtK6F4WYhYNwBmgqonoFfUqg6Pzf1wRn4i
aHTJMW/K4fMrPLAOTDTuZBgv8HK5lRKcxycANB8lDfrprjZ1WPPb1PZpWr5V7jJwroiu56iGuVdd
b/itnaLZWWC98MfEQtT/fVbt86O+0vEDpbyDiswpSx1lRdmgBeJvN1/PIaHVsVjiQW/JEqiv+zEr
UoucjRJbJ4I2srxkp9RjY4Lud5byPEb9F0zKmPQGKV1jxFthCJ35nSXF1BtvPu/7bw73uXGsAWjW
61LHA0QWe61wmH+sBqMjyxrOMppaJa7TazJqdiZax0W1LDxcow7FBkOCOMW9QdqeJsETEA7dhNaQ
FdqM13iAqHMk/mL9WsFSnSdvbfm5FAvqzo1+o53Fo1ZM/+nHE/ERiT+bkjkUjN47d9PTrKx1KTi7
YI97cvUPokH+rm+g1cJnOv6IXsJddMsR6xDNf5cyKydMGSDmkZHsx6xjbU09BLy48pz/8cKmCNzu
TU7yrXyMfugp4pF+8b6AImZhPAWdszP12aRqP+EF4Yh/kAe2UtkAcG/PY4pO8uL61RMSp2EEVK4O
71gvzr5UxAQGMB+QlpXFai7zDiDbLcG2rH87VIK9oqy/+9hTnNL1cyDeeP9EahMN8ZLIvdsHfma9
mgwS5SXnXpxz7/IX3idH5ahS19MxUqd+KbW3abl0hK9sZKYzSJ8YYwZn1oBnQz43cEaOYOZtCUoW
TfnILwcHCiQ0So6IT/R4BZRHlYbPMCEmYKeSeF1PmNAIZUldEUB6QGBD+kiL8LjuYYaJSVKqbZZE
o1dG9xYG8vSjFDRxlITKp3+oXTzdobgBgyRTMCyYfKzng2jfbbE99AGC2cuGtIV8QZ7n+VnqnHwx
mHsUkY7N2RUHI8nrGxY1Jxj6rpGSGAHEJW/ytT80lnbdb6fYCgk+LabNsCPBLhhMPY5JdiiTlQ0w
PdR6RfeHSUG2aW0izlU+NKxmDZReYUSYxlUMH9muN0Dnf+UGSH6eDag3KHtPOrAMyM3SR8f2Acnq
3EpYseJ5p9JclM44GZkMGBY26OOT78EOD2Rsz2Z/VGccColTDpNRTHGCbihgDTsrvL5deJMMmcZl
z7CqXMeKt1HIVM9gZjLrG+YrLLDcfiXZuj8mOHX5BOPg1dAcL1eFpUF3iJD+gtf96iahN/0+KBV9
LQJlBWQqQ0ZQj5JlRGFSir+Om2jIj7mX/iULlOxXxK24crbJJmxzlZH4qpe6LLp4/yx7PkFsWB4e
r3zPo7dkSil43ZxbRRqnv39/ijkWOM4swOuy9WBYhW84roJjf0w56NmNIANfR2mzAqHX+lhWjhGJ
fWJoRTieMVnnyb61cRW5nwb5q1fCoCtX2kK3IGOZbuLu10W8lSXPhQm9N16N/VEf3el9gCJb/bah
++bjBZfrp7mHiWAh+rU3LR1BCXkki/+iWPVrCVo0zWFh9N0RPB6qeHKuCQUtq0zc8sWYWcMm88rJ
rBB8Hx0g9K21vadLrHehqF2XAfUTtFwBh/4b1ae4JQ1YvSV6Y2qmHAFtORhl9qspgR3KQj05KuXW
Ev9cIhAiy8QyxZD02rhQRuPwGNkmHY/EwHcl1wpMxnWhcV+Rn4ivBDiuNQ3UaNRgWdtiAUvYP71r
KQZlY6eGxF0x3s951JVw8vIXicAR9XVu1P0RNaPukddEhIDGd9Jkj2sEqR6zfKtphSw6vQm8yhJ3
y7IHniyQ3YpJYA5NgruXyeQO3DfwLYVakaz+hMBifglwPyPckmhv0AlI2z5JETfjg1F9GR7f2+kz
ETQKf9wy3RyyDBc1D2YJyVQygvtyYghUp3JsqfvFF5JgBqpoUhJkMssT9BNdUIWWAbjLt3ogLFtP
8iLparl744UfleB9krJzGT8WD/DGl4dvKcbZ0OdGDno5O1BvCDY6w84WiEgkf6VmkAYC3Wy6jwti
rny51v6htJRrZ8YrWXpbPO56h5Q0Hxkv1B4NZf+BsulgBAdXOLGvzQHb+KZy+LblxknwP5abkr/N
/YM1HZOHxwWTmaQYWCM1C77BuuOR0e5sSnd0W/DwcWgsQlGvurwjPr5RobyB8atYrob2CmpkktgS
8Ls3biN+F5qgsCe6bcPiFBBmbtG30jy+wdiX+7zT/g9i5OYXXCVnb/Jk4fmS9pK0dFVcMvxY/EVz
jcC5tVVu7gSn/AKen9IoTw24CQUeeLheRs+LT8VFFQqTlGlev+kilNWtCYmgD2d3D7t7gIxTwTjq
N074ix/mB0d/Xqu79Tgqzx+X71Lwyc6Q5vlHrGoDhEby1Dlvhe8Y3rgUyWJlDzUmjRU817qIfN35
bEk9TD9wkAFzn5u2v4+n5/mFy0IIwTDfliBPWpPY6FhO9abTiULIv4465ScsOgxnBgHvBgbXPVQj
cHNIDBaq/b8gLAWnlMg8mazFjANxzP4Kwjnek3hiEpS2OtK4yLVTaTj2EmEPKja/tCCdQ8J6hKVO
JgjeqQJJ24mQkEQmt683qfwAWxi/cTrRGVBQ1+aLeSvgbUNZkJCBqOYDaRp2Idc9SD1PvuknF5Z4
YjueBJStqT5pyPgM98e034SpnYXgEoj0QOuPGXDRCI/d89FUofs0o69Wt8bfcHsE8XqOtjGeh+xn
xQ1kX+DuaXpWVWU+YLwm9g5+bB/QALO7PapMo8fqYgXSuSyBT8go2hBDl/QViz0YQS4CpGkqGKC3
N6SHw581d4sW8AaFHxipyDbqHXKunnGHipfqZau7JbG7iaJn1YwPmuk6FYOnlVnJGX37y2z5358q
J/Eeofp60ourz8lgAfMO6zKfcjb6PfqdJOscEkT+AwulnMZr+gmUe0f5K7vpWhy5IfhXS3wVF+ax
Sh1oCAd8GVqqknl0Dm3S12faxq/g4x826sMagsYRqDzlrOv2CsviXqqknblUCbTnsn1/qO/7/oKx
tVn8sRI9kogF0Ok4zybbQN2hX45v2vToQPX7T9fFKEoOLsYIxXp469RtK6Lric7VYfUD5Vit9K7X
o0EZsfqBK1dKN4tzYV3LjmXcKpbSiMbT2beX2Cko25FrxeNftR9x9SB2vZEG0mYy2IqPhYXyRetM
aNoH0vfvyhQmNIZxVXRetVrTHq2lA16LBRFSlaMz9MUsjN/nTKpm7jkz/CpGrNg6WShiTOj7DeDu
E5i5B28fHt4qQuO4Y+5UMtzsy+5E5gOf9by+EjLvJ0+iAWKwI4bFfY5ZyAaSWpAqg06RhxXzOQ9e
lB7PUVIR7vjMWVgsDX1IcgAbwjnOyWr9G/vqQR/wq2bONF3MB/PG9HnJkaf85kGiEU/tG4PZuD40
BXdWQz/dj+I/mDkE2b8+dSe4xYQh8x9gS3XBx7U+K91zpMUWlYC+J8ouAYDCqaSxjhPIB/OF3cY5
eOmhXp4VdZh8MVDp0UTNG+fSvndItT4f2k0lGaKRQ4xVmsdikgEIw9YEfA8FstRXrbflqaOV/pNc
nbo7ciliPTZzSWCjC9NvE8zi4Wi04do9K+TR5vcinE6oMDFZVT9ToWt+4sSyqWfepThTOBS4zCWW
2IjS6dw56tUoXc9BClbPnDN8eAm2F0L6iybs9vr015RhedxGe3PY8z6s9K4CQhZCOiXcCijpfD6O
zf/Swo6X/tYTJAfCtQKww31KX8lvn4Tc++lG9GQMH2LImldDg8zSRx5ev1iX2Z8Rh7ao7hV8GMzi
Wjb7OHzFbjUkBuKPeYNbXdcOu+EU+2q6G4MbY3LNRhjb69GeJsnFg18HwrCVtTtERiIdfsSG9m9E
hdclhUlWSOxz8MN3BFkDyJp08WFE/HEiRB2AY6QT07TW+cNg3DjXGqPhlOn347yTk/9H8kXaq7Ch
zirCN2Z8TbYLUZy/3Q7dSXbT23ijAZd2SGsbc4IadFdCWolou8CF5Uf0Mv71TleZLytDXNVbdtt1
FPLY6RHtjcaQc1Hu/djVi/wK99/FzOO5+jht/IJOjK86/bD9vq4a7MtZcUvXEUhx8cOAKotJIpac
UIreIPhdiruv6KZJ5aGzTx3dUtSkHA55nkcyoh003pVL0sWHZyHs8cgZhtQwD1e2hiZpAiTnwaU1
5UeZUUwa+u7xe4m/fjPBo/k08ePwdfdvKF+8Za+LqajrCOP+MY/PxHXuySJ2L7XrUSehuBikqsEm
OMoCnPDEwURs+XXal5/VqeYm29ec6egeaM44nD+qqoqaCpJ1fFYqgOJR/3XzsGgUUhgNkeVQsNQL
BXq0TtFn0R9RiwHbCiwQs2NWJxWyOrKxVz3phYbbvf8Tga+WwKtti3qQJKlFT239GwkBWEbZ8XEi
NOl5GW+iZmA17W3NoYUnXIdP2ZZJPImpcND+V3N3/xrG477jkhuB4RY7vuUuJ+Vl4reCzJtAjvnP
A6CsUCZ9JYAf+UHIEoWYVH2hvORWlXc6cKvoyTSXr4d/HNFjYHR0YbxEifiVLk9oQ6hAnr5krDXE
g7p2n0BZFOhGtPOJmgVdEi3ZNswPWCF9vfSg9X1mS0vekUx7cyPzFEmRkmKehrNx02vsuNqsurwF
pGXH3wby9XRPgISK3J3ihfnVxxBdnYcUiIZgbKoN1vgVPx7xDGirh3mm7I5eJiEFAh9za8oADASX
AXd9mArCsE5CG/bCqN0C/ZkH51G+Di5f5xoTJiQyXAVpjB5fjIiaek3GvRTP+Z0r0U3setbP78no
mSPYrYgArpII5CJbFtE3HXy0e2cUz6R0qPhPpJjtTNW6pnlV504w7D9RR5K/ChApdFfjuXst113x
bpVmHi39tG0kiu8IfM8sfBsR7hsqlR4WzXun6uHQ50xasGJZZ0SzY1BdrVfq0OiDvbjrxX6RJ5tu
nVJPDPGfmWgKm5g+9x7lKQCtFQw7Q0/JEDw4B8HGnRBYnu9kRrzxEsqgnh0STI874e+Sn6QtWxIB
6sT+Je98dT5tEIN4iM3b3D2F02yZH7tMo6dE+wokmjw7vdlDXm6mE5ndSlBG5HjuVVLLoikJppKP
JppVgOQCIpWs0vq6Cq7lO4dbK/gSGTJHuXP2tCp5w1Hs9ZCkDKokDYv9gFe4SxXDi16OT3VRzOaW
Fbp0tk+Ja6hqs9OBFS2NKRC5FbRCuAIucxi2d+HvJ1C1zE26C6nz2ZIpap73w0Ei7ok7tdeHFjJ3
oCbpsvc5QRUpcC41XDAfu/Eu0peQs4WO/Vx8MgaoT6TYVSNYmY85uvshAdSRysiP5eLrF+tN6xlu
rGcIVqDvveNmb5wF+TcAhy1GFg4PmmjZ5ILlQzaSKtKw2r1e/7T1aK1hx0olfmddR2mRwxgdp4R7
XSv3yYC2YH45E1EX+LI6fEhsS/WqloLnvYLSRQfzIEHpnZDQopk+i9+RPdxFHk9cq8pOcv99Tf3t
++x6kJVKHEl+FrD4Kly8iH5WkOjyOeKPGsxTAcTGt2syCp0ZpzeyZ0r+6eRdKklWzMK1ZfDya/oE
u2tPYvO028jFjwKQJ3+TLYD7KZGdR4TA6k9EUR2WTKQbuh/xjNvtTjSRur/00C/QS21SvUv1y5yq
u0C7mojQMI4WcDpTCd7ytTFDR8LYKrjlicn4jNkSW5Iion1Rwp769h69eA+RgIcw5AdUI0Nxni4s
vNug13CLWTVDmsbM9TqeJ6iHmM2iFcm4aPf9rK6q/3eWcte+8emSAR9wdEgjpeglXt4s+zGa3O4L
M6ysGKtVrVwMWHbLGDm03W/Eak40JDq4JI1Ch9/bWktj+BfPZjUqOFSENLxEd0m/UAtQnFuiv64o
Q8wIUGoGhfKzGi1VJysZMk67HsxFEI5Rc+8RP1WO/23dPSmFqo+jj4DrbGNjWzWRh+rOk+fhK/vg
0yC0vDGL3JoOIsCFgknaUco7opOy9qdao5J5h7sRw7eiTdfawQBt2hJhdcZwD70J1ERH7jb6etlp
b/xvke0lkqDVdkF2G1bRZghkr1LB7UgZmQHPDk0IgNR2D+Dtjf7EbJlZsYCSf/BA0kdtyEjS/X7o
kEmECiwte2lKw4WVFvrHCZAl94u9x1+00o1ksGRYQ64DXZtu1FkruGy74jaP2L8riM/zGsH8W/WQ
x/Pe9PKKbeehQ3sLNJQYZ1yPuOxdsP2ywBcIGZwSUHLrUefk8ttuT2yzAyrJ5mPPby+zIfJE28Da
OPPCifQbhAOnXsbBNSLM/VMAphBErL5pS1oegppGyha1heF/22uV5CyUn23sDq6tmyuL6f15SOWR
RHqdgv0UbMsEOBx2jpOzLD4wXVOaifnH5R/AH3PGFwk14y+nm+alTluuHqVWt0XOVxcESi1E0f5f
wC4lm6PoueXwY92NLLp2ncOfKYhd7RtT3zgx2PYqnvL77lgd9k3wD9SjACVzJ9G1jZkv33boH5kk
61JiKdoUrVaS9iVI5YIe4+6cTDlED/CJHNtJnengq/ThtvuMgJyxDuRIClLYCgLMhBoqFwgPv2A0
4+FUDNhSDcmXXxmsVNnlNklqJAFvYt8/4o7DSZxHy54o48jMMHbkYIlpaBq059/qlc2CGHYzdiH6
iYmbQf+DcNlJYMvfc7mUuPtANwvHUH9eQK7wuIuw6tOqIG3w6HAwbLmQ9nWosrrsdHVXSF+SSmw5
5N6/LOFB31hSlmxdLSyrk2zg+7cqqKufgAXeeizQvc0e5QOU93d83MHk4AM7aEgnrmXEv06DfMyp
C0G91+/xof6BnUjqLzuYrW3MNGhhpRhqT4Hsi9xDCX925BXk4u/zNLtweWbHrRvYaIUrJD1PmrU7
IvMDvWFzAjApf46BY81PLNr6t9Xo+X8yutemkB3fwkd3t/O4yrHEFVN5xhB2I/NEMFwk84f1zK+b
29P7WJXiR6XYU8JRGJ3wFgm8GHfClmMC5UWxl9gW/WnqGB4r1rdhGwOXjbU4hSxdWuBMr3w+AiYR
naDoX6n/OPeAGfu+8qKWwmQQiP1Kiqk5dSnbHoJ0K9SHD2AvytkU0AXRsEtNSytTaT8cn81hPwte
ycz8N85GdH7mfB0EzpXwOoXfAQKXc4zTxDAW+xXytozKVDOMz+48+VXt+GD42nZ0FDd3QClNuyQf
MgVR21BdqmaDOylJ9YqqeabVGj4M58eieauj993Eoxs3durTvDQXmy3uqtovqJsdtj2zHmJFrt8+
1jn5/t0xb6948W7EF1vYpnWN5Izf/fQi8FM8fwEGcpdXCM2Hcpm9BeDpJqcWEMBhvuICQOQCJHyk
nOewMEpOCVcue/cX665BDoRXoTNAgPPX5flXQ4HfX0VFO8ESSG3rRhSgvyUaO4l7PGlxO9xm4idQ
LHozP/giK24vnAjWt9i4wFRNkrAzxQhCoJrHmhmvwleYxB8LIjQ9akDAtv3iw8WTi6jSIiNbZ8Yj
Ui3jUl2Gt6x44NJC1mcXdBi7pTJcs3mYN+dUh+mqp9uiCEypeWY0QV53F77cTqjXKfGH4pU1TrV1
FafAbwXSkt9C6IcsWKWIXL6yyHJObRWLRTpC4dScYlYbJItEU2d76JCwB9hsmyF0Y5UorLQXhmEs
22NtlVgS7Q8hzTj2myqa5U2nLFW2YvvLWXO3zr6y4t62GhIlV0e/LBegcErwmtE2kZkMcWA87kp1
2sZfyRJtqedjn22/gHZvHkfbVBrDyJp5jeJSQwSoiNabQMgvk1Nx2grENB2Eqg0vp7kh1xQRJNf1
PJUCBuRmkCxM4in473PoC8aoaS/N8LvSkpZC1EG+PLBnoG1wUC9jYQlHKRUoJeRUsVbX3+jjvn3f
l7/EnarXNxdBAYAhQClcozUN5OKKE0bO2yM3mIVhzV5gLmay1SgKvbgdK1dEOroKz5vKtv76xYFH
b1R8nDHduegIOVpH4C+IYIweiQVfyqJmteAC3EDuSmu+G/m6mBh5MAcnKLWiwhFoWCAMXqEhHd2G
EwZzVzHSN+23fMSxCxu2wwLWAIS82eXhY7K5i3FPJlK1Kq402KmUP57Tb8g1Nc9wCR+j25ZUiZ3o
5FSNPpmYwpjYk5lwh5k/Jw87jShVktpQh4Su52LQl9Br5X03jA/NfREAQLgeiQBe6g3ZhGzjDeHX
dt1MKyOhcbg5jPAD4sJo2HsN+JIpV7xJpoiYNRvCvQa6c89+zZ9gOb6fWK5V0I+uNcPWu843fKHn
RvmqeyBa7zyLsK5xXFCn7ZFfKlggzEyVe50xMjOHhT67nueIBw2A9D4iXjaHTP3xEkcCkMBoGe+W
Vi+P7RFoRFC24AoGGzeT0JSpQWGF2fsJAUjo9c0lGRpjZCQ60w28hxuuPWUB6ZNVz88GVfATgtuq
WyWwOfKXvo/RU2JnUiXQK/zKoAgZ08QKj/vyxhQypQG7zhAyJcWgS1bYkULsALCH55LzXQdmuW8S
rqrhRcvu7JeTmRw0SwD5+VLg5W0S+mRw8J+a/4TUBPa/FL2+Nh/bF1S2mBKXlHv7FodRu7i2GZTd
8LIawFKVn7jSomUZI73e178RigSfq/oT0oTWMuzIwAgthMctioR4QSWG7m+wA59qMINvNWuAR354
PA9sHnjm4PcRy7rEhMI98dyRtZpoEiMUtf0+t88jvPu9+ax3GBl+8MXv6iXWmx/0ZMB0Pvxx5muD
PJlE3x9riCZJFv9PRMkm9Qrl/LLyxDIrRyu24D6tBrtKt/c7kjO3Zn+38l9BRx/WgEFaePooXFpm
93anKx5ZZtCnRG5k3yO6UgEnljAMlXEzXgV2dwbWc5ZBh2dQsOTWrQx/Z46JM3vYkai+wG3GOohf
lknFVKaABgUblyCsaw/SFRRvjwLd/NVFKk7r5XCSJD/RwW3tn5aUoNXP0uHP8iWMOs41qaYFKkiQ
ACLc1aLLin0g3v9Z+YPPHKoJiWjph9/RTUaY40qQdg7he0C6GtfbJmw5AyAYEf3oQQzf2az7Z/ux
WwIvPg1hMeaC0qRyA67rCQv10hLr7shscGkMeSGg35tfswtkeuK8vCEXazI8fsf4Wkmz06LLwQaY
xOxxQ/4eKz+Zdii53bIZCq/tLxgZ885XU16EqlxlARuxGk/SGHOYRHKaKQ1TSprFc+y6MrivKh9P
zDslAJW9P7dBy6LhLZzFgllEaOsiFuODjExrBnJqcs+YeV2+PH7qdK5TlxDj3IBTB37WpVz2p6hX
DH33axLCUpFST81EsuZxA1WvRs+OuwclefsujQJF3u2BGYbWQRogNVi8RDlvY5agCCifUkSQs10E
xzTasm5FT6sYHu5dtQQWGxTErb6TP1as7yP5YHOPzDVCTto+nrx5NzkHxeZPtq1A8s+Vd7IPn8c7
MVv1fTCIAlizDNcjmBiwWjVLRCbGzfYqqFKH2th9bLnRk4UuT0oNo8PyxU1mWNAZXcPV18QsXSVu
Yosg4wiJUQweXup499vrOjgFmcnVj8iZ6olCQH7Fg/3jxcDi3eA+C3Z5I1P7zEEbNp6RRwhCma1u
iTHFiZKM3XuoFmYsVMc1pB7U3SnQCLLPkbn2obYRvjHQqrbGpPd8vmgcnlRbKR/rpn0urwTtcCjZ
dSTkeRkafVx9/I//e3a+2aelU0LO4u1q+c19vXKkJutrr+FfZbRo71rBaYEOwpT6OJSAUkD2u3GN
5MD1YehuPXIA61zLw6DhbTIkoCgFopXahEyCXQauJDdiqX0S4+w3ng+k/xo63xGNdJ2mafF+aTnj
opydbtoZ6GYyml1TI/O6qA9llrT0F3dohA2GVHAmdwGP4JQ19pyvrvqUDnMx4N32hvQBLpyVO5v6
aqHAVxdZAVM0+WM2+wROz0MY2MOSiQf/lROyJxzp07x6HyKjVtMCPzQH137TzB/5bgwSS0NXVJ35
s/dG5lpuDoZY8KNAyELUQWN9B4YRzb9MxbY80MUbOr6Hu/N6eyXpSW+UrXi+XB/Z4afrhvD2kwCY
l/9foFAz/0pRZlGtuq3EPsmRCc6umwIrZ2Cs4mBnTYSB5JMdAGkH9qdC8AaLFvyCupSayZJWW9nb
7xkloPvZqA//YhfVqifeWM8SAtZmec0u45JgUP1RzWeuxm8nhNyj1xptiDTF+u89xWSeYCttejCJ
ywtb/cmwupx9QUyGe6atmAjetSUDHwFtKnxH1jHm0Jyerb6sqzkrSjOONmd5Yr4JnkQiLCM6DDcG
SeyRxbwotemRwlXheXu/k8zYItjrMlTHQkGyuNFFhExoc/ffa9jQOT77Cbc+fhgYRFxAZ7S72ArE
YOZJL24n5VOyw8zNNXgdIkmo9RSxVIIT7X/jZVEr0rBhq+HXQynzvHUaroQ2uE+SF0m8fKfZlDU8
MUmhVn8V2E8QYywuFilDhyPLh9H77UFjcB5CTJLFH4RuE11faLx6WFXp6gmYk1dcx2qMjO0LgxbW
QlvNF0D++gI1Fn6JrP6eG1f/7MAN2Z66B3/Otvt44bDhvopioPGuCBNpaLhQjrhA1mVL+nhK2CUt
IHwvwEOgDq7NJ4sOYHqgEebfXMZ2L3o+AhekoqNXvEqL2ECMHxUuFWL6V2BuhBrR9OAfxp9WSNmy
O1dGXSCncYssyCBae2Kv9v/knpSE1xHZ0gaBFat2Ne/vBcBqoU9mJIuNs4QOptlu3RkwwN4qeJpd
F/OS+a8wVoypeho9j2Wjs/LPcyFOV7YpoJP0TcAAdd8/U0MNSKmisUDX6DTRez/WHJXGwnTapGWp
ZxuxRaEqY07NCShZlRRr1sVW+9cd3UMP/sqrMQegYEiVLNTHBt2Nw0ET3/C4iDuPR0X/PH2RP2Gh
qv+CZKb/obOhLszNS5v+DC4p5ntbQnt3qZKUQQOML1fUc19eyXu3CyMlzFBkrCS2aJOh0Ur3X5dN
KHxEyW5yGqO0zaJxPi1m5sJsFtaAPlQcV5Je+W1ypSdZaCUH8x4lEsmlU/NjN2RkTjsaVD0yyoEm
BpbBE+fhJjecBVzNe5YD6a1TnOpqHWveWvjuQ+bOjCQMHO9cb4Tf4JU1nojt/rhIvgNBUiEgpiuE
m+JFgysiqZwfottr6DYJDO48WmlJh2ueKmvLbysZEd9lNqYRfDQXrZZ4ZwIL6kDHiTKTMDMaFBWs
ujqw2/ZJ8AeOiLjwuRwtWwMFYlvzIMPFnKZbpnQ0BrcqaNOSYmDQ9sSC94dM7h1Mp9q7bny8ZHZ+
VnNb+EU6kQIkJzyuHgmuxNfRqatTQoUME8rt+pny1XIp12eeaiKZtBXrs1r5DjICuwcZa4QC7iZi
G6uqZBo3huQCEc+Iw52o8TARH6s1600WK4WYr2omTjX40iQWCgzY1fpOdp/s7zFTFjlMZyHPDl/v
e4Ut2+F+tS3U677MCXQtxehtiqvheBasqZQNcRUFUuHgPlT2GuxCrooBPWE1u1BqY931MDSbzfsE
bUkA2qgyI+pmAg8TPkr+jBbYI/vY8EK3pCXW7nEzQd7UVXlpnzstlrsT3cdgDoJ/rAc2OP2B9uWA
Hfk2E5U1p2v4qX4KFuUtHQO4RwmOyPUkPst9/riN7oHYf//gze6puqdS8LgYw8WeA+lUjWvj6AGc
79cypuxCzKqvqJ6bHqXfupYUv1XSfoTIgRHUjb5lfHNSnChD5LPZeh90lTgc2CP8SYqwB7Cx6yLx
a2C8VK4HV56ftJwVzluwUPg3DC7kZIqW8uppCLTDvRV+8Lc0HlTsV05H/tLr1lVOv55D5AKt3hwm
GZFA/vwqVx1Si8Kp+cakBJnfRwSDPdurs1Q1DXZk0aAc/pLpwit0j+bkPaKnoL3Abfl8GFs0nCgr
BDjXDAhWDiTPi5MkbjG26KDweLQna0p/QfCmw+cvzkMTPDxpKH7mJ32+yrx7YWqXWFItnDCLixv6
OSUy2J3rVVo0K0HOrDfBhvrUu788dy9CTkLVXGOJ0iXboxrD7SUpVDWhLMN7p+5i0w7a/BlLXHYe
nF/ceK/6nfuzCfXb76xKwGjv15mD/LgkPOwaWzXbplLMTJ5Y+A180kud5g/+6nAFoCHVggVa6XUG
5tnDpRxQATqgJZu0VPcr85b6ukWXp1ejKuzrdh4UVsbvo6wa5L03X39FsyEUe8FetGAjYrjcO581
domXu7U9n0Sl7PggQq8GwoqdJWO5AxWtw4fdV3kEPGD2/LqHhMIgGqMmgeRoJ1ymwQZEMclIZ8qf
Lag9bvxtWO6+eWe1b4zXCumCSEmENjp9hVnSCndkOHGQJu4kn1TRMx2Lor1TRT1XreBut+Uaf6hm
8kLVGNi7bIHNlnEBkrUj9fz01MI/B/ivPywfNBC51YNbufdoEseaVwt9dM1iX40RAXKCfomdjHMr
SFcmpokSKgxDwT5g7vrfeLJwKJwBaEoBpeA5UOQsj3CJlor9CRQKZyEjTm7FJlSI3hw958niuYUy
oPmvHSGkD17X4zrMNL/epkWwFAgIA7b28cuD6yZE/Wh7bYldKP5p8gqwFb4Ls9q4lghU3qKCgOoO
9G43WlgWtkMbGoyHc1kq0ll6JB2OgFrqOYMy2s/s3YtU7mR38lA4WPt7tLTH2KOIdpjYB/PC8GYb
fA1Dx2cEuhcomtzNy7sa3Dj1mp5Z/iCCpO2ot4PXrGUoCrRW144WNeCgnmczhJop2orDzhoi6nB7
KbAg+UMZOpCJw1PyV9nGx+II4w9yc16EPdMMoOlUV/PYj0YO4oMRhxdGL/eeXAYkVxWnkj7bSBDM
AIh1a85JybO+TvSMrLOmw4BA/iQPcl/aAcyMft6bv6Lx38k6QPnJ3uyMNqljWXiUzAQvhvD9DGRz
FE3Rq2Nu05f91OD1TDkR8QL8l8SOzE91qMJT3+31z05OJT3rBZKA3ieyYRcoIvPv/1K2Mff2Q6/9
wUhMG11dL5uTu/C7vuPRfj9F6VrLnHYr090PalNP+5kYZdDaPS0uWQUmqAVhxII4GwzbL7oNkuIQ
Dltl1sqctorDpoLIuUJFRGckE0psp4V25uqYUkw3eDPk0u396exB6yKYioEAwLbqeDs6Aek/zk1P
Ktw8WyrtpirIu/LTzYgmW1/EkuMOsWp7S+I62prVGvgrSNMfYL1W+TagN309HQTmrkENkllzCTOM
JpnksfD/djYeaF6lkqpLCDTAWYK/j0zSzt4r/gppFe/WrZwUf8XAIrB1Sm55AsmD3txTXoRfrlE3
6vbb5eC9WRsQVWZMDmilVFkMAtlyThhnjs4H2WVJbYdrFK3P/aFL1+2H5yo77EUxyQmB7++Sw9Op
lqS2m/W/mvA+9H3OWKcQqgKCFmi90eDVdiz9K99Q68LmeQfu4UCRhWbMt0H+bjTBUWzNBDmdNuEL
5nKtzBugaNapAseubLN4mNG0opfeOIBu2GBfJ+CN87Cg/hNUMlYXVNNuMzPAbqecrtk1XXJ2dc4B
ro9AMi2kwsUpliHR+St+U50bQyRkHA2MAPJ0rDwEor4MHsZp4Jc9mg2Oy1GdtTgcoxV+8EVRwI8X
Dm7m7SUjAr7VnvXbwViG90sqvkinT8kfBD+bpJVWvTx7Rr1qLWrhopNUcBSX0DgAVlkfWvukoiWy
HwuK/3//8rGGslh6q+rkQNCoZ4FJzZAEJ2ouP8KpViOL5GGfeFWKjqTm7tVp771kDJCNlCSy7J8P
KoMB+masyB5jC/llYYtF7hvCiwISUGGA3IOyts/nJCJeo9+GtBvlvrAmi4Sp5OxUsQRuFLVa3Mea
ewrNEq8kscbpZC8JAdL5MrCMrp4xiQtpDruZH1vKnZimzzqlwfrLbd1ngBqvOn594b2sYpTqpVRT
w4A274dbFsG98TIa7B7PUXkvpIjeNx+6wdRCxnMeH58gcSW5f1ZdV7ev+x6OXrcuCF/U0Gd1qkZj
8sKTZ588RzOH3/O//Svtu5AbrVGbsB2xSHQZ7ByLzD5g42lPgs+wTKWfbPNc1ErRo+CGoMnJ8t6t
6h8Hr8OANfW66FraMVTlAk7AvLsy51skb/KwaFd+EyMP0KSYL9ZgPCkK9KctSLI5zcoI9+aRIHHq
b9vvaHORQeHK8pjD1s4MgZ6ahEX4meJTeYw2t0aQjsdvLqPawLCw6DBrRjumH2e1vZA6di7T0rof
258Q95E5e+8w46uHeLM6YXu/wkKQfp9z2KPAMgX8EPA0KxrmTmzjBg/g3aPEhgGJaXCLIzfOSa9n
tNATxbmBHIZg7ZTmpxJPoNLF4ZHPDzA04k1Qcirsyl1WL0OsBvQneZqdOZSGY2SKzBoivICj3y54
MPfItcZGaH6G805UyRgZ3BrqpzER4nAQ14+vTFCKRiaNZqKKhKhith5/JaxnsaILLmINCMXQ97sa
Q+P+MIcU3igCKlp38OO+s7rdg/uKTRXAcuiz4xTKGQ8+29hLQc7L6JgyMVKjYZf199XA7YRT2rlf
sTonXfcY3eDTWLxJC3ykczvdiKMMlSseyz4s5LOr3q3PSs32XQKDLVZoIWCwyot5x+8rTz/yGOvx
/xsItk0o4Fpbn/fBPGdDZxJSAwKUSuxMXLBFpjZyskGZq5heTdzMf1IFnObZ4NaisGftpkFoJIGz
zqaZ5pYSVqlcMBY80g8WsWPKI2clxJ97hZJydwPaTUN/Kz1Ymx/L6feLkT1E6isTudefINhM4yyT
b1Eb6uZKe9z7sqiw0gV7WV9klN8CONMBb4cp+2lyu3roWDkCrtj3y5jDSRtI8eWYA7SST+27eMkT
8pfT4QPTb2vLMXlbFZF6uGSp8gu0pv1FsEK6TDC46Q353AV17O6B0yGHc+nqMvOMaNx/dpYPu5Xm
McUphnaURgFTby+4MNkkxoalPMTdeuVG2nuUllZJTF6VwcGvAMU6DvUUOpJpGZtZz9F8eSpxvzsf
dRBjsr57bGDEjzSawEkHmxtGIn/Pt0S6e0q/pmTTEWATNRq8rzJjmzCHKdjHnpK8tqnTCmN/HO5c
WHslLzwbAuQ8/ceSqvXU3TzKELqrogv8jzFeINrtIYFmgRFrSx0k2qD1uTxU9s38pyWbRdkkK4Ux
d+UgD0DX4MHw0WBx5Iurz/iJujZBcssGmUkpGtBhZiypxI+UNb2lhM9sCySyStzVgN38qVM1QiAR
je8tEHSoPza+PlSEi6lRWFYzylEuGH3LDbGYFJVHiv0jn9HEb3T3/6v7X9XYA3UR8teAHn+4L18m
ZkEkKRzsoxyducSvLX5j90Ih+22QND3PM9H8jdGa9yiklqAif2cb2UqtlQjLyEG2/J7s3wOS5syB
vWxJZlpy33R2zRVppVOgRKMqzIGDSD1otC7IBJ7ThYvsJzm2lySswGF0ydyejXuFdIGdoSFoeUtB
F0Gz5uJ2xPaow3bjJcHq9y6RQ5PETjlGhem5QHhDEf8uvS2sDLxAtll33RkS9B/aWFfE0VBYW7xc
RLqLYD95ONvgvF/m6b72yYAVfx0jOxwOEuucEjoo9Q7BMWir/LKrVrNWTUJLgsccXF/5qghrC7PJ
KULm2uOqWOwVntsLkFb6Wh2TS6T0WBjG5oSsoDouwMBEAZRXc9UeLvKiHN0t9UINOQwkB5p/5ja4
++c1H5Q6WjgAUrS/GZ+SiTZc6scJ/y9mPLY09FuDAsZm1bAIzdvAk1JwvN8VhHUMxSEg/wqPZhmy
A2a5Yn8W+a3Smwk2DijjLVIUwMoqUKFtzNVLI/CrNrZ1iOvLiGfWZvYrghdcaC48vtODceCui40F
FcFnuUhZixMySd8cYVU8VZwzbXbVLxBRs4b/PyHv2qZoi77eJoRYNCzjUFR6LVmULBGGPlNta6cY
igrSuwEGeYqcfUBvevNrGqZB/KCqRqt6M1DiKdUtIlcUp4ugUfdEAr+sOag+yx/fFNjO+yWGQS27
BLrwMmpoNdQDotd/SRq35YxiwRKQBYqy9apGz1mHZWrxAPR5HFlviJUiGjac2wTs3lMBkiuF+Pst
ELIKwrKJfE5Gbgg+48Aq+hTlQ5tJhvS2YZO1QX5UPvAQ03WgwK2EoV8CiUgTsdm3keH7eV+qwijg
drX0oq6IJpadv4huvYzg9XbN3yjefcjjr8eDbJ50M54jmCUuQgii5hzzOuUcSDxmJZpqPrkSiTB3
3XbqvIzVuOaDVGgheA3XZT8W3tTuUydxyHDJKEfJpWGmDt1f8tmxfNnPV4Ww93LRONCqNKiaV+Gi
TKzT1iAfMYIXHsEYkNsFnkaId6ZYCzc+Thu882sldAg+omU4UJ5hfNH23rU9SbfmgvmX38uXZ8Bd
qhpGi8dU3Wnhcx5zJ2rPcjzJP6F/D4mkIRMOmVUFsl8Z8pm2k+XaV5tlnSluP5PhAVt7VWnpFj+D
m0BwNvmvQqN8aBhXMalL2uciRkiM1QqcjLcZg1pLW/LhaqqN+u6D6YPr3XQDj5ii7EFqSlINhkbO
TZ061pUUm8P3cLTI+ncO8dHOQwgkBDk8iLuPOlDiKR5zEKPI4HjBTOkKJqLNHAjERFm9VyPIu/Sf
r3Rzs1pwfL9r7YwdOIarB3iuTV8NtTDGaDkM0gUff7dED68yPXQGACvQ7kNhaSvIFT2w5e9rZSnA
PrTXWfNO8W/FBuDNG/3MHYNOuEurDzpIHckTt9/lC2Y877XIwaCI8PsdppC/CLtwNVYaO4iYW+N7
OItb4vfRWdlH5cbFWYVY/3lHGYekOf1H3Dy7ipk8hyLgkRe2VLXEywQeNpsg8uKwmeSlzx5w4uLy
aIKheUlBnF4WdlXtUBOfhMMdLmyrirTEtZkfBIR5jrdtVd/YY7NzAAUcqO7dEKq4iRPooEGBxPBK
DTFGZOMZxXjRht5OYWL05gUQkWaH6AZMtEEl3ikG0oRW8bocwopD5gxOmVMiu1YJnSmYrrGb00CB
WXBDl/yIgxY79lOznYNixP21L92svhNdb1TyryHJlovDqUjwITLSbL7JF0Dt7lmoblf30qEa32wG
s5171OCWV52QkIUNAJlOMbyGz8YNZuGZrkzTeumj/+iBsu1DlsAToifys8igu4c6OjavfUindfeM
5Oi8A4zCYIgMH47mCCnLH6fAEP/+9nHkRCtRmm2Xq5mMcKe6t0sl6MBSXCkcXA0gEqPavwx/cGRW
+p5rgeXOeXqrgdXDrXzPeSXHbQGnwOBgtKIuY5xADJLeK/Z6Qh8F+V4ncWkZulQF50LSno79aI3J
XDaWdWLRR/zzeRdzxJZsmKjLllnF6TycLg7BzW8GklMF+flofkhxoJR7dDRf81VV3KRfbqc9kf/2
bhRyjeWIvZuNu/Gv7v8TGWf8lHI4Ag7X4cvkWwcIw0ezeJVum9yu17wxCShSzeGVu9C9mi1CuznX
6K2WRzFUmi+gz1HtV+brKijcOpntJClfjBqyNcLojjb/8MDrmY0XlZlqqNH88l/BOoKBKSu+aHEC
AvJucQCpPsyfA3V51IRKER3/iSLX3IzRIyJhFzfcgPzs69I7HltJUyYseCMb25jXD5FK6H8wu+cS
+gAFz9JMjNMkhUdbma5LV8E+1omkpVWiTU+uZcUXd4dP4NzgiKYnQNCBmG+ANRngV6kERI8uih2K
anfTxLC2SHE3BSKRq5HnBfQYszydc7scNJ2tuDHuzAn/Ar3w97kiLqDNE09Y0xpgEsG4slxxugZf
bnhDTmiZnVoeDwS5QJVqHOtdeYZjgf98RchUaQ54M5dHRVs1EoKYYgauD0gDRVajQF4/ADpUiq4p
pYehHHrnsMw+FDLWs7pIytScajsczL2HqY35RNHfguC9ZxG+iTaic8NQkSF8ZyBIKH36oxu8BtN4
sSI0IzOpRe72sm/LDaBp0q2p0Op1Du6bsOLMVetvDAVU5WTC0PEzg3gPDDj02NkiUOmxdiTNmcx6
hPHj3zRl/WKXyfv+16lkfiXH4eUPty+1DQvQQJyENotMecY2aB4cSlXIK/Lz0tFNubBqkUTLdda7
TuOSv6WbPTGkkeQ7YSvRg9JMMECvdzttrNql5iOB7XXImanwavEqX9/dmXEXXA74rZoo4x+8pr4d
Jde1NOTgjg1fCRm5wxqg+rOGQnThM4nAjkw9TXb11zjRgn3sWka29ziBVXlGpPbaoQTx44bftSP9
P52E6G4iUb1dlBXgZ3/H1t0LJeXHV8OH2aGLy4xRNEg8DWLxcDK2HTqJvXp+DfZDJp12xMKTHNeQ
JkiqN1JNLHg4vrk+TYy3YpIpluRuydBLIBoVLoVyRTkrt0jCjXeykIcGwuaM9gw4xWjMDbPxMl2w
DYtK8bibF5FZkAw3jhFOST3SO2o9wpwTIMHnwh+R2Wey+irRKZE3+ozRowCmWMlkvv1QlqYH8kXZ
iegTTm9TJK4KYqyCoqnLEAbZRrpsfpyuqDHu4mxQHYyhXiE8J4Lr6D5gIySpZisMtbC5+Z3hmXSZ
lWGpjJgN3Jfv8TUUCj9VlmfzF+xnuhba448HN7IPki2RNLCO9vMF5fKTUhc+pznUiAckggltFQtL
NtMqjJfer8YsZEOCzQiH53UntveAtPLIbKoGnKt25rOBKo8A76jNaStG/Ey0v/VrfFrj5umwWhDK
i3XassptuQLzp/jtx5q0T8iwPF32YHKbcWAmyRhRNnnDO5vClb9NOR/VqY74U7x+SnZcEa24wMsN
/85BPmL+dWiWaUnAQamREcVPnwc8CTKzdnHlJxAAMdN8L+1BCBt9yAnXP7/u5tNPoFm7Mw+YiF0/
vDmU17K/w3QTk6NUIn9r3mQ6irYRwIOfTxdTuJxCES0AjZqCxx0YPb7HtCt55TNf4dNgwWdSVn6Y
W+gFRCtVcie0ojY1RuEFrBtl04EqhPAA6SVRgV9TQBzFHE9ecFb3uqR+8kv32kF7ELFofudGHo+G
3cj8xLCZUz4Xj5dIssVIPAVbwGumtaFN612zYqCjLjGI7DGa/jozZhz0XAJXZNoYWaXxSQHu1EMn
lBpp5GZkyBfkaWUA1yYSfWL7Z0b1wHAeVi9B+0yqEfhBHCkfzCedSFV9bekQJxefgn8KtuqV4GLJ
4zJJ8S6km+CsPsC69uOHj0VjZEpc0hxQMw2SegPGZOND+ce/E2kiq/2qehTYfpfdRdK6JX1uayXQ
qhlP6c+Nu647erFDNsaumMAu34j+N9YQmS1fS4NQ1sL0Aqo98Ao/5Cwj+49XpScSJu8mWn059PdG
6W1A9GbgceyKaz8awUVCi1XVFPsn1Frbat+M0l7w35P7hJPtefr1VV4CCAnK1KBMCfAGKuD/p1Nz
+JW+49J24sLfl8r+O30xI/fmKPSDoCTtyFPIYKOogXXiiqLiGYdlF4HYtwCBoAzXq+6qR4x83ktY
OU5UYb8WgnZBlx/UuwIrSpvLHeqLtseuBGak5xGjliDP3k42Smy6bZ/m7LQ1utlCtfW8fV9wj2Rx
WmLMnP3C5RNHubtst7AArrPHVRHdKSeobvm9HCPkHKBlZAWc3Cm8djXXxCdzpNSHjsc/540+DMLp
sQA7tYPSB/wbZvFZ1edGm49iOlyfGieo8bM3piYjBUg2luZgGSzZ1yH00w0DvKiHCS9rLrs58pfn
z0fjLtNyojOfk3HI27OjeUvZDX3sgomAAAg1zrxdzxx8mjj/wMvccV0QMUPAxjm+kHD0oVZuP9wh
Hj5dr+nB4aRiLt2P9oHpDjMIGmRKB2VeOSGIf3pgh5OshgkYYio8WdJ731ZyZ16WEfZZEMEIgdU0
wouBaXaKiPvCqGBGj8QcSY8upWPci2zMqKKDY4ntDH8WsSca7OcZE1OCvYRNSk73oe6eV0sZODdV
cQPsewyYFqRWKRpWVutNdC9HPd+ezU7DZJlErByqsqEIgUqJfdGrasqH8UyPvQzkhI23L/nA/KdD
wJPMtu4KUu03Q7STnHrnLm8N5zn9Nmf2fUCZN5jgyKoueQuHB+unX6Kp5tiavGpqA4oZC+gDG76k
EkT7sRVMwKbBe9LvqdrIUKqTX11TGKnxEOCQM+JsTTXl0H7tdmhlhOd/Q8NnwlkHXJjVfnegv5Qe
UfhFsRH7DPd8YU559Q4pmw4CcDS0Wkv9tJQx5W63r/hcARtUdffqkwYCpjVIij335Md2rnvMgJH9
P/D9u2aFmjJ88UnAOX1iYIIIiZTvxwGMMwuYHWFno010wwslzpRacAk+i2NtcvLRgxs1VuVqFDXr
f1PLVZVgi/S4ZOOV7fjwHDuRXdS2xbhKm8MzWUbDgIea3aPcOQbhVT+Ue17thhTRJHU/XqXdZIAQ
4KxjsDdnQ/OkQRLsR/OkbCl9Radqy5XCJ20sDG8dhCCMqwrKUCkVmA3eyIVTNm8l9g2hrBlHfMA8
ndgD65AzuZB/Jb91fMDL0u49K9C8wWKIqPA/2W1rnf4dja10XYYoJ+VoNyWiq+aGy/ECCXqnVFyB
ESG5/nTh9HdSpqT+0pBS6ysn5Z0nPCUEQDMI4Y/3HGlAh/csJWg6nhfgLsjc6xY+30n/TB0oghVR
KN2ofynXQDhWK1qJTnV0zLnkLYCdyPablX9t12d6HF+NKCEGpkoA/kooD2+aP/kglNdk63Q6DcNZ
KMNUJp/yYTdjPnNU87sNHmasv7JYZEhFXjfC5TdbP8Rw0aBF6PQ3b8BcdwV7Oz2u4Nowwo/fHMTk
A4VfYMhzfC+mwZOr/Rg7zYQCwVj1GSazfnFqJrP/CWprbvH7E+xnk2tE69cPzTnQrkLqKsRzd0sf
q1sqnmqU/eS8skvnF3CFIu6jNpzaLtXMxjiLpGLE5PWK5TALYMhXd8P9wb5f9kDiUrypYJTA2eK8
Fgd9qy55y3aCBE2YVhiLiBGleIKd97OYUvpQDSfmVlz1N/TEXCDsm0y6AqPL1GITxm1VvPbSDfEZ
V40hhW+6JdWf4jlqxWJaGa+TtVdUFNGW56HouKh3+kYsysqryd8BW48T5KT9TcPpB3vt7JCN4mGu
4UFcPSTgE1ff5wvRmDsHYQg8RpLC06pMnQkwGzYqE8cdVLHjTOkJ8rFYzz3+2k/T20ewuLa/bx9e
6maM6ryhU8Wkx8YD0tgV9QQopzl6uyyExWGmAnx6KQrp2ailkzt2SstKr+ccqe9+x21JqJPI5s7b
HruhyASQxpl4umD7N2SwPTCElt4IZp9kD0cHfxWNrjkBrREtLbCLjeNZAvO/T4sux2zKFxu7bnHP
9qUmsX0kUu0+2XICdChm2nUndc84wrKvU8+/KKPbYMsZKk7x+SxO0QFlt7ieXEZc1NiBb6O/wy1z
1fuFEkAb3UWzj41nER6JyRIgZ8AgLPHvsv59jo4MNeeGjuc4JQDABmPplJMnySFau5WjEB4sgyfH
qTiSH598neLF/k8f/gKRhRuskFaMxG8K2+blYctxxQ+OPYbssvuCgbkmYRYOpBb10vefp0s7S/rI
0aGXbt2bb0rhI9v/8zUCH1MFC8Y4IOTmhvDwOyyiqxkCwcb02Zg1ZkVLluUG9f5AuaEuZ2MXmqdA
ElezKsPrl/ZPJKyn8q13rh2irKvw7K5IVZMqV/uzpkfzLW57FpsxC8tKjJNxYptBr4Ubb6vQ4kri
7fhNakkTzRYpvBA/rxbuudBTLjN918HN3pGmwt/S122t2+LipJY21XEn6fZOxifdaycIcmlCnPnz
JakSMhhnUdrec/imAaoRH4E6c9zGz/Ccpz1uucXscHyqNDiYcRo86RwIlaBDqfo6UJyoN2NkQ0M4
gW4q3EMgYOlTqSTUKVPnZUjmeqBXgp+ggI/xPzaR9OivzP5fNbWTy4QG7tbo7vivqasHsDCoPwY/
wsgQgd9O9YgBaCv2vLaA7en+jcsJ8pVYs5g4HsrJs0YHnohPVFRh+QSZ/muSsxOlIhC9qVnW+EKi
XYb8BzP6tEDRl42hYnLvPEynip5erZ7V6dGZBVKPd5daNbz12ES8wHrErkyCsHKJ2j2tMHmX1LK3
+Hpcy0WqGHvocai+zfWc2ajHenHd2hIXkx7wuToD2IBo7hoxC0Xfj+y6tuCC2Lddy0YRNMCXQ9dp
f1KlhTbrpYqJcMzhoBYz9S0RF0o6UPJT0rOQZLl5MUR9V9bjC1Hn6xQNEd1Y3U0lNWOm18SardKa
S8VlovLtfwdpvbaEmUUIi2xllc/rmrv7pWePMwzhnrMTyxYgDMO3vHsDH3oS/rVpZ6PcXaYTmx6z
ILQOqzNemwLZjd9B6dO3T8JOvFK3663UbA3VdNrGRe6DwyBRJ5LecjlJyPqjOer6x+euhhG/dF/V
OdrKTntVF+uqob3GwLUBA+5vhmv8nHliOfE0jU+lcsjCeoQOVayhpoiLgNDO189HTURuN7v+6A9L
1CTwaOpBaYvQDY0+y4SyOQOfESQLM28+7s5WiCJx0pAfN+h/Nq+grGH/rcCx4JZfQUsmt3vxdk+e
tiKp/Gf66dZ1m/tYzzKso+oN7iSN7KhseUOt0qS4Z5EHgSHbpe7srNwHHgHPs7h0OuwSTvJ3disX
UskERl8MSOtu2bw2zVwiU7VQavESXoK4WTdFC+gEMkZnL2DCgREQK0F5r783FM0q8R3vH3v6cv1e
xvVmuUTi8PG7TZdfmDG7Y7XLIF+B0Bh/jX7wOXl3drZmGzC59seqE88yPfRzUD1keL/w9m0on+34
kmbwIGE6nr2m8BXoFUJeR+QLIw3Su/gNc67YgA0f8f2b/TLjh+a1FpPMyOHqUfKWDCaY3yHpiZbD
SdhkjfkiFyRwWL/DLAUytgDzEdeIimKWYIhrk0VZ0OxydK6u+KyJ77+R+FUeFGhZLcqsBoDDZBvm
qhFhb1vRneHuRwcC8ySx/8Q5yWU2vzXJYlID7tK3HB4vCl+ze9OxxbF2cS5E4FCX3YAewHmZnO6T
rvMbNonNRG5Ot/tt2nJP3i7eK8svyjUBI/D7AIe4p2ztTQ49r+V3sOcvXTlG9j0k6i690nLozanI
42KGkUYQkwvmlE4x6dx5N/i6NRimyyAJD4fZFCRpQkCmJQQ41RtlQWah/BTgmrxaRqnDiCCs1fzM
6G2v98262zW3E5en8WOAmOGcwVry+zeMiQre4a+IQcZveevvl5XQGVD6TpD6SPttX1YD2r0LBVTw
MqtqStboMOirw7xt5c43sUOuNk6EJvwJqzMwpQGGK8bR7WsBRSG/j+kBajrKOW4rttwstYo1Lo3S
Nri8pt9vTTFA3wDttpTIjS/BK9cqQsLxmmixyZ5bPMZHdhr0u8ckUckZl90YRIzZiz0cgdAHx13Q
Q5IsnbpQEkIMlGOsaaaQXvklVKoCdIV2seVffV6pQJtX1fQlGVS8ieSDGtPIc4/5FINqy0+r+EoK
mdiMpB8qfK/wAkvlEuoPyYrW3v4ytgtEy5LkskhDZ8jZGo9hofVPAVM50E9F20wHwQiV46rRWnxV
17L6zUmEEkRpgCpiCbPBcCAmACWLLaSwYKFz/REMs8ls4bvQ0ILbe96mfDogW+t4e+16Fss/cXod
eWQ4Fe3Fgq2/5a5GcTn/5lh9hni5z2UmffTSbqy7066+JWedOkEyJ0X+lntk5ZW0Guo3xo0j5IuE
gXkjqCBPVEPTMz3AGhkHOEke3jiCxAgCyS4GQdU0mg2EKU64fOhN4aLKF2IoYPE8Sa9NYnMS9+8Q
igHxnpU9mw9E7nHoqR1KnCIazvA8MjnDAXAHc9oYRt+bWz51GnU41RFIGCVB2s0Z4hW+tLWX1GN7
evOR0UqitwtxqTRqY2u4TM87x3wyAhHjthetOB+41KhCkSJZ1/n26iXTczwbvOYDK7Zx4yAQYqMV
/xYBZforLbjxnBCd+ccDpDWOMS9T3Dpf4kLpgYPEs/ObZsXeOb3A6enXIn1MLjh2iZbR9AMmIEYL
w2qSPQuxI8/V2yZdjE1voGn1AYPbWD3llBcNHtzU2FPt7Q/3HtrE6GRFpj270USDJ55Hj31oatHT
2ngQBzLWMP0Q/AjZd5i1HeXEdEr/OXYkeja9gQpWkuF1FWbMiWZV0JqVhbJ2EoF6cMQtf+4esK1J
OimW3eu8Yho0m02aP19D0BAPnBZwFtczEdvavDuswWYqMlLhN4Z2oRooJj0vTMGWDJQUyvCZhz1w
B/WK/jCGWjUYXlMq7/GOSBXkGlLSMDt/zZJmyzFeTk2Md9UR4nC1BxSoLGmKDaGcLS7XbUQ4pbvO
+r1qclGoGw5fNRtVFVVBw1Owfd0yBRSljn2nkRsSMN9dSyAwgksu6hXFFMteKCXqwYp99mvx0B5X
iViPNVTsDIShAqsNs23626skK2+E2Ksi8rVoDugbtl5DwrgDrmA17k497kfssCRiqGoZzNwa253Q
0Z+XySdRAKwGcsVOp0e0IV42zyJotFBUfMCv0zJBkaLwMN552eUVI/r/mI2EHfcuCohSkbvYv6Le
QxqI6XC50F/qrKyy78AOOHwbBovdyMrZEo1dKSCs7zwFRQVxawhLboo8+eua2hJbQVRYdIpNQev/
V8tJqCn+qYKb/nKNmZX1bZ0SUFgiMdznk1jU1LPAo7Gzs5yAhzdQa2fQdnRzJRJiQFaRq0IoZiqY
t7Pa2sJ/JHFP7yNt/7jYw0itsCtmIqbkPvAItt2BGIpHnCfyGHSNpCRVvDNMGCTwysHCTf4FeKTK
FooKqmfpFYfoBmF0Atx/sWPJ+3Dd/aiz2//ByeJzrmJ4rI10/eoyubcDtlbTWazIrYgfQHbDEIVc
jTW9RkshMHydeR0n+hCPupmRjbJyCgoVjBp22+TxoDUR9KLRW12ZeJ98W21nvt/ltsS80K37aB/k
m+cmJ5YRNNLtpY35zfxFJn5XaJrH+jKw7ohTJEg/RAY6XyjK7MXIF20rmI55HeshznuzvEK7iBQ1
+u5yQj751KFuFvcA++MDsvLOvqYT+DdJTGYHk5wHw1dWbKLYYk4u0lDYqhH4hPCoog8QCiN8BjkY
g2GwtDUgThtZVXdYYVmHICTHATVGhzRzzExuqwTy+jR3ZHf9MhjOtK5JqP8+EjGJgzLpejZDztfo
F33ajluCAl0mxenErQpg3pQ1AzzR/lim5gelRmPxrTq69LkH4OCMqfYje8TAnD2E4DiZ1PpjYKRG
HC10larkxGflv6iIDV9cXnLC7BYXjIkbXjYDDeEPH1zjCtZTUWpqmnVEJC641Um44weuCPQ50gXi
d6mSlLGKjZ6OER1q/GWa9vBpFlFAqoq+LQEGaLYHvd3v12mPip4Lxdl8mnwZGVeyWQSjIsZFQI7f
17ToipVe/51CT8APo56O0KdeqqFZd2H/n4+oTr35HqaB2yQPimuP17o+WRgik5fo6PayRTpuW9vL
CsQsK2aEhSz0q41Ji3eISDISofdCyE05/I4+BJ4RMGdNl65UGLQZbemmMCUkVyalh31aNrbEn35f
wtT/Tpk71GH+OsRfSrvL4x559qqxAXT7rpZaPhECTPCZS5blY18k8I0/zZ24P16ysGwCTwcfVuEx
/fDpHMVhvMCyC2cl/BuSKxfgo1WoH4uzaSuXONcfXvbe4ULdN9eGg4oBy5R0guaQQSVWSPBnPaSc
3vvzW1Y0JmOzYaWcQgVCgURBDcl63gEsHFgVDXtwOwV56ZS2c7JqVNCRtaGXNjq7LTjOVbg9sddu
OZyR0AnU3iURXcJgk3TRFY/Q0Vb7h4ykj5dX231mM6WdXKpb5aGPz4KtQ3tZm0InQWTdumR1PxOF
t7TicQnDi6PHmSVqy2G2XvSEc63M11cLUg35hVpmE0n/Rnlv0v3ZBEBbM15CyuaQV5J4s3VyR0qn
kBLD3R7YQQkfjRArqWKZcMScugUJVS93pM8AwzMM/RjJevfcfS8DTYeuLeDr5STvhIRKkEmfLkkm
TWCn5DhXDyvm+ETTAEkFBocKQ/7JA0WhyhVr2/Czo0hXQQjWIf/haE2JZy7pcWUtGkcHb5X5+3Mt
Bl5ZdQ3UiIaa1LdG0OrN8kILzlk1yRcYLkRQI3cDiVXIF+WaNzQoKud0zk4yyyA8yqubD4mnTrzG
0auCO1hu2WOueaUUlgeKdOV80Is6htwCKYiNrv7b8GmCDp6v1TRd+WdAZm2wYK5VOApHJ6hdSaYQ
bgMT9+0p8hW8l5QYCingN2aszAEgQS3EO5+1lufS9E1Vova7/8BhZfPmde3RBv7RAYtXnKk/yzqt
FP/9W/0ULZSqd07Wiqe3ZS5lrL6TB9ErHIwTiGhxJcI3PnnufwvJHDjdRfUbsmfgOhP42nRsF4ih
5YpI/W4cikmT1I+Se+5ncJh71qoDp3toP4Qd8Is7iDfVG31OnjlFhuxKQ+JDDGkxXhhMY4C5AcO/
wPAzD2tnqT5hhK35vbTIGOf50pULpIBv85bDvrvxcnD+lVWKKqXNCuoZChZ9GPcNxCqAeQ5tWtqI
BrYAIkoTs38HBIO1zTHRBoihgHDXWJFTlEuNgeV06l5gjImF3oVNZe2q7ogqjkHprxigPNzbiZiL
iKBa123OqVZ1WzgHqkmchZJCIva2fuW4CtXUvcsxqVBbC2aq6zVWDsMnfBJNKUpZD0Q03SkUkUJ7
ubBwjYugYgX5Vrk0F/RveP5ViiAlqP8GSmEBuD8mima3C5ffqPh7LYRPGYfPoVi/bbc/DdQFCcnH
umWZtZqjeufC7li4IJMkIrcEsbYEK+QtgyhnHGXvCdyBCgf/ABQ+mGPHGOpup+dhUpDA/yxAvpLt
xETMMS/3OgF8J/DvnLahpjQLHsMKVkr7BtdRYIXo+vz9itNRYhW0hQLj/ogQUM2FWfx1zamseA/K
vfNC2QhTJs7xjhc7YfNze8TgazA8aok8wEdIA8lJazJsCpJd4Qb8EYSy0zteJjqQUN4EG1b4FxwT
ArOWUboNkziGq4KUbXdN4gt+kqKCwLU7nvUxVGwBuw/0Cjfp/aB5CQ1EUC89oYd9NxWzYa+ZyF7f
KZBqLPPYyIia8lxYNrimdJBnNIWiWqvP3GnXuZ21H1o/NQRbByYpfK96Kw+A9XNQhcGBtFq0BYN4
o0mrmP/jEHv8+iuRrz74gQSIXwP4Qu2snG+bBscuWjVyYJfDYHaUzi9c0m+g5+A2VgB4a4eBSp3l
7hwBUO3/lUZHkbGSiwoTpdkGGd4BFEiSPRrxIl72H+x8oHj0WlNo7o0Fq9DcHML3qooKaM/2zsUK
A6cKqiDolnxRUWuClbhfzD9Sp4ig3JOcvA69/0OBFhukkV2jkkbbITBTTDN1At5kIgzZmQX5rmWt
yrmcQ6pJepEhyEM1ZpPoyN63aeH5hiFXCT7ARK0aBFWMp9Gp9/ApEbIee13xDMgNnKby1EJ1Ycnb
szicd1nXMgQe+oLJEGDamCb9A8UHyj+KdthX+rxgBz1ODHT8eDO+90S9ErFJIJKYmpuLEpuUJa1r
+MW173VDmHNjdwLp3sIHVj0iQ2VLmILjnD0waOtLt2QF+X/ascIA0cndH753YirTEWKl8ZXXz/Vp
212qhdP2dtLgsKD5B1dGAnAfLPH4LfdhsL5URLvI6xqd1ZS8uzFLC4vZsnOF5SSKfDuXI2MFrYI8
hSg+GyhdE+jiP4Mz9l1JezMVlEtRMld6Hq3Am4xSJe5iZhcBxkksCwGyg7T1UomFo6+6HRm9Q+Bj
1LGZPGn6JynEm6dFfCBCHHjQkhjtmjy/9sFu7k/xTKnYpezqNz80fswgdjVS66KKQcoE37Cdwrf1
4qShOcJPlBbxRCelHQftJZIfcK01x0rSXZ/1hM6SQLrlD+46BPO4ZG0xqKHYU5kYMau7JouvsgA3
b2UbLca3IipwYbU97OUS7D1TeSC4bhPldcEB+XI9TZnj49HmRemXSVRc8yhMGQdJN2rpiUH1+O2y
UNcsCC6ExfiK4smAGVntdPeVaCT2bsAgjuoBpZ152CxytkRtIFFR3pvLo74zpw0R3sHFkvuyzA0U
Y6GZmFaejyh960lxWaIBdIy1oFtq1IaxYv1qQN/5UOg8Urmt1Bqkod8DQaLmG3NfpCnJelBDmTpN
ALAn82W0QFz1f2t6L5ffED39bOKwu4uAVbvclLacwKCqU7xsh2vfaQySx4hR8jSx+y3YoEN+9zyN
bxMUfN28mqu/rpAT+V3yVn0h/+jkUG3C2owHVOYf8IB3ErCEIqv8QnQJ0YOhTlSHW0wPuIuVJCka
Mt9CiNRqa9m3s+Yw88Wz/bJgzRG4N+CvUsKH2a4RBstkhN+iTUdUDl6SypHlvgR2w5d3+jNtYLw9
Lxi0hQFWGQGoW/26NBAT3uUmNi5V8k4Nu5P3TAu7pWzO59mEFS3RWyhMlOGwb0/4CzVP6pkL7JdU
C5Kdxlk/njLMnEhT03ugvpO/fBBEj8FPGSxIw6/EsvjazqYUMpoTJrXfGFycvFLhZIFrklbrZDBA
gx80x1KkO/zGP0gRi4umUhNOn2dFD2JpbDN+t11W5d8UeV4Wt9JYEwKZydAxVgSyV3HedhUmwkQk
CqpxeQ4SqirGI75HHoDQ/PKWJV4aca6vdAYTqo641qkgAIhytOPbIqQ5VR740RzjoMnPxmM5jSRk
GqweeWmJSF2useXw84+9e4sOE4k6H9ZicjEKSyTwnDwRl7KDySHO5xb1mbwnkWyqqsqtaLGtMwx/
xNXfs9qyAPGmZiQNTgNE6xhS2v8nwaVl3u4b5GOoNwYMifReIr2+M8Oc8b9nOKMqi1nP82aIitLR
/rPaGEYL5hkKeBOIqERA6Tbl9Xw8nNIu4puyIkdDZosKYTkuNqgfd/MQKyfPNrGUdtK3vcU9rcvx
tR+BQemyHwkqSf7kR7EmigSStgL/qaGgBafe0fkCvxqkcg5UNzBJqEcMhlG2tWx0mIGuJM5NV8cB
2zFBkQXDszMl+1nM01Yq0Wzgv76Hko6v68OWYa1pwB+kV9NM4HKXOkQAuO9386Eg49dog96u9GC8
6XBtkpMna4G/hkJ63qV6izNIpTHXa+rN3jeLlpO6ZzZxud12sSavxBi0lhQT0aYS/Gccbgo9szSg
KOEEMse5IZSRUuaTI2GHRwnIbbdAXm4EuvwzuVoWOE6C3XCVHosUIm71BfqSuWUtvLkOjGB98mIC
ss/AeeMIE+WuvFPAwLTpB/j12V/JMqKnVQ74avQ+qKi3eN72kCy54AFOeiabD+nJv846vWdn8AiJ
qQM5RidgLa0pSdHvt9gbeta8bIuyqMeyjdHEiDvJvD4jv9VJDB2EARPuwu4yKjRZsR7cubLIzaAr
GYuCEHAezJE8Q530F7hlvcPrKCsde6NJWFuIowEuA5VGSTTcX2xCBiLTMmvAT1hTLQqueL8yn06n
l28fEh/iS/yAJuT9g7+MeeV5XYqUmO0a58nHGDpToU1fty7WCVGKvfiyT4os7HVyQ8wn0EHzi29o
mE98igy8rVijUiABd26T3zFSnf8NmajAaV9Wr32gHskU4+Ax5s35MyguPSAI47dxFlZc9BfbJSAX
jBjYSS6ZdU7s06XyT58oTOc9nc39mHmn09pUP83FesjydEjz5e9AEpNMzA93p7e3K9uj+fODlpnq
skVd5tC04QIUGGOeuJBB9dLJUfxLe3FUZaL8d5Y06hiCN9qJFU6C2mC5UVmAbiqV8KcWu14OHK9K
3kAXDF8BW43XtnjN+f8VTIIsnCv2czjMZaVJPNUT/6GPHYuiXaW3rLmROoKr1X8f8+Ne/mm/cI5T
ZZbviPVROcoYF4dFbnjiLF+B1+AxiXZ90JgwTGWutNQRj52S7u61YRV/MH6lDodlyYhKT2/hcklo
FLwolKz9Xf40k474eA+cDR+7QdggXLweEenYvLdjCJRW41c1Js+2Eewnoue4hkCbD9Y6ssdqVTZb
EHr0D4rePw59/dCjEKI2qY1m3QtPYXkUK+X146VzoB2QXmP4sqQJGKUy8pjzClGUqm8oEbxW4cJk
x6Vidl1SScBynIl2i1z6PU43WXkbBs63KJR21BbxxmkSzpRvzJGx8qIlc2Yj9vrog2yKzFMzMtDB
OmjG6ju3sIXbXv7rgprGAwp1mrQEQnoofCZXdvbtPd/gMz591STOkPSTlfXdH0tZWeGcrsaLIR/m
E2y1MTlbjdQQE/BOzZ3frokArYmDqHtCtnIMArsjuCnDXoZh3MiDMJqOdc6isl1oEmLcwDXL+O13
PozGJgrc8sTdYiKK/ERArr3e3kkWPXasfz9c6AKFtJ6yOY+g3Gp0biX6T97XoX/l9bk4ZUcrHAUg
6185wLdpmY4CR8/55Kbl3uLkwITUhxuu3Na59jDgIu0hfMFFeQPHACjSeLVR8+NdCBnO+4CkkxR1
dRvct2oJlzCuoDdVvqSDeP2q6ph/LvLMXpJGTCcUo/TvLglV/5HqZIJ8GiWdYOjJ1Skqz5ftNcsn
a237QKj0DDQyYfOUHvhikz5enczjoHO6HVlGIQTIPZv+3iCYBzVO6vqAYAdpGMomWpZyZYZLKs2i
dI3SF9uESaJIBDv+r/092FuYNM2NV0gR9HeaCXGbb8DXcZpfPl+OIALduaVftFgWL8rL2Zwhefpy
5ZddqA+uAsiHuGHSn1LS6KVL9NaM1AgCTpQs9ZS5zJxrCSxx2UKRJ1NEzlSVTie2wiJHr/4W2iq0
CLjQGBmVDIyk9a9gCbXLMVirAUR1w1J21OEiLdxXHQF6Q4/gdqpVM3yjTtyiauum/9aPmCxbT+w2
ETlTKhDivb4h/NIjvw22XpYrRxIgkmMRSicSBJhudTwZVp09pMQlmJ1khdtHGnZxkFWrUba9A2IG
/8JGvHiwv5ixbX3mYFMwO4nRluWgpoWjqM1M/hLbxNrKZnjPlXCZNKsq1m/mD6pNeHe+eWPJ7ONJ
JmL4iMefwEXr0bI6wJbQc43Z1YUGv66WtiGpQGsKro3EGFqXzCJnqnz9gOUUI6eZ4wQp1Ff9Vz1c
TAFNTt25vZtoFGW1WI/xQrTDCTmp9lyWnm2B25a2rJU/EH7GZM4khj8GnmITmI69My8B99HUD3Nq
sn6bRHGlIZmmrkfA3F9kb+JIMZz7xjoFvgDEBeeSUno83U3E02FHdgxgiLVnKEeiBaOLmmDqPxc+
NBrCohwCN/VSByMfPgBgsrjQ5VZttf25KSIL9n3P4wSiVcrxshoHtsIz9l7MQjnytJ9Daa1/IZt7
TySkZtAh43xj+YWkRCSb7LUZJAWNz3orFT+INlYcUh1yJ3sD1SRonsG1XCw6j2mmGD7ww2IwdrL8
n3NSzIun8sjiqjyaJzIlfjDjnrTDV3vxQy4LCNvRRznXuMr7yl59+VhyF2s6IRWonqz0P9F3lliv
avgoupLP9eJV5Jhm5uZaY06zVrn+sO3pEoTDtxkXbywHAK7y2l5ck+Klw/tnn9bmFap6U0vUo+Oz
B/P/Ne1zrn0zSO+gkWPB9n+m/fGf+klOHmQEdbgdiUCqFiLMV4PFEcD/Z2ohnE4jnyOCjn6ugNCj
GszS69kZmsywRmBsubVBYzspRfZljXuStZrfEjyP/FJzBBsH7qOih6yOAlxYDvqyiqQJIJe+u3Q+
11K7OUMbnC7FpXPHINrbEDEFxMXMoldXXXJHBykCui7qFYAet6Cr/eVvXDp2lPoV6iSMYjUcc7Km
ezMOPDEF6cNOJ1kAlzK+Ci0W9+nXuS014aNOX140rWHOl8xzm7TMxnZPXxrtXu0NcCF2tviU8maH
2fSlJSr7Wa2PaLZPSXhr+Q2dQBwe3SbmWomZS9C05uRWsL8NYxtmnUTTzYcQZwFMCSn74dDNqSEz
hOQY8PYQ2lKBQZZsifHoTLGA/JxHitjJI8m0UkSs3H9D6tsBgteKfRpyf1KJq1dcmOlyejBLrRb1
zn7cpfTbrBeVAlqXb4X8WSzcXN0boZHSuHd2nswuHgcyguukK7tqr91I6qXHJO1h1k4OVjvobKrl
pwzjTZYovceUiPAEFRIMysNBkAO2hW80+2YKRkWzGatDF1NB/rePSecYKfw+kWREcb9aH+jilSsj
lwRN84zV1PKusQ8oigm4/Zxhsp1tPYZaMZahO5yvAvnP0a9/vdbTVi+GvZEf9WbtQOWEYXv9B1xe
pxCitKLlDek3Iwi4qIxZSnhKelXTcjT6j/oVlOPkql57xP7NHvmgDcqngVaIMiaAWQOsrWskHGsa
2S2MppjAFN0K94nfH3hrWT+gdK4tmUzbOMu5FufiS1GrJmehAXJsiNMoIy8/wROvEgkmXFXHAX+1
Z9wT2neTdhR/QE/5SAzg3Cp6Qvlv7oqfyl9qxx//vXps+Ih7n7vQLB9AYWN3WXFsA6sMwOqxWqiu
sfXTv+IDcj5IW/N4/tHX6eQl/xTW0VeNcH6UH+qiM0E+OS4hpxN3I4HBTg9VPU0xqqxWxULJ7o5a
0sZVtWIgO/sSSv4NGcZThtR92CLlSMUz0vGPe/CDpH1Tkop9HfyXNkVjrk+CqezAVmOGQuDcCn+J
y6Bb/HhAAD5od8FTI4CAaozEkLChR5qfZE/6VkcpDT54U0mTqHgqqY+ICgCG40jgQtgvvuQoHVcd
LVQ0KTMXv2iPGkRUgVuPBeDv6c3KN6KRG1nH0RsMDruq6VREYssSuSARWMorGnUOJkAOkFHTWuIX
8ACqVZQhQn2obraNnbin7PwYh52AnH0iqlwqwSc2c50UCnRxkOFAKIvCpgzKF+LbYusZZg3tc7nO
gubEpwD+6mGggzBjiqzDEAPhvriGUMMheVBdIUYdAd7zM9UAcy9zyfzQM5DqDn6S7sKkkWzKycdT
Hb6ynSESnpff2LfmgrFylBuNUx06tdtWDY5t7kbYGYntSo1TvmUddD+9X4V2W/AW+Zr9Ekc3LPrb
BKe7YEJ1Szp9SPuX5VLshnwk3XUL/V3gQ5/WG+vqjC6wNMK3VExMuw2TDb+ZKZ0PDf3Lc6bttET3
lmawkXG2Y8nfSkUb4T2c6spYiPNmmt0Zww5VGOWJZ1FB0UClb2N24Nxf/3IljcSobnhK2zXiTZ+Q
aUh8yNmpXWC+XyIfzTGvn5QAp/OQew2y+8T//hDZpPvD3HeUKhOnTPBFRxxf/PfUW7VQ3f6JBbuz
Yjg8cAHwAL6yWQEK4LWgG36zkUkqLfBlnHfFvjqBdShHZ0bcTAkCrvGH8btq1k7ZK9jiDoiqpht9
XgswIG7DZVgP/4nGLb7fXrywNaRrtBRPNbMUSowke50KiwD6MNHjd8WQ6wq5zyQqLNa0zv1TIJ8D
korbpFJU7IiDN/riujW08Newdb20Hsoy0httngqEW0FQ93NBe/IQw3V5IVLcilOlYwSYXDWtku9R
uFmJDDePDYvvO/p5QkoTeoswRliGeSQfi5MhDYIevEbPrwwq8TCDMFrzVawqrduffOVkqhbF0ICV
OpFC/j3JydEBCcofyXxa2cyQ3Nzmpg3Fci6CG8+k6FyFzv9AtIOzorgx/Sm1uHHY2H0CrtlqsSpm
5mg+XjStJnOCzBVJXbyUCcvEE0CmKoLjk1nSbujeOr3wWfUpgr8122A0EEeNM1rc9Ns0DOJ7ZgGh
DNA+eEACdELOQ76JNYsAJ5UgG+c5OgvfX5W2wYvM2GQZ2l4U7VHGAtM9w9/RRwde+XFsRzfwbTC1
ug3RvcCnQAl8drOscVt6+MPQBaQGGI+54sAWmEDer2mkTF76qWgcVvBjkl/FeadBUb+S/vnOZCi3
u5bBQq+qfcyjO15/7ZgHnh12pNhFKtX7EMogCo2ChYcjQvr0Spdb4olj3UznnudVZnPk6lWnu/f6
c7prXjT+lDw9AYb5ZJgdhJnLnOlEr4pI5XKPM0lJyZccKMNf9c9gmUvqym4mxqw8l5AqWHEMfuI4
TAZeDtzGQvZBXIEoLcqlJXK/+94GDiF3mNVS0RoBkOuKcZnV9MtDJ7oyaxxrTqz0wqeoPhM2WuWf
po+ny28O6Gj3/FYQ57aobloe1ql9n9W6yjxFU9vSqe5Fk0vPDnUsLFhlTsGsdPW99sGS2vL7tV1M
EArexqZvbKtIbQ8XSvRRScqciY8MTH/grFGAXGwNZi9J5BsuHMcDQH0yLvI2dkibIMAD80l98AYI
63GIyTYWN01IT8uXA5wWM4XP8YM12pNOzJ3mPC9WTBBWQVk+CfPDgrhQ0vVVufLapPdzULonMaRb
ylBKbex1BkeilXtcP6Fyz0mkVo/gVb9qigkEkFeq7exgdH+GeKNhodKcFtVwKy6UyTlyvh9a7ngG
95KT27CAyVVBItUh2k5UATSjOBOjXORC06REGlr04bnr9S41bHc2wMFBj9L8nJfsUEu9uRjAyCr7
eDo+jFKdvZhFteJnLcfe1+0l5GpwiJI2Vy/TsO/QkWHMdF1BVwQucvbPTZIx85p6dESJ79FyW8C9
FR6ypFhuCp3drABbm8++YAh3Hq/LGNcMoZRFvOB3+g4J7kA762hFyZEjbXvwy4ZScnAFxvdSfC5Z
erK3te8CF36l7nUSYo6c/yovrhbvt5s0qorsImGnqhp57fdXr81rFqz12BqciFkWVx/D7CDC1ZQN
0Nf5I5WfWe2oxtDu7dG5nc1/RQJvXfRSVUMRTGmnu8T8tzZ2hOK0PjGknsOrMfWGshQOXEVlK9Lr
V3CpS8trx6KplUeHkNjQPWgkoU3No+039uXo8jhbD6Ezs5Vz94GtzcpDbvsd2JajEC/J2E/VU9Ju
ehLb1unOTwonCnj3+pGOfYgSn4aTdS4PDr/ZRDvFR5vUb+8pJEz2CXwVIJdLKEUSRL7NvmPoBL9M
bQyWIvWc38KTX0pob4v2d8Y8L3FnEm6r7uWOOqw0Fr2P32/vkhMW6k4fLQkfjcIRdXKewKVKIL5B
RjHEFWH3Ob2UXfVHWsjGXCUe6rGg07xK4XyDlKjVxPFUy20PcSOfzrYgOlI5vMvamggEDhfvbV9F
3L9SI2WB/A1ImhYw4j1Aa/Z0SfRxEs03umLJhnqWqSC/jQcZJCau9f4m3XpF1VwuAKqJtaLsr6UE
DhibrJ6KrVwDTJgZq2VZnDMSTYJtF9ftfs2f4VvL0iu6YEjvZGBXvdbOAGX5+92411BkxWgc257n
SU+wmmy6NpAPMAWH1+IqPv4I2jLqFpAVu9orFYVHysc02T2oWcCJD/aVyR1ippJpwVZ1mIlEIqqU
g0PMAYNyxtfPgfFvx8VplpqNCqjxFSB+MXeN9yb5Eyg2QY8LyL0cHvUqtMh6PJRwq+PZYbj08pvQ
70Kbg9SbW3Lg39025HBt4QjIGWrIyqXd5lb163r16vTIoVgJPkcePyAG5bSpWlIIxsDB33MDemD3
Fb+TFHm+XpY4wV4I+uMn4Y3g9M5tvSGLutn0AV4GYSm8E/sB7k1jO9ay/reR/uI0AcKc2K312PFq
g8djzJFC/OtT8S88cbC3dKqGKeZzUXqNVRaOe2kl+NJNzLqWsnT1G3x39AJZokhB+I/1fIljSKzN
Afw/xQNcOIpitjj80zjmKBIrQ0yW/LL1yiIoRX/p3kMLJgJoMzIsNx6lhSnfpaSpnaVgKhlZiXj9
KrdR9qaNc3eZjGLJKBKfcUMm995fn38sU7N6PFjrnxPZE7ucMqSspawF1l1zFBAwLYuutNXJ8qQg
vn53icDf1M9bEMjzVUcHGEGdGshMYjqfHjQFIl1RMrAUEvUjGZSujm/EnXtGamqoYQRvjxiTTHRo
vhaf3ocoj8DUmJ6JDioe8B9K6wE5bAFIiwr+UloUEmbCYZEt4nKzLtDHyPThnam61/tFjvfnckBZ
9sVZK6Icu6OcT83Gf6WWaf4TwfVMeCqIsOnSMvVVr1m4dRNNy1rZHRj6exm78zaAlA6EaeLFsX02
sJkWnGXxy4PLFho8z+XsGrrk29gJIaa3T1qKSQozCYnQhaekQjZNPpkEgq0nJKqlinHqU2NCedDC
PmF24WijZgdnlpXUNlDfeqnLtNtqznVKoyJOQiSPfmIEvFl20kxmv8YUvQ9NpMpuLOLJ8Zcdalh6
BQ8Uf5wKbZGHQnr1aD06OEyRqST2+94lTbIS30va3kpkPffM5Uo4DOish7X8dzUSRWZn8oCFquIh
qjcGY/lVhMLivlmpz/uzzdAOqVq41JjKeD/1jICCdGGFFj1vaNUu7sxmGkOAC/GvK6mNP5eKC8aH
bfR73r+vwS/Pn9qNkdsUcn6Eo5TPmFgEFXWGg0KaNbGYwVh5SYqCGWR8bDpAGM0dhHLytzuuC5L+
9gtKD8ZJUMNutrqpn8IsFHRozEf2XB/YT3sFxzi1aGJz7scsKhlDjS3Sgx1lpPc/AXLayWvJG0Ot
vhMb1mJ/VGiUvB9MUclpG3hmHbdMpN3QqHpweHGgvy7upOKbQKV22UpgAaBDGLmIMY1py8xekHcb
uHLrQlOHBLNnUPL8z99yEzyGnPHV3wXmdK2s8qay+JqlvTAk32lzhoMfS0d+xTou1J9IfKIyMfIk
Vrp5GOTe/hpWZIcOzrMyFC1ldxcIlNFnAvpVoC9VIxj+rC9VrhySwlW0XlHFKQMD4pEysL8L3gkH
fusCj9+vk3ppepUFtzYmb5t5vD7A0uIYgbCcUKVBP5k6RJiUZkQcd7taTvzeiNs21ilhMIBqJniH
NRKvmGI60mEoxV0Rz9fLamcSoJw7IfazoQWxbgoCfkLKnB+0n9gfqv8csjwU9jMAq9tTO3sS8iQa
CGrwUGM1pTNVk96pdQetbr/Ip1KZS0MBaH6XIlawtan6oTKH8O0FspCIuuqyahXn6n7HVWiWFIBU
Bm7YIsTGwOo7FbO5WghrVzwXlf20sLb7+Ucb1xfqPBg5iJvLAc/8MrQa8T8E/wWTiuubqox1U6Zx
Kq5aZDDDbrwnbnQd0aVYmQcA81+jrbAtCZkaIhTF0ZsHkdp7fjlSr4dDlXWAtRm89/N0jiXYbxTo
DX7auWwUpeaLZxBmJZvW3oKcV7TAZby/H9hvCnViANDILbHpVsOmRld76I/I/19a6M1X1JP2yXG7
PA37zjwrJkAReXBSjaDQCtNFuLjmvpxdaP/tWg2oPXs2Wxr2h/A+Q/li7ZaZgvPSjE76QcAH7itA
DITUQe+k0kybON3qOVIzshPOzYjPdAD1GkzynwUDx+suXiEOwZsvH0Pz03AZ2/2QDMVIy5xuVO8f
0MU0M147y5kFaIK1GzbcvuPgMRcHNIq9ywDtZxquPzqGmKMWFcnAAWhqcRXaidGANWKjIIWAREVe
XpBgdvEm9jglLOOC65aRYaZYwlYt3y61XqV2YjNEiY/1wECu81iddDEf5uO0wz67Fj8848MRdU1v
leysJbgKQL7pCD+EgOHSveGduOInrEfp9eb2CR0YTVmw6aScZH8u9NWFwlYOad5Vfns6gqa8Q/VW
RWjmReEEYOfkHF/JEOpAmoGIFAPrsL6/5gNhTsUnbnCGMxMnfHGTfYtbQ9e4GFrIMM5UBp22hFF/
R0qy890RpvXvsD21Yq/Es4vzS1lV7wBzYBWZNzekGfx21KAXQYv2jM1VzBkWRJT5Z9NXZIjgWifF
0/CE5ZVtcO30uEgS1mrLqg3MSInqt0zqwwtgSLdsbpZIH+6sIW52Z+aynz57e7kWvnsHfAaiIAeU
xY52aLOavUkmBCZTHg815qhQKbZwJS+A7+q9HnMMrrdWrWTrM0OMV8/Kg4E6Fo+IuQvp06fd5cDF
itpcFiBenEecEyoDiqJqhuD9WdEV2oOweBO6p+J7NaqCqIoZPQ7FnABv2C8xPE3AVdvEmKHnvthQ
MacboPLSOqN4o8CgNtMCT6sAQzovHa4rKwHDizT5FzLRBO6iiRoTEaKAQ41yMOmz3o/L+WVc0H2E
bT3P/98MoXbKislKXczLpOrhMKqwNRt2rudvTNHa6aSTiAa7H4pzfmGWz3h0ieSsBu6b7OMEPyGg
OlfzKLCuiChifCANGnENOrO3f+aZW2XUQIRuvsFGMxxuVU0IeTYD2EVyuTpDo6jcG6ALk+VOcgLD
rPhlsot3mN+4g9PvCWsrIqMeRjiYceHR0BIvKQaJIEmkgRHFiI3Ha1bTsnGvVj0kf2OD0cW5pyK/
ZdPDpRBv2kztTtoY0bQjhw1uNdgUFgDz79EbcpuweF0c8A/TVjS1WzkJqnQU5p8+ViRFzNOtff2H
xSZWHHuDAeu4YrqHP/VrlWwkRoydOqUDzCfeiRl6BScZoRvt5iMyl1DmtiyW6ey6DMA0qar3uVz2
6/wKkc1MiPDd7JjFL7FXtuuokz79531qOq4qfevs7RCuvDJTyeD/sooHgEjh+eoEe2YwA3YmVQ1l
bRsYh0ZISAiGDUiD3awC4W77YE6xdyTgFXThAtvA4oFlowy1fvl4fJ3m1Sk5HhnUFDFtm6SmgGJY
SK9OTZLAE5/nJX1gHR3SPjY/djZ2nIwbB3ikQfgg21u4N9EeRxppV3X/DfUBmGgtaw2J9jlDj+O6
aYXvWGFpQWuVMm+ZvtyLBn6pO04+LFYIslGxKk5LA43H4qjBWNyCSHb3464Nb+R7faejfYSZu0nH
27TgJJHIfowr6zYcBO+yYJgmiPwxqnpshYDFBul834K5t36pfAgmfsPIeLa8P0j3DSizMvTbGrep
RauXhb1+RgAfyZ6+k0IhWMQkryVyc0ZEm06MzpZNp8BFzzhWvBISejMt8Oh0J1PRzYUIXoEtmcX7
iuQUwDGOy9q9rwHXC7m7vGQUf2PFNmgkZm5cn7JG+a4EF+V2mtO5SrmZO2TX1+UWM8f3Jpqp8IDI
BRCMVNefi8f6sU1TL3+J3Ad1dwBaXUgMZNWHBhy4c37MzMvvEn0XPWLZnuae+56quLoiuKNuPP05
ZQ8d3rsV2s3MGjo2zRC0En8CclbwK/v8wyFmN9HR+pW3Z+CbefF6ssU4Ch9A1gHcXhzvmOEGNNuG
ltaxaQ05ECTWhnkB9tZLPcwQHdUdhAXcmVchWNe24nT3QSsdIrogzicdCcUFNc1N6E9WqvejOzyQ
exw7iYD3HOjHarWieViLdnHAVjb/7CdfTylh1pFkrAD3Sjk77A2d1dxtgAWeg//7dNLme3T6Hpl6
L1PlChismBPLyHCSKhi7sIhdMLhdIK+gWABU9dIqb96LTPUdcP/plAtC9jsyAC8AmWUjpgr2gkNH
7OpQcsJBuIVHhE3FFEGEBxVoAKY7rI/PZBDW3qA4DE3GNdgPfT4ckTmlvgtVJMmbOiVKkrVjSc85
oxGgX5HcOQl7cblGE/fWTnHOvFFhFclk2HhSn0CKEe+PTpAnFRa+N9C9/GmANZPnNAMGI2s5Qawv
Jllk+PILyOKKvuC4gOehhUHO8ZPmKLgO/MAw2zQpcY3qgK7TcI7j4/DzsZFuqOjYNcwL8/9uUwR9
zRUsE+LNiuBJBc3pEep4oXiZu9EsBhOs7OIe82h7o67uggKco79kYeAndjfhzmdKABr1xwGnfBir
bFfgniLUMDTDXU1V8GTAGx7HBiOIyd7WYQZXlMolhIYw/EubYh4HjE0iRFfvUdg3H8lF6xKoX32T
rwkkfhyu2roTQewSeUkCBlPx5K+PYo6YVqWNfmIpE/pf0C4jt43q5AEHW6dSUx3fo2tV9r2Rv5GU
Za6Mv29vQUK8E8i8ZztP+W8RtNlnuU1hcF0Pysy+xm1zUHAutWGpZ9q1ypcp/qlmtGC+RVZYezX2
RGgug4DDKfXrtYbh1dLtvTK2OheE7vQ7Tz58kYTpxX3UguMt/RUKeeBKYIH9EXaMI2cMW2ObpkH4
2yqcxEAGFLh+q/IJsCmOUAMoGgSTLN8TTvDAXzz1lQq2SwPPeyb9LJzX3hg3MyJkk89wXXlOF7gB
bvl/xZ2XNMcTKxfra9LToNECQXLL90UW0aYfa5Z36xjJYzRjs7VijKhWEVjDVBk7KQcpXhKP+Ac5
DTwprpONYj81i0WDyhRKkJKz8sy9EaKBOmys0Q/8lNwnwoPQwy1NQi9Oda+J8aSk0uXBFY6ciPWf
U5oI8SemN8ho2sELVsuj8wriQACzaZ/nNxUpmL4e58y1nYNT4yedPAwB/U7hyR2EG5dnrd+aV7Da
HhZupCKgLWLmtY/n3dZbU0/aCfessjZDN0eapah01N7BMBYOUqTGvpEL+7srBVGyDF0pRXyD83YX
pb4MxoMon5FQoTpwOuxKYfWxxIZeodwiwo2DnCmdcY9D00Nouwj1Hfbb6nGyEg8K8ayEB6tv5J7N
Z/1IQQkfRTOBU/xwldTbC5cQ2jz29gD3S2zkSlY4lMcJgtOYUR2HSvDPDFyBrTSAuYcx40NrlS3p
+R47wHqbG0I9juHredR2/Q5X+jMoFq7S1tturAqGSiKyWp31mH1Hcvac2rhBS9Bu5lonwJtwwU9Y
H5yTZef7WH480QEct3eDYAALo6/14b3EfKDMUOsr0+Te6K9U808t2CUVadxlbcC0wM4kKSa2puph
5wKMOtFHetfPHi89m9erwVOx7ea/UVwrpvV62Lx+2GgPdqYVunhmsAQ95rsDlt+HO/RA/+9xWbtG
zy3Lx1ue+h2YRTE3UrRWkedvT2ch/c1SDKQxGJPqXIzN47WzJvYME8qPEs9FzVoLRfjP3VBxyz8Y
DrGxQatfgU6ZELOoRaF/ZDw7MH2cjGY9acEhLT0Yfm6bAg3BH9sKGj51n3CJask2bdxze6K8opwG
EHAhAgeV6aOMFTbyr5/P4Fg5ped9uiWyWKG+maeKLQUZk3lPxrbbzMxswJxDk1YEGaE5oK9hCsUE
lolDgg8xN/+xY9CaonFnfGGMWxFHSi4sJhuO0wYqHwWqxxmtHuZS/XavOQbR4pMNNbryTb3qR7+C
AitJNrZTX+lGrCsY1k42hapuEnLMmbaXeT2nV87oe/+ChghDtI1LF9//2iqUVEEWUFIy6E0VsWOK
ZQsdXxkCM10JM/L7y7ojV4rcwL69ANvb6UFVS680zzh1HJPK+jUcWyBQFIlK+80q3a52qyebVGjv
5JJoawhczZ8dxZBomr6gjcIN+vRqV5DkEsWqK4en2lzYJLYarTr6S41xrwv+GeAlpfjnkT6G+2bL
xyFhDRualdka0E9Q3QQVce0zbw1Gk9JWooTVJfZhDaUnuz64ythIWTgQYykxYxUEK4uLJVmRtFQ4
3jqMhKHqJtm8/4JmlNVNQzrrNdNcesvDC8PukRUMq69vAV7nJAtT/JuyxMXDS4l4rmULuwLh0lsb
1Q2BGms4zJnabbBpICQYfKW0HN4O4VvAgGcHSj8qIkgnC15BE2bTV3xSENhYn89u5EQp/zj2RXrM
uiYMB6Uug46SRS4uWqed7mdjfu5b7DlKae3yCKny+1VFT9MydAcYQRzVSG+c4qLdJd7Kh5llVxQf
mMWuLlrzBqd/V3SRWJ0nPMFtRa5FIvo+us6Mr/9AGem5AKX0K79SyUrZ8SnWjeiLs4lPHgDHNqIL
TrNf7jiFM+zeZ65CUHoBbVK3pVN0LFzOHZWlYaUrFjCuA1oJ9n6SR7DYORlYV89+a9zhhXQXm2Us
lyHutkjPktm31WbzkysNwM9XSHGSDezplnYXy+H1jbd1ajevoypNMFpZeC0Z5yNKpn2AV5D7OuJU
AHobGEDDgNsB1i5PjfXQg13ht8E2AMfizMbfchhNhyTZojQcCabeg6LUL8SidVpAXgIS7Kzbu0q6
CglY9Q5ScotgLVildjg5EnZoD34DpKPnYpf/1Z6jXyZ0O1MoJ0IuKrKFq68DIO85VMFyojRhn46O
mFD6S1c/ZjBQx80DEnx/Zwhuhu7T9OD9wsx/wn8ahtS9vvmikcnQg8SA6J4DCANDdK4ASoA6Z5mA
Y2lNXxqlq8JfXBgqhb7jdUoGE4tyyB4lkJSj4OK9VMiFcfKcBkx2lHg2ZoRwMhaXE1sTZB7FrPPj
tTM+zi0ULzGHdsXtrOYWhjcfH193tv35yISgYBaTxMNzeGzj8EI2rHEnxLx9ghtG2nBzhknn/pTQ
qMVrZ3Ycd+5OoKXWlysKccCaQyqme8eL5u5V0a/mFaCz79QBfgF08f4ooU+T7ZCccBvGmb1ZAZ+i
H6hV7u1ag4kXqdzm7gs15l68Z4WJ11Am7xZEjj0g8O4VmDqzDY4VdjUz3t+03wMnaFzxsrwAPQR/
5WskUVi9UgNz6dn/CWIh4ZgI3vSDFLHZEtW0yaSomLobsCIMfMYQoo6GhIeilACQvgj4Mn9FIu/0
mtvhdIQZ0/KfrZZz4IK7aS6zqhJ87m6T3sCbYl29nFaytQoUHatkAdZxB5uuh+wYWyBpIhQmQQLb
OSiehkagOWZc7qqIw8YXmyB7wbMoDvfr8vxxBxzSNuUVR5K+ATmd75T4pbRsHcemb0Mz9NKifvxc
6rVtDPCBmJc3Y4P/wts1MJ6cxi1jsIxTpk14TuXvyCFgUmRCmZv8BOQeP+8VrSKP1TxftLyox082
AWRHCk1zmAXLw+Mnip7MUEMHsQDCA3DKnBqXZ69omzZXa5nNDqKKyeTKqzITzz2euXKZGopGbFyy
+W22t9bZOpryzWPpnGq9NtQufBKsp521RGaoVPvYi+id39H/s3TxDLT7OHVlqluagXIiN4aUT4Vu
O2F6r8D2lHrnz/LiR9pOYaF40/I7X+VJJJnTvLymhqrbBMEip/Zn+tK+znuAtXOqYXxQJmrdz8bN
IWsbXJ27gu0fUf/LcR1YX25rscSPQnr7CHz6/k+2mKVFR4EkamOXTgGsIic/S8ailr56RqExSEJ7
uDcvHXFUhPYWLlHGyIHJcpyjp9QUDKL9MQO8DaIDmUr91O5sqQ6pwzNTWa8sjFbepFLLT4Z9ZgGo
2aoCYmrz/Ni57K7AedfEbOkUcOd5uMPR4ZlTObl6jpxXkX8M2aFkfmTDYL/HfVgsnTrC77Ad1EU7
eRCFTTVm9Bw1pIG8MAztmK7ZljLyo1MKsizxsi0kIu9IUBolgEFv/Co4zvWPr7lEk8SrIbc41Oj0
7U4o5YOmyPuyh9DD6tt4uO5Z2b42ulx7XeumsBs07fXpVwP/YyFEj8KQA/IhZd5YMFHE63B6X7di
yQumcEV+AHCitVEhdILqccS+QYNLe6PclkAZ/17LIOPu7LBvEP2N9m9W6DzJC+khnfZ6W9zC89Sr
JAFQVNT/tmktIbTCj06Zlmp3Q9mD+E5jSSHM1iAevWNMpBrgnOXr1D9DcXZP7tMmurZDHKOw28Da
id38mODB+zcY8pyu5qc8dHpd2O42P5RtfVOdFU3sVtPjYhGt0R71oL92MyvHuDFtzBRVJ6bKwN0E
9l/R8ClDRAhiJnvmmaosoLtCHldYi5GfcNI0e1CejpId/EsOaieEprj9xXL1mDd/JHo7qFtE4QiM
7GMpDQKojI03/xlptryScO77yDxTubT2IDI57sTVdciZkIiB14FsjgUgcBz3pAkxGl99qZ4qVaZ8
jmEYGsJWf0ZrOtzFMnqNrLafmDYshLpRO8etsYKQkciaLrpebie1lf/T6UoPF1PNCqJAyR73GdjG
BWB0CCI2g7upmmUbF+Nu7tbp+BEyZHgo968j8NyOrjHUr6fmQMyHB/4bs7CKGx8AMG+XStcc5Ati
LCpUKOSKU8YiElwPdMgcTTwOt3O0e4V4n4+GYb0rqapPOZypPBQj335d3oT0//xqFpjrxCRuWnQ0
Jf8kCxYD3mApDsCHL34JCGI/4EwyW4AWXTFrCGf4YsZlu2GNJzTJDqA+drWJ0q6mue21k6VusWhK
HrVDE8VkbWV/FZj91K7zHCjH2bXqL9VUvCIDrHxTEdUmn+IQl7LRn2y+S9fVlQ1sIXV/LYr7HmA1
t+AJs2VrgyDagWVpC8gGjuKG9dsqotNISQiaNlf05HF/luSQdoZBVo+MBB3EsiPPCsAFBpRwns2S
CaTDH0apD813hmPFUsv1F/1a8Wq1CQX+ExoIXJEPv0FIDjvwqxmJlkWrOizkUzWlrR7dAPMybJ9j
Usyi5y43ng/158HW+UsB7x8gc9b9bRxA3IKR2ewoBFjW+sbABHMUKRew2VvtY8ynrOPpRTq3CN78
4fukPIq4xRUfZT1IqpViTKOz+9HK7DYDEIH2MgW2jAyeGHwr5e47FXOjMR7rtHTCZ8eNdXnvc4JW
RvEkuKq8C6KVtskijEnDv04SinokT9UoOTmJ1NekzdIBThiJPlF3eguLjRLxVhF2HTyqk1yC307C
h0WlwhQPQhcUyHlKyHzte9cK8E4evrjAvj2W9dsrbiEwzqXjtfHoqAz0KPX3wcdTiYCngTQtaBLl
f2S3fPwf+jMSL4vJqk9tSmtklQQHmIuLX6QkhIgc0uYzhVZGmAPCTx1p3gr2b4J4gH+w2z3A/8xa
dJ0NWtgAaLxdV9ilmmvSLhrz7A3iaDog2YNzSzqdzvOnN4bqOsUlXnv8WVnJoSH1YdWo9apFXcjE
VUpgyKdsLladtbg7JIV3mV0oqgEIdGNRQ2B0CeihexqHHtergcQ2xAiCQYcFg0TKxEtp/SMPzqc3
ccnQ1PKa9Vmr54k8suS02xA1goyPvqQlNJKqeklLMHBQrCb35AX2/NjuBwctbaXTNzizb+/FYxT/
CyQMkNAERsPp2Lcg4lwQVokEcG9hOWhY1ojUf5mAeKIWj40Zla/22PgAseon8aEEdAOK8iZZUc1e
5Qmzq8lp6OylqVPVl8GHYqAdtL06N12mN6d5yvRE6o96PV15GWqT36F4fMp++g1TYHmsiuzkubP4
iQo/ORSJjpH33k2RcEaxF/vbsAHAgC7W+jRBU00rHDHSGbeUzdMWV/X03Dif2AziuIp6dwIlEROD
emlHaxA4nf1rLaTg03Yn80722GkTWImQtNv2azl5HAxCo/KG9aBHdqtFospJHL9pmKEkFSYc4KEd
SVM9S/mycwLzvaj2w0lgOvQMrUW2587s8Q5mdLGj0WTn6Ee4c77VPntWtxIOubYU1TwoVVKq9hct
yloNJIjXQtrxLhM9vRwEo4IR0J48l1z2RephdalBnBlX4JF15NFHmrbtDfGkxvLJa4qkjoJuAZek
3vzD5stPkAPf0CZAlFtHKZ2xuAawyXNcznTE4btD42NTCdd7DPs4Zt30vd+xVhl7RtZw+qjgAULr
M8jNb1M6EEK/TSMtJo9Mhnz+OcWHv80gseRNTKLtxZxBzO5UW55GtLI4Z24cv75H7nFJrbYdImQo
xOahHUniG6UKb1Zbfdr1Zz8gt16fFkmcsjWK6VxyEeG3kdCX9wWy2L95FjEDe16AKEM5Kn0+4vd/
ahx40diioy1qJn7TX+ZFFKbxFilCuMJ0eX3903J4OLTWE/aipiZJWI+oPfTUmrPpUm1l4OjPen3k
RTtU8hofpIRqGnX5roTfeCnBvXS61eeJqjwNmYRBdl9R0doJWF5IscF/AOhsTJdbNFynaAmzOGSp
OSSmbhpLYwEGTWuvVrEKGakQtaGNbz9LwOgVOMhBWuNiIbwfN/qTIaEwZEG0qxl8MKKl6LQ3oXdK
wC0fM6pAurM4TpX7ccaXxWGv5oIYrE4hs2N+uDCoRRtql/Bip2VNUrcZvmMcuqxV0EhekafVqsxm
yTpRX3EViibwAmwoAhq51TbbLRCJRFH0OVtx1JyK07rl3OV+lSYNL9lr3UkFCDuOezgNUNEBkTBp
onxczRSR6z6KMdhDlDt9i0itvxj4wjHFJHV9p5W/cLdDtW5MUDSBBdnTMTWFxah/deN5eB5YesRw
YXFV8+fu5eYvKePDMfqbnJVKM9WQ267aB6a5CpbvBZPvWllDzomYeuBjt/7l0NgHQDY9MmCkSl3M
/IYA6ryK/JRO1XHEHf2NAeBdSy7IA1xDdDU1ns0KLmuqlpowVdBZ3B2mHyLHz7gdk3vKwmJuTQan
qy+SkGPjjR9YEnJOazcG4cXLqJFNPj8Hxoyx52BUPwJcdbX8cx6ced4YBhazj7oFXn2TjvNDGvuf
On1hqvGHOr1iS1XLSvUHad8i6RWZxYAf+0hGryyHHSVzgZJ/fo5oWoQcqNke0l3ciCslwY+tmvcL
DSt3scaykU9UrquyJPggjct/YFqdigZIBVxQjw/5sgfKaAmyU7k8kpwLHZTobj+uBniIprnV6Gxv
0XRitQr12w69hdckOtRMdse7Vvmax7jye5R0NZjyAaHm7wLfoMwehMDgxRxzg2ztGSYCIR9PL6NN
O4cH2cBvQGd9zy+DgCsAb4YQ0zcwwHVHV498XG7RrpOfQbsrrfcDjS8KIrl9VLIrYtOYhtUCb8Y7
vmKIjDIXyZBCS8wAajRY9jiXXyxByPRbCNnQqKyCR8YsJpZHMsIgnOXZlPGR3QnWeQL84VC6so2/
o7mkcvhtjPPTYpSEyHcv96gKJ5XXQo3lIzYfWga+u++cFA6TR5Fgd2iNqUvSc5xncFBpTH7TYNWs
zFjwdSnzo4/TxAR3PoVULI5AmI36KtH3Cf/9oVhI2fMjaKPdyBD8dv8FvJR5bhiUeag4hibm2lVE
EY3laO/m32fEcqPyDkPwkjZ3+IQjtrLhp9JQH+BABjQzq8lrKRUbKDzybmFjlsx+7cesMC9EZGhk
Yc4sjY19G1eltimE1lNhMBzhCWGUT2uhDotR9+i0H44lhXwOanV69K9s+BjLRVMPGd5GFl07PK8A
io/WkQywJ8sR4ggOWShJ+RS1WL2sdivG6Z+Ke0hwxIiESQVlMeADFEShRjkLeplQ5/kA+3EKqRbK
fap2fFcLWWSnoQAknFi/Fx6h3iR+/kC13fDUyO0seD/k7VBkFg+kAAEng0MDYpIgtEPRT8RIs0VE
HxwqLcnni/TwZXpvoeZr447+IWCLPTouwrF6wavEyX37lxdH9qOc4EpH+AP5L1PnRjk19UqtLjEt
shjoRZH2zSdNsmg3SdJaqzxYBCvKnal2EpzdFkLTTWH0DT3cEZGVpXMCQG91wTSiwNaMGtgRsbSB
S7rfe8MEOG3YBnQgO033z0BYGWfA6gl4sCGRqWQH4BWmJ1/diFG5nwAtNo49Rhne7bNEK1VR2/yq
ojX+iodKwFAQSifWn6x71FUvZETep07nbiSBpNcDXRD3O3/Uk+uisD5y3p6TsOK9rSa7ZsPVshCC
ru7I+LaOI4TaJJ5SMlUftHXFnlA+6yicWEV62pSJrDOcbEkXb0AJK1YiUwPSywfHhR/Y9YWW80RI
cBJjfAybQUGR3YTUaw1BRaLrXiYxYqcHs3edEZ7V1UkGo82kxXVN66Kw6WUUlPVZ7gg5s4P2om+W
WT4wCr7T9hTj0D1muz8nq86pybkPtHyzB1AR55c761gbWVfDPA0HFohjoNokG/veAboYifgyYJeh
If08cOIzk1xhXlJAfJtCYV521l7ZWmBkao0JfnNNMn8zyZulWw29TrcRryPSmnPRtHw94wEijvTX
eo9IhsYf6TIgwZ4yVrsaXBrr69t3sd2ynL0O97ckFjNGG/OgC1KSENnnI+NVrr/8/DN+cCEIYkwA
B3rvV4MLrDA30HuusTC/GsjQbEAceaQt4Hz6V/5vrT9WCYqNga5lUR3qMVV7tJrTkpuj8G8PWX6R
TgfVZta9zKgRpkk1pSv2BClTb5VFez0uRAeQgkS8VEVeO01g2PMZ+7CfiS/Kl6Dxj/dVIfHGo4B8
99cTsw9MYpyjgFh0wCHFYMaAD+eyV2Yi2nJZvr+z3nZWNgutuic3lDHpyDmrIdAflCV9lCvoTdlm
lPnsiuhscNLc8fb0LOkXhfaylVT7NQh6aRx3VA/KA+dYkhwyVGQ18HVJp5LBY82+TT+0PZn/hEzD
wbV8Xs9PVi78B25aqf2wNVlkPvsxELS8GIkBAwbF5TK7z/or8RMOcJx3FcRgR9f+S2qI3usFxJB9
g24+x194X8+UrnIBXCIVK69z7c1u4xVughZk9wiTPZxyJZm568cQk24MBa07gKHzQjRl1t2GqtTr
rajs7iD0s9Emcg0wb+LjFLClfdP34ihz/CB9EzWW4j5PKzRJSWY2hpAT5MavAX3qBPA7rlCy01ph
9iJDQQgPcQWzQ8Zv6n4ZV3CRZ8irRQuECvcMRhqrk1skyFaoTK6lpmQYA4pGq1JzIurpsF4rfY9U
pCRpTBr3CtzfTsdRKxcr22lOuamANjOR7ianJcpx9xrVur0WCxM1DxJzTDo3NBBmm/VaBJViQUpB
RKO39vtt3jr7w+oPNUrg8V8kxinzGJasNKSQxjLKpmqPvKs675kCqbl4T/l6v6Vc9gM5L2sIg8mt
nt/7HV0uJRVkBCSOMuuszbxeUZSi90XiWxoAc8xSXRusg8aL8Tf2Hc6Iau5upwfNtKPQi2l8DHiD
GCpuiA+28Pslu8N12Mdxa8r3NhENXRNNhZ1d2DsI397GK+kgmT/kCBIzgT/HgOrpcMUd9HMk1E+1
l26HLf3RMJbt1e4gzVryBPp4v7gzJ8R8BpEEGQJUM7qv7Lv/uRMXX897TRw0/2M4KcvDhQHLjAVd
cHbYv95qCAxtIUDndn8DuWKWIGLUYeONElxqbItx41m/wZGXMWpeh25nb1oMtVpX1nft6OPV4V6e
+cUnCljnIGv2CuJU0tsEgc4Eie6Hx9T8+ykCa11gIShiuAlVIJgT3v6lpp/yl+tvb/Ejg34XJLoR
pU8gv2OW6NWHQ+AXE4eK4o3UEicfYu8s11w8BTiT+/IwPetfTfP0YuNaSnJt0CcVW/LXK4OKAr1Z
ALSicKD9Qw8WJnCTwpmQrwYOoQ1meqp6txdapN2a7UwuKxUwUVlpyj4UJcREBIfjLFHwhp4xcW/z
1fXrbx1dsT4Kf/EGHADD/fxas6R3QAAayYUo0J5J4Q0RcWfXr+kDM2JpZAbGKu1/IJ7kgQ2EyNJi
YpM3UUK7j7OqesaCiTDg2yylYoc19CcXkZE34gIpVTC4OXGgVJI+D8ZfSALgXcfeaJBrOFYiUWqr
8EcRLG6ZLbLVq/Hjbx8kiO8XmjYwtLNm6m88N2KJ9Wtr2OlCmbwBAz6XaWRGAog4Q2NJIsel1ZHr
seOPR6Th43RvCNiQuEWBIyIOc8w8o7dtGH063Z4q6O1LqC0oaKwsNfpgUrUEWHMwQlsCCWSWuH76
a6uwAWoFKgstBfExdL6/AhcK5icy8wtSIPNVYEVZOQuK+pAouS69BMXyjd3ve9PTI/3oNMmxOxAV
CwCacI7eodzllPX/Ylr9APzK0t2z1trHPag7i7mGmTWx5JrLSS7EBgkNg+9ngYDz+vTU4DOAdtEo
Q/YviyXR3ZznQkLjfY9RY9DHEKU/H3S21UBPfPunkCOt/S6g4uwtR9C4DitWiHlydCI/AXlq4bq5
lB4BlluJCex9FQEQ6X9Yq8O83XDxPJb38RQCBbXFQzHnNTHT6Dsl3x64K8tHplqnxY99WZgImTSH
O/VrjggUz/lDIJOeB/nR5QbRATSlYV5+feqya0hrV8nbGt9XTF+4foK0qA9gX80lD3n2Vs2Wc/GE
bKE/qiyNVHvD5jHH9mzsYVDHIgRNkOHXK8hjlc1BI7TEJQ6K/4XlCAQ6mPki3Ry3KlixIFXsxaeq
IHibzPZTn1ur2QD1sTTS5JMhaRaIJ3kxKq0uDQJUoQHn6LoFAQ1BkBNNK37ZMcV+5RSIoCGdxbcA
KADaIkmofm9q5BR0IIjDB3TX43+lmLxBTS6Vpu+/737wqpbqWFQ75FI/3jhNwurp1rIar+QDs/cC
KXJYg9zb/+hOe4lNBmKdMdbBtMFPLpOPsFKnBnq8yNYZMUXoJzcB8c4wHkfN5ECEkyghhVcvYWEy
I2HYQpGIQzc5rRh94IUVZhO0r4ynSLuH+bFq0QSg1sgzQqIP/kcpswm1MMWuSROrXbqE1s7yfiNt
cFuCYAFRoFFvrlWgtP4MFz0waFHD7THHs96IJz2FuaFOi4/X6Rfibii0YUt8FJfTo/g6/LIAliDp
XLwEsdB1U7BnkHxXZdkgJDmFPV2PQtzociCPVm5zJCzSHMvc956JyrvpnkglB+KvjQ3jORDiIXuQ
zkG5k49rljhi+ecZ46dUaQXoKLrfVodng4jIPXAQUi4SDM53y2VEB3sqsUX650+0gXj/vzbDiamv
NGrqO9Bvk8uT56HAeldqz0B+FZicGqTqmSAFYD6NQoYfO2mWNt6w47uiNZQIZtORt37I+wHZLZFa
O0rR+EV+KFvJXD1NYIIevpvsW2ElowpHR2Y5HipdvYuQOGnj/OJxXCOvOzA8Ja7nY1OWxzBpcz9U
ZIL/2MJrEZvAn7dNS0DpOMHa8cUOaVkw0wPO33ITXYW5npRSt4KF3Xeswb4KZRt5YG9iiUHOXpjN
kqD0Cgf46gpm4tW1RbwqVGo9LlpScFWC6qWJjwbb8euSzhedk1dUleAxhp1QuSqpzdPutO7XOvuG
c0vbYAa16N3yCSfCIgUMYiIq1P2OMr3a+TypUTwV9JgWN5J+62sSH4s0x0QqQRrFZ/zQ/SOEWlNv
+kiEU4sS+Ha67XmOXT+qJXJUpFn+4IOkZqys1aVRPusCM+mfta2ZUGeewIKCWgM6M5Ljcnavx12h
HGBuv6agSrU/cP9zZZjL/VBZtbhizb7TdyAiX2fdvLkKKv7SzJpJf+kxeGzFJDQU9O9HXHlgxvGo
obdH6NBMo5COY+4jGp5ZjXGI13PUCuwTuGBUV6LT3bBShUUwZrBQjliP3gQMr5GNPp/74m41up92
ry2hD5bm9uiJE4WSku9dKNVZrfi/yZFPwKNwsmdEYv7/j4dbcjDPKyw08OfHh0bVJTgzJeznpRKz
kktIZUeh/uBPQyzSB/B1PlFtkIq/As7gZULCqaB7QtEGcAcgk/REEwZMX4cXT95yV9Ivi6V5WmwP
doCn/xFtkyDijhIomKz2wjMgI8yKVpt/dQPT6oqJUmhPuViix50VzAkcnMbZBqL54R6jJ8EVhnx6
jmt7FZhpa3PGcTdFybVCruRHw4bAhhRQjG6KTXPLNCbZ+BbCkFvO/hXKrA8tBJk9EaSRUSoRNmpx
iLZYEplR0iD4eTRAp2KkXlKbpEjqjhb3B4tQRK2LaSgcm2ZkNJX6xaGZPPQc4f0Ayf+H+jBmlOkc
B+ITP05p5oJ+BnEWrLCTsYNIbl4a6EG9P8CDg62G20m2aP+eLcu3RXTH4DBP8Wag9M1cH2jfFoFN
9hIgI81/zH8YHf3Vbs+r9paVuIKBOzlxXcZaqsJ+CWP7a7TSKE0Mmpu/bX/+FA75C23xvppwZJsm
nYq8cuilkgQnFjsXa98BO58fL4PNgFJWROQiwp6t88dqJmDwRDMr0IdCQctN8u6mvGynHf8H8mnd
CaUWJk+hatH3l2ku/eFM/ya3X9LIJqiDR6pQdxv39yjK4TmEj+J30vAwKZzjUiswBWQeLcZ4C11U
fv12mYnZP3l6O96ChC0PNp/D+5I2/LuNhkmHgqhSiFPkF/wf3i/txC4Q60gaakgCF2GFDFHqvVs8
cGfR11pY5IqQkb+06e8hEbYxNeuTL825w7926oYIyUArulX/ISLcfTV4Im6n6Cal0Scv641UfI7J
8ywYRtjmkNBNPhp0Zvx6k2aGkxsamHk1CvQIAUuAwlc5HtMc7ZU+XERD8Ttbg6pONUGTzVnvJj+G
PrIpqHBBliEPOgpFw/FqRfKdmy7wUt4I1VodjFyOD+ec4mFcd7eS2sZo0VZogMIVoMcds2aSOAxE
WEHns04RkhmlwaLQbgIxEBY0zKTKzF2UJf3Qnzz1ohftTt3HjWoA1DqHK65fwaw6VaQ+wpW7DIzH
KYtC15JEhtGczUIGx0ZwdEjwp0Ohs4I2vqg4xaCB2KKdxIJFB+AhO3jVGkJt8IQrmDL7OXuKjdCp
XdTcK3y99T49QqALsHPfjY4P1SaiZtc57etBqqbf9JM5KvDPz5k8iCX60yrPP78297gRkhINzpV8
ScchRR2LwkUU9u3VQQrZr/CqDmkw/L3XXt+/rt1iPflGsjlHqnHIRwhlGRypMge7KJR1xATPrPas
7xryApr6cQdPRvVD7tW5Rl/f84l6XUXWGIFM4cveEqLTEP63ZGKbCrDU+MTZ9WiSvkUllA4uSny3
uKtJ6ANd/geLdzbCDF/+REmKpWKDqNM66rx2/7ULeRFT5xAfYihWs5y1O+T/+HcmRsQYbX79vCSa
Y8Ex/y8NrDNizbppGw7wZ1ro9akdY1jF24z/7ACQYRrcNYYedwIRNvSu9OUf/K6v5l4hjRbTm1gD
qwPMXg6zzAq8UPTMeQa29ZaG0d8q1Ciuwp/PGs8k01kO9Bxa1n3v3QO2CUVg1nb0AI9PmzvlVxg2
yZhVWElbjq7PqcOOLF6jgWbgwGEkiwpNzZyb8l/trOkjjL1DI7Kb8C7DpiuPXLqvQE0CGg66mrMf
ByJRNO6FQaz5X50foL14IFWS72p4aFmRBJ5DC3DkPFeNDTiksypKBvfvP3CKv62pkew9FwZbfqM6
7w4PcwP/yOgIPsdnBOGmM2H7Rh/iydmtbsGctVy/gDkdLAwfNiw9geIaoGVe2cz+6GbNPcvohEiv
EG09crmVAIb08w8YJGq6sO884iN2dAAWgwvtEE5dyTyW4Z4TMQG4qNnKX7P0tWslQ5nvc2qA1FU5
agTk6zSJBHi07fHlavNpGSNmdrHq+JkU+UdzZQN15bpyn/7Gep4b0xP6wKlowb//dwxvIgtYZTf+
Zb5H9dAVMImCN/kldSd2p0JrCIb5S8E6AwnNtKlqeLStENs73Z56cAWgxGFDPUmEHSwNBU76erZw
1oF/XnOQ1RfZKKRCWCGSYXZpj0chuDfgY0WcKD7/rCbQKSeW7+jSBDGswdrNcJk7O4IEbjqnuhcU
34CG8EG9rDUCQxbhRVTry5Gc8gx0YK+mSfa7uNUKXIuDu69BAA9lYSCPtkVoT7iJlBo2GazPTZUT
mHmSUUXCzovwrS2mvxZScdG8DlaCBExp5FO2GwS3M/6uVk9txogKaqOE7Sykjr+Qb54d3u+dVrE9
k+zEaOOC38+UBBYyW0vbHSEuhw9SRdt5GjNCC7UuSK1LxwPNhzq1Ndvp0nZoi7gqJxeEuB56NCCy
SuRBg9TxFWwmSg6EZyTQvus4ElqZQf1zHud41GVsTxj1mzk2GOWP0MNr0q8x7sfIq5p4NV3DvLz+
o2wtdR55Kis8Rf8BpAxMCsYjBzLXlOwNR+xgMxMkIjrwsWus+qrGD06dwSqINhvBkU5Cj53Elk7m
71A3xTLDvI7bsWjdAMHyyz0LM6+yWtLKd4dTlLUDTK2cxDZt1Tvzq3Tvza2f/+jrIkY1G85YP0ps
Y9q9w54FcjVRpVf9SqzeilRhhLEIjg8ukVDuEK/jZ8cVAZuZNa0/U+gnTX0Y5omaVbAMUtrmY+VV
g0Bbx2tK/XJnCnmTqsJklLg+/wBUO3T3KtJX97645qY1NWk0coCYrfxoomxJI7Foeyo5MoHohjKW
2Sc+mIM8aoHzMyiqxgJANay3RrGUBj2ep3V0KnNhCT9WSNPeIDkV0DGy4q0i9ATe+cPfH9PSSABb
pQI1DtnRc/ntnYtFsC/HAQwyp5soSbMA4S/y84rgnGs3kzIRoCYMbDjlzoIlWufgby9Gb4jZ8SF6
b8SYZmRP3JRTAyjCUXmNtVcXP32o87LSVoRTQPmhw/DPRXAcvjHg6HBBqZC3O3dpuPYKglIGbciG
rkjtj6+STeG3t/vT34XkHOTmrEuEek95VP6a/H4eruSf9IeyoAjipM4bgkce1haPnQRcqyfCTdRh
MhC0HVsLkDkUZGm8pomcT4/M8RDlLOxefRvpmoFXBUGqooy6FvH6HURpztANe9d8SiNsmuSmTeGl
RM8nkf0WrFptKigPXH7JQSR4ZakIcUTUrLey1kbxmHMR/+T6LD5z0D4PSO/lHkwsgzfKs1kMgEFu
wEjBKNLqP3sj+WnoKtcqYsEaNyN6yuG1nFI+5f8dHJIkb+v0ZJPN9+DSAYLODHalwgVL7ZJOFOOz
fegNXcKE+JAvXvxT4BujTYcTk7nVm5FYNDHTvD/yK4evOVGbUT4hk2ypUpf8FohHWtz71iIfZzlR
DaO7+jEQ2nF+PIeW9cZcCR8JLt95f8hfIe7FCh2My1XdipTxWepq/0ZR+mUA0HNkcUTSwAwRc26G
F52sJIl+lQAZt4ELfZBJ9MqMtMdLjoZmWzwL61jFn4uDjl4WunOd7rm4APnnKPOQjOFbcxpotTJI
fWhnk9ubUM352BO0C7Mq/WsAopT6g4BUKpFBxhoZHx1+H2TXq3BfP0D5FfK0YzQ4HVxcg/ARLgTI
0NijwxEkDcB9x1KqqUGrbAN0IilepulIhgeQZAaopWQUYJ71l4eNNEzoQ6tDh93SLcVqgNqrStMT
Ak2HC6P6yDN+lXXTIebPN6AUmLT1eh3S5Y60RDOH3IX599/5wUsXLk+1tqyT4QTPjpNKXMpwSRKf
A/Q9pgSDoIFOv3rL7oiSmk7TjZDbXaBapetW2u+7Xsl8CasLV/6sbCAeDTebvDTagPNB9LaFEQX3
jil9jSJI8H8hRj5bwWp+dDu+B/IoU+4We6tS0yjUzDXdAJE3iaXfH+dmiZEilglBnvczeeUInDH7
cJybp3oZy9sT7YlnKx9zUL8ukl6sEIU31AcDnAo9z8VpFfoKdPma3VeIqXd1jSszBNb3P0bEoLzA
F05hkH2KDfvx4SZvxBP+IV4v1MV/BNMLzv3XwTFMAAgGDjFi0xA+UNSD/+g8cEvzF2Mp8gh+xjkp
XU4m/4sx4bJuvLfR+QvK0XrgSz9vazCKpR+Cnuw9kNDZSNwjip+vWHw6WZk26T9uiNs9jui7Tpkw
v9GxkJ5m+J2TM04l/jK43rkElFZQa4/8jvnJrGJ0UKu4STEZ1Sgfw0LSp78w4xrcGeZGkI3DMYxM
Yvzao7gI+eDTG/OdvS1jlcMTyXubwqsAzwhnt220HhZi9Gt/aO6tatuMkZo2lUd/J9iXvu8El3gL
uWoXqLASRhye08QbPGQ+7YLDLDxgX9mYwOU9AL/p4okBP2h+UhTWreVEDRueWim+RO5/ikWEA+mO
p5lfRPTfwNgMTeqle/gDZ8Bsb/GzEtzTvmwy6D+vBFYiPZy7Rq84qHh8/CgkNukqa/7sS5SYm3EW
+xrop5e0h/tGOXK39imxNyQc3Fzogl1jXxZe47QE+j/iw+bUxOgecLuExJhzgbbctXC85FrlBnRd
d9AQLpIaI7sO50J/qcdlSqbod+n9JGf09Rh3pdHDeXcaoKrrcU4LDJpftWE2KlxuCz1BksqG7XUv
RgBYbgh67wjKs0gPzGtv5MZhFUa3dCz79b51ccyM4ou+Du2INAMboJhmD+5h/4l6tecQYCfp95Af
Q5eC0Osa2kUtrtuq1iA8nVtl3pNFGtvGJKleOZeyEnsKVEIPxp5qNUjdqVHC8lkqsRhKIiZv5OLi
Ht2jnfooUqoEcZ9oKqxK2pBs3E8Z0jjXR8bhDObBCFqKe2g/NHfaEin4ZMVvZuI0DqqGkFWgVFrF
dn95PpDg8uNMS45eLDQ1Zz4FvIEO1wWqLO2uOL0Jk0CZySf6+dNEyeCMr7pBNLH9rR0gNcsYY98c
eyxxbGVRePYpKJ1dT5iAItSAlhWak2am1yp+bSh2HVpLvNarx0D4E/qLt3cTE0z6lc6hI29Enweo
fIkQvwaTyTmhU5TxTx7t6rhaJY5Xda0x3nGyH7xyN9ZKl/FnKGLt6tIi/yPjCfkpX0iKBzXK0pVQ
6s8UxhWwSzPZC3zIr0fcm8EXqw4VKQ+voUy6Lba7tu27dzzLlGWz3W1IMM+gvMqfcwKTALSSd16l
+YLkVzSBly7w/hSknKu8PLdefTiACxZTJyaQZ1/noBt6BTyJNbPX7n9MdBTRyMgGtOWnf4M19ZVw
j9R+NFBSqxLFuxT1H2qUd3WSGO4wuiEfCflKB0CDuIfw/R27rkrfn6hrGKLissYeQJkBKdvkFJO7
75klFw9jVC4fC0lYopAu1/c3dKm4UClLxzOTrxv6K5eycxFcZReaz9Iv1qTDkOAEsz4XnB6Smm/k
RpI05I74LGWOh6ieY42DOzOYXu8DP7Wbv0RGoUlsSjev6hKbVk3W7oUN7dTA2iiUQ0e5LII4wXNB
p1BXRgrhTTXVWTlD+MIIyGosee7kEil/UFOrqHgfXUe7mfXwblRKB3xAtM17u98qw627Xj0hmiOH
Nj7BLFZYNQCF8sMwuSoTFcOmDZoXoH7aZNRabxdB2JEtvWIBxoez3fxjN9c/IGybJpbfWoA7oG2r
i+/yxDKiaseLEpsJFVKhluOy33l/SVGtxoe/nmZtdO4MeswxK5/5Lo8NKqEwgapaKFX4QKgzSXtF
/AxEc/XG2v5Dzx8fJ3pDH0ASyqcqrF5CwQ/TfSFkNv2RVxMO2gVU2ArnGnqU47Nn/DBfY+1CyjSM
EXPXgaVnJQYNZJ9odp6lWjmse9D6KiRAgShUKDhUmty7+ZMA0MPTJw2Fgzl01vCrbNThqbJnVL06
w8dy4bN/gGBYM8yU0BhfXAZf/YFplasx5XTEjyOydwC3eSLVUATBHkHB58Tty4DKecoUuZQL5Jgy
hHS+8wBSXFgHfuApHTkxRdl/iCW/hjIfVLd4sqc1B2jUtRPqxSlswXzNzoyMwSdEgZLSUjQxvmhr
yxV7NBWpgM5acfr1vv0pZVk/DT5V5ZpTKD4Jz4pDAN7+B3thqCdzWKUBfgU6I+poqT9NuoeSfKBq
i1F8X0/oS/UAbHDlDU+dtnd7S6uS3WHrTRMDXvQIBU5BAyUFF6Jgr1PyTwj9mS2gZM2ftjOZJdEk
fttAFCQDo5G9mbvalH30GkammOnyrRh3nOD6dW2jv2SUyXnu1P7eczjZY7DQAS2lVID97f7apqFE
+g912qKACQJAPRVJKFK+/mn0uBQjLOrGmxsK5NCduVYnqFb8LzgTZTDIbqs/+VTlBC3VC50XgqOZ
faWpxSCe4zGFXjK9iy3trQp+ytpa0rnblh+XeR1uQ4C/g5SBYCUvr31NcnWtDCQ+lXZINLGAD+x9
RpoqAfN1Nk+E/d/xbjlqsd19hryupz2FFTAtk4f9sbNbFKo8SS2QozXTeUmfKaXWy5BYsQn2ohp7
E2X5ef3ZVpDv+UUo4rWBw21XK7vlITTYP3rkNLG4XgNzBYGP0WayuEUat7m8Q0wPuaNFCmGUhQ7p
GotI/9nTglE86XoC4I+aXtrnx/6GCpj9GwrXyWztJnRwSUoxK9s+FAfVywTwB4LUsRZP6VVCCwZ5
qKuAeYhiFKNXD5hRMhBt/ShqcS2csPdnKNwRIzbOnFpRyaFBYgZp7emH0y8I67AOnGVUwjTnZVcT
1AeyZX7CK8cNDZqSqCwlW9M/vaD569rMVogVOPvpiMWAm4RlO9rq1/Lv4YGCT7wXwg85K+xst8zA
rWECFrATbjuSHEKi/gCcRsXa7/RQ5mtqgGKfqeWgJNOZsuDevJXKX6GVOw6P/A7vBHOZXNE0acTA
9IMs3XyGDoi3yE8uJCh/zfC0/tBS7fXeH+oCUe3BZu/UyzJyJy1mJWcqVmCFGWkh6HuHNW3kRxHm
daFqKKywj9whHRxvcZF/5q8PnE8CAniRWgTP+sAwH4QuKVmPAr0NVKSeYbQT/krkC925iFbRasQI
3PZzZsqRUHY3sKMPKQ9v6QZ/cBDS8MhWbzIP52glpsjZjniVMA0tNRZ5h2pjdrQSh+EUpVU1l69Q
yz/c3JrOMoH4vsxVtbSRje/0g+QmpmcEVFO79Mkjy+ED2QyZUDLzD6shFS3QeaKmQ7E5u7yYBdWX
v/Dt/GvOJNWXqv3nFV5bWqZgbrSHsI6Y7jjQ9LFxqeYf6uzp0v9NraEeiZ4ZmcsdiIjdVg3TpdEs
plPZ+9do1RL/esbT/yMw1qIktQpYmquSBRV1p9AGqFStRgBigsTiBFv9rdzjY6a6AFK0yUGtNAM8
bUICX6qOmoztQrtuJ6h9Eh9yOHxlXdmgEdyuSI21OkqxaY9CmJzhBDoNPkT8zw9bTPCB3fJk68UY
ZsGWUZ52HIMoLwJ5d0alsj8T9uNeNTsgZkTjnsD4PlaMhD8ejN7QA8R1FY6fjMfo67JsX6OAVKgC
Dc+I/aVYLVLt+FpTwn+5ZQe6gyD5Z2zb74P9I6BJjkEGya+35Lx44HH4gV6U+Yl2treqNm7ceJQ4
2Iur4zhl4xcAiloHNm2HFJcqVE7BlJgFP3ZUKnQ1UBYJoipGFOdic/qOHuoiw3sZXQE5UFb5gW6v
R+sZBLb9jyueMlI+XmBWsQl39DZMN92QhBi4Is707+MNA6sWClik5L9gTfJQyYmsZAqYr/XsaiVD
arD4CDoveaVNR5QivWh0qeSaOXegHMcZ4n/btH4Jr1n6bTxTHKrGtmFVu0WN1EI2j5O1GzfTmUNN
WgijijOFV89Ma7bAAYxG24Pvy0hLLZkB5GSdxyRJmhlDj9wXzxj3g5O+tu1HMQ4zLVgvQAM9wxgJ
z8KLKfUd8RI49hVaZZSwhklb8uZEil9bSCunb64CqxbycIWc/0QeTtBxbdyH9mkyASmqyA7Y8LAy
cCAOlYwT+dyG2k9HwYJLNXZNidl15xDxRaZqGSahTrnZ0xvcspF2Tnh/giBPk6OSPWAgOSKN+fF3
Jtx46hAo7+Jw4ROjGMKDOHXhVLMkqo7OYzYcoAx6UZUs0rNlp9UzwtgL/p9oc8Laxo2MYhcCXR1y
kHD1ZRzCA+gpmsAPOLLQFzlvU+7I7eJEbOAsETZMwUqxNc/ZyGMHOEMT+QltvEpEBN7/KIVrMmiM
okuoqwZh+5IE1Rc61fpgArotrPo7yRWcepR5dWBtVWthFY+NZdgpYfoM126ZqsfmN8OeDamC2ZDm
1KAjPnuLpea3VIu3vhD+FRuSlK91kj4UnLEkLTWy1/LPLkaIcT/I+fswVuVWhXGKkR5zzdpDdNRr
HHurc87OV16ft3HITBMCOFhNcxk5lOucOII0sPJfl2pV24VAT2zDMHEhFwvnI6lFk/DqedHxq3n0
OG7a5dVsrzoyg9pPN52xAYt8QtO/REX59czVRm4w5QvOEqPLplsRJb+u9im5ee+dfTlRbqbGmUlp
tYMtLNMF9wt7PWLze2FcYmLIOEz9tal4hh8tFpx+8oALKl33KwnRBh7EmMM5UcAOOtTVNXekT337
5TWx++Rgf2Wy/w3L+U2Zs2ZvR4ytUNZTOI0oGHC5XUpbbXWawgcJG/+N+wmVtc3gTQjqUUGvJg2v
3hTXHnIVyebZWUwnq0lRL1Y9LC8QL3KfUtG2IDke4V617f5K2muxIlWS3z9flO5IBa3zfDBtO3m8
nMZT7zD8ft0fOKkc98fFp1TKhyZxvcwcNKoorgylwP7KC/1HpoLRmc93bg2/IohWgHGnRwz1WQnZ
a9ZVu0KngrSn5g/HfxGuvdrjTFTJyPVkItUjGb1eHVvmWQP7jhDoBVs/ukq3FsAPcvtMGa0+1klY
9dMaY3O7lW6vj3gXeBvV3S206yLisGDn0CQZqe887YvDP+zA8Qe3KmnBxcXo2l9Xh/+2XMcfRTKY
GMNAlmMOJKMPpELwnkLEZ1ldlSwWWeRTTDjiqm7GnHdwh+tz+ctRsPhbQ+Uo+dy6+0BS96KgUmAM
aGrvEd4n2taGmk1sIZeIsaE/U+zqbpu6LMuVb+3p8BDZZwwSPwDO2yYUz3KbvD5a+0/PrdSQsk9s
9DwPmdszrCI/2GAWSj+tR1Gfbi15IR1Eoy5JGJ/3dW0eTdE2MqunDm7ucdqeuEIl8EyQhzXdX0ND
WiuGyHAXBd5MeJLX/X1c984/FPhq19oLjPTfi/NjWPhT2teoTV+G5PgAyu1eIJNwYRhwPXMqv6bY
a8TfWCG59XD2s7fzbmr08wHzxaflxEsrO8HM97fQAtGzSGn4JI/lrYwBQnB6BoxGsuZ3u4czfjoL
e7IqqWwRf0luCRZUKOY4hAAuspnDasrp1bk7BSYIEU3YFHxF9U4AhOHlHzYUxiCDwqJEYY+ttsU+
AnlTDtOWZBvmA4P/j7Z2QW+QfPahqOcxVTHaM1Rlh/oOd7/9Czmj5QCSTExeqVlm0KHK0q814fKr
mjeCWkuFIwctbHDMuD/OedAMVa3K3Bdory0eGKyWlszZqHchL9SF+4Po/KLvu+lkZTd9r/sIPHuP
0vBJuxIX9hbtS6DLsEJiNv2ahQ6xrgJuHWv8GVUTiFTosEMjb1GK42MaDTLoy6iFUOwCzoVlKeGa
6OyFpgDSnWDjCwmqmB9KH72zEthgmYRm0eVeARaLuf8NroLyceFsIZrqCAugmrtMRztvNcztUjc9
7WqZBl9OdtJle+s7MjLzEgSqFHSTqGC6iggz4dh5b8pffGGs06USBFS/gjxjWMAWwm2MGCKrA00V
az4VCjjy0vcoOcr8qrDtNF6L8irIXBX/OqHKpw7aligz9TjhgfR/4iIK50TpdThJuZOgi/otJaZo
t4NfZ10Gc1BC8pVzfFlGSar3tqkyuEUxys7zhAhwwGEhBNJE3LFTFLls/uFgOMAxN0jgdJVEZwpQ
g92Xczyb1g8Hv/HylQibVJsYYJQtJDGWvywBMdTsDNkQx+tHOAPOn0G+V9USClE9QW4IQieAlpbG
vKgu7Y9P5cHPQAv2QjqplwEzTAPx3InSdB2DtcT/o0AqzOvLAVia5kfzahofe94gUZ2uSa9cStmp
rwtVgfM8ZJmV559hJUgUMXRgA2/BqPhkGMmksrb9StUd7sAFGOEzCby19vGaM4MbYALV/vV5Q6cs
aUMRrxFrogI+/Ba8FFkkxzoCHU/aYItVzI2ZD09vgYplvNucOK0of7EakJmIDmqnAGxp/oK4ojtw
xwGTIDvEt0wjveBmNYKTU/JZhFfLOHoPF/SQnccUvCAykhdTr4+pIcH5FJWwJA2mMLvlIwHCl+tH
799X4HAxhVU81DTg+kSIQ3DHmlX3eKmxL4AjQJKFTAbhwcH+2Lv16VUjXW4In3dVm+tZWbDfnf5h
82DjuplekaehmcUgGfN+2+bwGFHH1nKtC2nMA3qmSFrA6iP9NBi2grCyCea7wOnVBMYR5vkcj779
mOn9fd2VDHKrmvDKrI67huoJyCm+zLwdWWb83kfTdfBGqUwHjfb4B9JeShItvscy8bkhfXFoirQA
XsXg1zelKVBp0bKcz+6dGyuVSbE7vu7Ya9CNWFNKXUgsMxEUyXuj5RiwC2vXxNJGmvvnENXh6RK8
86ADz03DQOJ72XoS74YpI/e59r0E4e1IKYIXY8X3Kfr1DW2bmoWxPYOIj8V0GBd6TBr7vGsEQAoH
X0nI9H2pUjKsbNz1yDd6ZKzb9BroGDxuA+7EI+YPfm/8BJ+HM2GBJDGaTvUePH55jGC9Pbk1is8s
efR7jmp7VS3ipD+R5yXymb8Qy3HbwexGKHEitCKM8pBP7jvWK39GZjQyNf8vwVwu3HKi2vpYGJt1
KfCKV4llupj42VS+PDuJ+3aB6EGwHkw4HRuEpk86qodT8zto7uNgoH5CTVlWDaxxIIq52QJ8jIkn
yWpb1PHsdNRkRHwA8gisoLP//4wdLNdvAWaEpcJ3ADs9OPNjpvbFkTm4LSFdv45aahZqUZwthjp9
dMoJKsYy7TGsKhU8KiViEogccYi7Jcm7OLrKoimycopWAzeA36Zcxy6FydoWgoT3ZXWSScdHdqWO
ArFCVNlgG/T6/9pz+uhyaTm8gb2KpMDeMBv5XhgEnoy39my93Ovrv3+Z8bEld4l3sMkr5OTeHwEE
TyU6UozTfGrGq3Z9HoXWBKXju1jMKAZoro6b+V9woxVSFyEkqI1juRuUAV1uh05tZtUddam54HtE
VJjgnAbNor35qtomrgLR5lZZauPgajoYdSsf08/14A+2A0+/MHViCGghXA2Fa7zMWeKZqbI3wLPZ
wKP7POxCQJ4b4OsCxMnGCJm7YnpHGtvHVSDUROXvmpzVKY173H7Cp1F7JpFvB8TVYDhWwONoZppp
Vt1VNn75lYuH9XgS+uqTbCJ5G1iwyHnbYLIK1y5INThA8uJ8HHSWkrKCpU3Wj1p0KEtJSBt1zQ2N
M7GzUPKnuJrX62RqVvldHTD6BmfEUt+tK5JNIGZDqiZsR7IZsmdESmkGVaGRgYkbETY3dZ/BDHUc
b9MdABv520tv1nTiijsNbz5/+5PgY2e9QkeGJgI9fYcuqVwZlQ+nsOjvZdXIazfMKgS7nQMaKVzZ
YMreyZ1BsxgFuNhhf0Jtpl75NWJDWgnZPTfXo4NfmylGtg0mnvNRSW3vz0jAilYtSujbk/MgxhgI
2Ec0ko0T/3+U1IYEJurBac1zZGDevVMbcA0xnPPqc6nhFYPbY2DYfekSeQlkpRbj/wEytSioxwkq
K5uBcNvzrjZSg2csYUnxu0V157aGjHAgGE0b79udWaSwHLoaz2livT8o9YovvCRSzRfHKbA4D+YC
etfNmj7gw65f+flAi/Nsd7XNznyVaOQ3wS8hSWNDLJLW45RedZ6gY9ygQfikv1Vep08zT8BjFRgK
9gIRgXdrrhvXS3lSKDdInZrrOJLBi6huhX9t7F6w2b0I8u3GOoiwle12625dIFGKKMNYZ30ncWQn
BYY6IKWCc9Y69T3Y2PrPW5Ey5WnWtCPmKHFedjtEYWwi3ewuAD3OPUFa+DGRep4IttYoYdE5OWYZ
ZYcqCL6kikjWvNUZZK2Jwl6eguVPBjqaVUFmkFvwtIi5Aa2uqRT5eRc14Lp3fThzywhrmlS2Z1vO
EexxuSagq/cycsh++azU30D2Yi8cM49Y4nVKq/Uo5Um6ouKKqHVa03zRIhjvd1fbF8RW52wFRnma
qEAPQzKY6Dy/Y7nTA+Y3ViaywlF8vCx/waaneCwOPP17/Aj1jgjRXrVc1BfagraFSELG2slKEXgD
V2wqTGv5lXjg/VX5sKx6BHQjT/NUUBZop7X+dVNfO9BOYPiFZj9tniBlOfZne4Lq1AyhHFlKvRUR
EY9ANMOYBoqS5R+/AkySBSJYJzgg3VQyqZ9UUh30bVHNC7iq3Gm63mw3XFYPwzE+8f0k6jAxEJlq
yqKwMEipL29jX9SoJlv4Y3h9M5ZOSwAi95biWZOkdqj3owniV/L7Nvj2gHeICFELT7QiQj+bXNh6
qFvYwE6TuzRXGdQM4+JNDWfMDS7V33FsUmvhP0uQjbexw8vj1mbX/oMUlyW3TLmeyu6Mb/uz09cm
4AeWORUCSxJH4RL9BQ0GtuTns+kE+z9iBZ2FD9o/lnCMLvCCib+JIxopt4e5Ai6CjlL/t0O2CusD
E20X0Pbr4kYWe4CszXivpuZnUMab6a+HAQTpwlkTFkqSg2phE0M8HSEQXZHFQcmoavdLQPmBtQCn
5Tev4SSYGusBiEDoq3gml+k3JS/EcEpfNHZj5kop7CT6gEvLz4neNtg2hiJl8a+y2is7jpdcRPMe
IVAZhyW8A1YtGtNdBmpYoa8zBhgvAG6RHr5NAHSwciWEKmyTPP6EgSZA/73FEt9X7I+k8WQPhA0e
SVhzsb+ughZbsBzwCG6Zd9LSdJ6TZ9gSzFFhTvVB48Gb9gJQnQn+Bz0glka9vyWwIfFQBwR5d1KQ
jMAGAzyposqdD4bCwQOhhqWJVUUTYYc0VWPD/+5eb3aLo/TW7scYcpIgExS5vO7ZkYw256VL1i1L
QwSeApXfW2WN2tDMZjG8wQ/TmFmPAAWCeGQf6SZ7/RjJywH8Hup0IhLzqgDo63ll5H0WpRStJu1H
6fpQ2G8nx5JaR3Haep4hgB8l6iPBZayLT6kQlk7140vW76jxa87a/vTpI7TRyc0M+LrBfBvneGAX
ek5RgV8Grk9/k+qD5hxri9rBJGGmIP4sdWzZ+OkaKB2L4lvIaA5EVFlZWAQwp2fBIhQxnRxI0X0Z
26pBQMu+kb/LH8P6pt77i/emGYswQgKNAi0Kh0+nVUhsNlEQ/vYEy4I5TvF+fs+3e/lFuWMvmrGg
GFDr7r2iVMvu9S2vWAaaFnkAWG+7ktI01NMr/1yHPdgNjWTo1T5APutYe7j5SKaqnX6Ntzz/Dpxc
Y8VSMA5UFxcQyY+QFYxiRcoKYynmEWPcxFvA6NV1+P7TaUzVWauyFeyqRUvelBR31JRYUXBEDIqb
SLTAxLd6nJsKKzfFPk9cuQzXwRDvUvft+afYyNhJWkUtfxi3ZAYaznA2ISLi50d+C5zwpx7ovvkx
q3/RJ4fQBrGwNRBtx680r4vAX6OAwEkc3gDhd2wxdL+XQtSLLsV8L5B6mmXXgSlnJ+Qpj+mUPRBZ
xYUbJtNQNCkcMAvg3VPATqnx/ZI6oz12eitJJwYnUMrsh7TPTSGPQJjJHvqmd8/odA50nztLENIG
FRWHCtl1Rb+vT9lVI+rURXHBsMyor/oSSZg9a3Kx2xTcqwvrOwiCrCS5hXctOFz5zT1CM8lbzEha
D9g7dvA0l0iVnfY3sxYrzuyjNgYw+PEKjhkK3hmwYa1w1jWn5UHg7kFZckJaNJ+kmEWmVSmmxocr
AP9tujHq4U2C2tFKIsVLEE34e5lxRsXM+KG4Xe2Gx0MdEbuVsx9PcdvVnyXusZ49JaNaBeyqaDbK
YyN1F4NG4qXI+J5v2pOrIgn45ne4bO2O9ahxqlTVax1TzEnTKdoeahZ/PpGqmyDOqtkAYknqoB2Y
nByABdyVrdu3RrFMmIGQbNn6WAMCt6iqgDeXwC5YyvjPKZsKvWWNMTAuhtA0SM02KxodAsoNfR1C
t32OZqH4SURGjS+6xlLrWs96uGIOr7JzKlGNIrk2nLDwB0kVTeVeeX+hpmUQZVSKioPdLuMlyVEp
HelxTKzkCieKkrCnO4EUosVD61rGBOMDiRb/E/KoxTweiKDKFuF7T/+IUeLdkwBDiNdHUFTXNpBt
U6j0wDkcexi/DFpr21TjMAqLy+rUj9xYP0XXsUubVU7pkEykOu+pqjj27PcSNhK2BquLampjwAJr
5QUOfNrXmWFpW8YEfxn+xseuhE3kWCINLF+HP8RxwImZedS17xOPk0qP2cAnjk3e3/nFExWlGyD2
0bBMCaSa/4G6xbwJml4lN//v89WzmUlW5XQ2dMVz99YwKsjLlZ7FSJpBglZh44uOlWhsAE5vtElz
QK6ynG6PB0CiYUKVKK31AIqUXEYnaCBqAaq8liQKL40vUra0tafYlAVVpWwWxv+6azBZX4DiMxuv
LcK5krPL8FetW0zSpZupFr43XITWTWjPzAd3lAsqWvf4XhWXHA7PDydb/aNUqFcHaZw3tci7wmTc
gJm2Xs1woJDS7pWda5V0TJ3Ef4BHZBwluZzkEAfwgbxZnav14BTfdKFDyI7Bah5PWCX0Z2LQ551m
arWL4jaB4Ix/QQvhwintqAgx/pOGCNisNqFFrXcqbR3LV2u4suU5+f3HCHmGAtJrqLKAkwBMnF6A
QeO+8tmBeDTcVWsaiyCGBY0HVPp1paXttRm+7tJV9V6IsntQtVv1+gQlDwAHUWxp6zC+qIyNqyE9
pevOOncBWqDnqtzPODewWQHfQrQc6fOHLtFxdVV30VEgmTgGOKKMIuRDpKqlD8TFPenxlF3d0fPF
2uMYIq8p0FvAhiXIPYTQLl8z8DnkQ/0pwtA69rOBlgCRNJdnu5GcQfEgdWBrpiOWSQZpQCENAJ/0
yaERTjwu/iMajK9LvTQqsnIp/tucxjhlBFPYD9TYevtg6ny1XZFdojtxAvgKD39ib8IHndFj2gTi
u17vsJ7XULKHNNzxZS7xWtBYfArHKDZzcskYVniVulRnUrzdbw3T00rDU2N8Kiy2wAyXp48dc8ZH
9v3iSb341026/tAFstez9dWHNwOvcaekQeS8WTf93FRDpt3U4oAYCt2AUh5AreMMA8WuEJ7EoOTY
NbMG2d0oyONGCpUATVV91pCUcPh7AG+Y67ukHXx8VRV4dnfNt+jG4SgNfSiWMrp3Ktnw4MjqdjV0
CYe4Wr0ikVU0jLdXGRmrnXWNFe4jUQGsRO5S5eFJXWhaHVMy8T5COdN27mZbKaTHckHAPgLRKoAn
Pcf2Fa0w2h+wG62FGG8TH05iV9t3h37sKog2fM0upR0Qi9QX4itj+exgVgiyShqsWzYXxOjUfQ0q
AG8el9OCmFwYMTGPRs798DtyQ/gt0PGlAXm658hcg+71yGB/mG8owSqEa1UZfmEngnnquBtTGPil
GS0PYayMD2FOmkuyBuSQA0KVhvl/1aLWW0p9OgG8jiZaOcHvqaaRe+Y7wAnu76Su66XpxuKd9LTf
hv7LUkp+cJ6IwdycUNbG2DBblSNfeJUbOG29HNfJs+OaIQ2wixVfvRU08Axpd93OdPcUuH9OwdBf
Jh889dOSYujBOe97DiFoqoRMeg/pC6FgerXgtiDmkzkeG9+UvtwI9upy85li6y0Qi0cnOUKchIYT
tOfcV6wVP8f6xyJRx5VP7VTLPoBj0V1neVGu2l/LO4ytcwXt+wcPraN/uEiPWIqGTzPhNg8EnVjB
yMfiuPWm178RcfpqfauOBvvgjPcDtIp1GRAnubIvRfZXQ1gkeuGoLmYY3l8Z3AuT3zI6JYEjChWj
4/OI63vhdLuN+UW4zoOpHtxt5m3ST2e+BxBR1yZzb2ooVvuEwpXrtZMmP0e9aB5RUph3has9ljV5
MKE22VRQFQBLtCL8142OAa+VbbAYdoVXCpHauzadccZj/xV74FQbjQYCee3apVEYPkCkMAGvCp0P
p8rC0Y6/hf8/jIZq38eFxV99oA3dNNmH0X2DbvB4ZLwZlTVRTO0Gq7PvlB8YsdToL59laTPaq9ar
QiCqJEiRualSajMXBQyTOy0kImAtMHsDREWf+E2netN9ystB4vzCZUJhRPurbQsQR4ZvmQ3YORxt
fUbQtLOWoTXDZM7WC96GMInALw22fx37Y3UgSyXyuRL2wPnHfb8g7WUoLKW5C5/fYlSSGDr9JAsi
U6bJH5qlhBWnywX3UcvAlLUUCvMJbrDqZTahVK3FPwf905UIFi0+accBtoMc/tEx+W3JAKbaSTGp
3HGzYjamvf+PQebBXVjE4Tk8IGlyaFvHpnwHG3cmWqACfu2uJQ6RLOHeQRMnOe+RQClG1wsT2eUi
8LUwo3moFzsCNj4U/lk6AwuimKrWolXr+q2M/GL2oMU8sYd1S9E4PDsoC75JMPQdp0S5ggHCg5oR
uJhaQCSHrWnL2au4nJ3dVXslkgXrDg3oAFb+CcygifoVWGbtNeUNHSIYW64KUuM7AvDST62qxQS9
Sja4R2jE1YCc0/nz6DYVwySulatmWjZkX+Qh1iqAiywWZ78UVcsr7BbXCOPnRokhHfGKux5suAQk
OwZUjzgUXmBNnaUe1bVztEWn1hdoFP2fI03OLiGNnkTWLIe9uANmVQmdXMFis5Bn2DWkwBPdTfjk
TG90rXL6AWL+gbtHOQaZxGdE/bM9MAcTyUnvA5+xfvUd3Y9K0YoeuZ1VfBisZwHi4YQu2uxIHv3m
DjgY+i0M6ePp6Rh/2becasgHsohgIbtOn8ci8X1dbmJKOyOrORc44U48bLVo1BD45jhOIk/tQ20D
nbBjhC1/Xqvbn0Z9jXTTlTRJwhz4dS2ZW36SvLLaZiwXyluqgL4s5kjaSrOzyEC+bEvaVBJo0+1g
HzWxxkF+wrU0nux69Y+l5mpKOtXeiwim6yMjFPkMq1B9mqEo9HoBfcuWNfanm0rsJVUfVTuB6DWD
mhzJ93rV91fAe/ocxM4O7Zw9P2B7LZdd1FZpXCYtLFYgfaGyF8VD6tWZT97sCb9PkveJcdwEYN9o
+R8b28dIBA1a8G8tSb/lc/RTI5Wjs6+enDNFVoHjEap8qSfgLLcInLefPHb8h4DA7Y/rCwMzb72z
aqYUa5xOKkSK+Oekz524e+9Fg9/xejSMyhwIWS8btrJ1xbuMFX1tabiPv/jeEru2vFPE2NEJL+UX
ua2fyrcOvGBKCEK0ERmRuKShZpPxL6uB/neSAC+TpCWM/jFAwP1swYlrARL7iRiiXoGbdrOps5TM
PWo2n8iWQkHZQhmKWyKeGamp5dzHziU9AicUsl/d7pds73Nn/Lk/eI+gW8ZEMxPS3nVr9Dz0oVYg
KfiTATGEl4UUATF0pEYI8Fq3IDWJ6ESGHzn4G6WsqOrxTJQUuPy7mJ+iqfkaDk7jLPpUQPwgKQsB
f5fEPC2Yd/06jFBecMUifZgi56WqSp6NYU4N4sgI/amY3dUHK7wNyh9k36qgZP4kFX2IYyppFk2q
UmJQjVBFYIDvK7hSqvkYEaH8y4XheJoZ5GXucAIEU0AWkfAeI4DIPSBLEl8H3H9Rz3ZrOSf715dx
pBJfN+3RF2/CHWPv4SvszaouTmp1pKQWfR22mSNlfNgmntKd7SXzIQnN87SeB9ydvag6YM1XzE8b
/JkQAWBf2rRLPl9jjzJAqmvmJnSUbc3xn/7PeBj/RjM9GpSK+DOnPaPuZp89Sqw2sB5pr7wuq28o
I4esuJkxzA/w4COe5qejSGMYanxsFlEW9Utb5lrqSu5QgNmvZwPPgLxXZntVd3qyZ9LWYriYYXGQ
50eEffU/Fl5VSmop1lKi573vHMPZSY+KRnvR0O0BuC7ifJALpwSkXmd2Lfu4rTf2D/stR2xbs9cA
WwTytO47XO0YTHEU3Kh8jMtcUvXYI66XkEke4FZSbwjvAJOkHwoiBQ938/zV/GTEWnm4uYIvj/zo
t609+gWOt4UkX3M2ny0sRManUAhPqLtPN3sPkZ3bysLMmrS0KUwN0UbxWyg1FDq3koiXsj7WvuiX
RjrDAI2QtYzJy2XzrrKZ6e9LIcN4DE9jsWKC9Ju96Mb8xHcnQIc20c7zG5KgSnp4CmuzSFftGNuQ
zRKhoDvMcgfKMHlRtNyfV4ovIcpfnAKBx7TmbmXuVIvOLXXEAwDGucXeNkTgG8yGiGsXZrJgC2V1
2aG2R/RfCuUTolN7cHkC/2wbGt+DXfyEONkO6PTuzqF7bbGVnVF6q7DodMkJaC6R9mqBGaayVvep
YjnmQrrBDJSAjWLBPA1H6j6m2L+jKrBi9FfbsmBiUSWOOxiozSSPbazrp+OoYpZG5URHk9yRg/M9
nFeSk8jTbAX9+dZqBGx26Cg2eJ8BaaS3vwtQlyKMF4FAokbvRd8Eoy6ApvshpPgFaJq71v1Jo72T
vQNyq+NPQEPsZbU/dk8QDGFIrurYuJ/e7CbOVCXNdJRO0U3fOxky139hhxgqbhIDk1Q+uJ5hCsJs
C/vqnNsAhmFGoXIiylYYnPouAymYG/tCPaeiZ6ypAJQSJCjLsspYvThqlQIqq7+IaluiCh/HmgOK
DviOlGb9+401y195eKXp6Q3Fx2VQUC88OWddWV7FqVBIMT56nmZopKfnDbNd8YqFy0kJafTh63pT
jZq8xhS+FEwvJvU9IsOARHFzCbKNuOSq2NsUgeVR5iPiPLHvbz2B53XCffvzuBQxdVOQSBCEHOFU
RoLMySAl0/QJk4ju7GRhs75Aw0S+e0dON1yjAO79oViwNCdBmZpz66nxNX7athFOBoG8HC45YL6S
APHcgBRBG9YCpSQPWmPpEB28ZfAUQiB9oaaer/enVaAqrgQVtBR5PTQBv7UBfPyAA6HfY9l6sQBl
BH8Cbb2xTRfT5ie/J2WcA6rbX3K8mv+MPGbrnW6b61/uTay4iPdGTCCe+NwDjhe0LaOEHHODbFEL
IllummxgKCphMkalvIOLWMhKQ+1ndnyQM4CnOiyOEiFGBymhgKClH+/htPEbhvPmCle1c2bmyCR1
nWDpxaWJJ0/qS5So3Jy4uZ/41KrwJ7Cwt2kqbU3e+Iun5V4eTIykONbyN6XM8F2FRUwhzJqNVqL0
tvL8TIhpKwWNt/XxHcUXrJAiDkWo7X2uebi7w6VHrRx37pleejuiBmcqQqXasYagaongHJ5KkpGT
KaQJ7S8d4y8KYnV4RJv1tdZ+I8KJ6BukWMSHlifKtCHAEJzhJxNq3dR38jPWNK/cZO0Bouqb5gKp
p9Fggg8PiSwXPKIDrPxjEBFABMrh4lnYuR/t0whgms4bDs7nlMBF/dcLAWUHhzPBEYuz5xDjkrK0
mAsZ5XAtCzXX8ld11vO+wwnYfvtR63Abs3yKe2vMu6PHuRS+y5mWwko+Picu3P55ZJ/2XHmmbo/y
+slgdP6iptUtFOZzkFb9LBrtk369rmToN4AovIZrtHWD+FeMPWUlfiNHmfkBvQZChmT6bum/ekvl
V7Vhobte3rNFdJ7K/mjr7RZW3X04pJvablx7WFgIEcFfSJ4OP2mmn9cuzl2xBazvFa+MXajd9iNR
Ef5hseEn2cZ46zq6KoeTM6Su/Va+7vmcg/5LnXbHgCKmowhPya11pMAve4l8Bf9XKDGcJetpRYRJ
6fPgbHNO4c54ldL+s6OF9fGSCpm7YUJD4jQoo14Xp0g6ScGLfXM9/mwwOG3N6VFS+dY37nP3M1pT
IhvNAS6Rn+FiZDRkwri0cbR8TMBP0yudpMauEcepnzD2sC9zBnKvoLC8WmnqYFtYt2pdetSEdtrV
q9PxzWj4H1oSMnIJpYH8Qa0dgkHWwgkTMDXa+G1sSx74zldvcj+ci+et2MR3JRofB/xePKuE/WMv
7n8eMKdORPZS7vtuGTgUCfMai/cz2UPQzIxwxfgikasDam8wEwTsplB1+O6STkkBNLRnWCcT4Mrz
xtslbPlDO4aAMDII23dKjOcBhH+8FkTp6rpZlnRa3+mVpIfIVS10oXwZ5rwTlags5ctMT+jcKFtj
53VCLiWJ4jfW2x0OTjzsONIEkJsXRpgySPUxi5Mpx8o9885QHVG3fJEK6C7rAtG9udITUvrkwp13
hmrrE56urOKGAIqBbiSDHRqrwnPZhwCqBDZe6kbgHOABxlM+AfAV42R/MA10fF4L/Ec620xubx7m
86YvZMMoOOvRAuRDibTM7BLsVzuosMgWUkakvVngMDCC8cN57r2haSWf2ys8qoWKBnhvUYWPH+Ax
bYWaWA6puuLZRDo/zrbErpzyuuCeDuZyT5nwoPHiUbSMqs+H9XomeXcyrHTAgeRnjVSlVWA83upU
ALJFRllWUxh2X+63BRnEXpH+2nYiY7pBxTJh0slUyKD8d2A49ExgOC9WCiie+28T0xhoA3NgATDN
JldeaFbQFZcmyQ3mwLPk5ZDwhloYMdgAx2ts2HEQJiTYDseuiO4H5Gy04LS1PZqnK+Pi6nsj5R0/
xXotzwDg2413U1JDxFn9V2wFq0ezzQaldgpoL+BqvnQfnx509thVS+R/AqtnNXmk22MJcsqU9SR1
/+BqGRdSETs/D+5AYzSz9ANWAsKCEc0yXWTstX6plOVhJLwe4CebJTqwR4lS/AjE5h5sr7Ub+wca
p3bZGyMox3PSWIpnfGYAMylmISbPnnCIjbLCy+1bpdZQq+nTcue1/3Rx3lhFn34vLYQm8hBVambZ
VyWw3t8Rprvxfdzj0l+TJ5yx9pobxWRTMhkJ+62VcG88l6OfVUlBOUgyuJ6nuqfKznnKJQMp384y
jtfcTTlkY/FtzD0ediT3yGUZbjdJiUyvMIWltV9auMjMgfw/EtVRMFPUErFZoeo/z/W8l23xvWm1
2XUmi5u439cl+7ZDrVpoEAO9Pqnf5ER20eoRgUbPdvJLEbR3/2d2LRGDYYjpGJKPEGfzqsFCjg3N
zRd6maNhD0KFdTphYf1LoTEbJr63D5sZ2WLwI4xMMlVgkh6KSU4xiMz+jMh3mwbZDomCkEsG1DtL
Xw5fpP1kj+VWSnvHiXJpGojYECZAkYwCvX880EwVWtQPyTlqgOWtkPMwI8mHM+hl8rk/lUnA+Xdm
Cj46lwdrv6AhByVsTILLPA/iCO/8mcQXdHDLKsp4vcxDEpBjAjSNqnhJpLVTtuK/pJlpc7AH6kow
dJ1EoLFYAcodD79Oq2UuZs333y5VmtDw1rAbFQ0GJAHM9irR5GhslLU+z3WdG/XxEszyPnb5qBu9
lnL7guo3SANX9x+//HUmkTzsi10QgNR/2sRBXs8TDl1Z4OJdBaP5yvIRSegXANVYtoWQTB46wSsL
34i9rLIbp4Ywf7J0/cMYQNjLgcNeR5W9/D/l/gH+vzEdDdh7DurOdX0y620Gpnd77Jm1CFRjPQBj
fk/9mBgE3kqkHgJcZS5XgjEMMn226gaf0cz7r3vfZEHNpbJHmCWzUTBoWSiF+LyJbfJeJjVNTCS/
kVmCtMUyQpEmqoPkpqbrNqWuhYSUCwEZBmDWpQwiQtW2B7C3REvEXNjms4OsduGZroyEM2zpnIEg
zuv/58jvvjScwkQE8Inu/FS7rMT32Kxp7WD3UqpxyT+IhoZP3BnExHPHhmYbViKAnqSaspFa+a2H
1lGyDlFFUe9k8FFjfqeCXcJ/e6zppjqaTNY0YyNPlQRSrDIXYD10LoPHEiIQZLRQLjBzyrzKzouL
PufnOK/pGfFLzeVaG6AdN2ElDxw2a/QYz4F08fdh/lHTpUaTUB39Wa4u6cZP1cy49jvzhXpcOdTT
d7Lf3a50eP4QCA+ugxzazPcYEMir9qt63xADWWQyuieVzvOknhJ2GRPGNmYhtBVJjdECQgwUzBq7
Yp+30yZsABVeWeIFBAno+N9G00iRxmFd2JCFcKg8GkdEzBox8cgRaDZ6HTBMEhFnP+P65rAIpfDP
p7ZoclZ9CAkaQQ70OxEeZG8VNvnOTB42/jZois44NyRN8vytA+Rq0oAoklCK1A8iJZwuuSZvMcgJ
X+98l1iVp/5kZt1D6Df2Qih0Cshxik0GfjAhMGr1Jh4bzfsVJ9J1MD9WYQtxI9020Kiv/zhaN4X8
MQjHUL95JlHO3QR7rVfqrMqHGvW+sA4yP0IBaXfZafL9abSM7kVs4WPugionhseudzp52ALU0Oup
6n0QLZjjZhRpUsYdOtWX+joOQ4+1m3GPCvFCz6pPx4YTEq+xMHm8989Q4bOs4v4hEI0fT4Qr9PgJ
IUkQQHIhtHwi4LTbz5ra185bI1Rzkv/TpdQc2T+M1uBk0gi+TjPdoijKyhHaCyIa25es+Ggr3Z6+
yyQfE15WQTCOvXF2Qr7dlsfOhmogQGHwEwmhZKy8xjjXob9APbclR1Yp5UC1pl32qwF7HSuCRznx
+4wajUdivPy2GHvAMuZaWRIRewrVJFQe/NtRxfmqDmgbfvyPMO+OjgN/Qm8PdGZxuc2qPjCtAYU4
Wi1okDBE5SRcPWa/e8DWmAKVlKrkVA3k6jgywVOCJuo0cloikpRNogM5kHu7y7viHGehoTiorRbn
wi3j4UbnOmTIXW4yUE9gpQraICZFY/WEHrtwkYfg9ofn9Nkks5xLtAcURch2aQ0HE1HU0I8FQm28
LROx2svnLt5GkYjodD4xbpAlDhltU8hDtywLQLdbbNKSakSEMIob0u4zn0oQt4Y165Zol76gF4cz
k08xdXDqqvbnDCzsl7aatJoXoMUG2FJ1edBv0/dI8R+kI4C9YrZD0UDH7tJRXG/HXagU/aUAfd7I
49I+usxIeMcDHxwxfsYy9YU2Z4jIaxxVgePcJRbKFs97z+7Xf1jXgk7bI8W6fuKpSYKySJP1wXfd
xEQqzLVcVc8t8K04LtbVnBH+Sg1f4rkN6Ghu9b/aNS6sdgDtCF0m9DHOZ4Kd1yaKkKUwnj5NdbK8
unJcWFrwtAxcnI7mhjhvhYRdgC0das8h6zixqwbvngAJ2e0NwoPe9GY6kLVQGNmdUJeaScwEA2B3
7F0qA2lVmT34ppIVAS04k/P0xM8dw5BzQrbdq+UzXl0H8FqEkaiw/Vcp11mnVJAxyO/jyOhrfrFU
Bw7jlcYF/KKI9vL3GJgi/W0HZzq+SYyySFgTPdy8n0Qd4EdcdS8E18ZyoLoUOmN6/AiTL7V24nua
eEmZVyiq05QJ3fx9SA2HFm+Oq0b2ssQx2ShkdtDpKUEVMkLwB9lkbpyg6o/6bkQ5ZfjL0rnoT2KR
Ry5xsM4GJppi7b+HD9Ed6efJCqZRfTRXSVKfWySJ/zuMMcaj+AW4i0DVJYGp4WpFW9CT/D9NDDit
XhCr93CJmvhsTlZ4VURKuHkidgw9htf0Sblxo3v9l3rGnNwh5NxaIUb8oWc/HBrTqo7ZtwTdvmwx
aDxyEoPXe3VqxiPC1eekCNH1GY3b3yRswGvTCyHcqAndrGZtKsnEVnaPN3h1w49QRS654ak8jsky
ijfPEURYyEGH15rKnjzbUGSKDJJstSs192oyrlBmxG/2LAVpdgjwlHKjlNacEtghTZxDobFR+i8e
e+Mj5O+/x3u5hyaBPqOZsYDFnvbQtVgO4Nl72Z3Lu9bC7g2CDLKponoH1ziE9iQCOkznQg0RZsRM
q9ofXVFVHoAbDpjThRceUYbFc5d34RkO9MmMetOcCOAAwH4Cy1d1TJfce1Ae5pAABwoLRyUhaHEB
kC4r4wp5hB1C49qb2iViFs6j6Re0hDx7/6iDWZ6EnBugPRdCXY0ZniApdZylXttmdY1lND663Qr/
rDYrbekOMr6pI5RZt3KIwsN1iurVl8ur9bNbtjQ1x+FsoLd7Slw9ZxaoIk85CVHMpgWcUBbUcyqG
l3oSlge/CzPAG2ssAqTXwjmiXyQWHyujP2h7Nm3STe4SQeFvUatkpBdn46eihW1vW7IkkfUfazc2
zB+baPsO2+H5QweC+TeI8QvrU0hoJ4J67kznGjYtWQKajw9cEFpLqqo/43A0R7xukv2DIsEOabeu
shD1aM64ZOU2MP7e1BOh8iUKKWC9bcGZslKGi8ZV1ltgITLlLVArwOngPeM0HKeA06penkIfa0TJ
qbNymlTu9XX5LDlZ97SQDJs2kLTVSYzCAn5BdVSFrqBR4lf3HIb0urVmecGuBAB04dzFErJGSYOF
5ykAvJ3meFsl+SVYO5DylGE1/kbFhB7HtzEVbhYBwLIkz88a/cO8mwmJflspkvs33oThlOSnB5Cp
kHzdsBWmzJ4z37/QmtViuRAQBdiu330ccc7/8sZTgXjd7/3j9qIMWj86wKTo6xgECMusvrgcK0vV
hT5dveLOT361Gvyr0N19QOa8jpWmmeNW1N4whfRUA4MmV+60SNCM2LtfINFKh3aZHVkYWXT7f61F
2MexdXubUwWawYZLk9tbHhzkAWckYFEFy5cPgdJ7J1mDjbxSYaZNNkF+f39XQdYzesKgggMK41zC
eIbIVNVhYiD1tiptgRwgkHXrzCa4iaLoCDSzMzjm2XAB/Uw1zsMUBcNrXiF5jQllxO58tnIFuzcg
j9Eak1NZwfG/RJzNwiVMF9YFgFE3aQmYZLRL9OxQ/u65trzmjK6zZeQDfcOFXQxZmb+5VkpU3Gap
AYrtFjupDI3dp4ZE9SQ68SljGPtrony/otXucG1ZuWvC3n9qXLsYLE7SXSFzkC+9WbtVnD67zhys
Q4wkcocfduq66uTUZe+FBRQ/J/WDaBHTYPbqz41AjQZPmUbPjj3mJC7QXS7jFankaBn4A7ba8koH
rifsDKkpCIdPCb2qJpHUbKHEUyWBz8nxES09MqJ/XxvzZMbWn/BzW0H4NnI1EIw0IikHfF7apvZC
W4U2i5MsmymIO99vMa+Om16cyqD5sVm1ncFy6+FUgh2T08ysHIuxInO/l12KrCzyvMr4PfucTXw6
ny2Ua1Cosc4dkIn/h6azQ7Q3GfWSvCK4hvQGur9GfzvvFx0nQOhGLn83aLKd2ZdKzRGNr/W4BBC2
HMZ5zo2a7Pi63WeLesMYR78wpKi+inE/+3FCgEt7Gkn8J/UOVyZ7vvnoUqpFmhyt6wUzqSA51ZUk
eIEV7FJVsjJ7iS5qzGQjsjhQ/PZqAKRRBO4NTpRP8b0Dj8RDLgyX9oj+vI8B8dYQmU4HJGImI+V8
Vpru/YG8JJRJL1s4J90VT36z4GXcJ6jL0f4mBEOxoGVuXOqKYz7+L6whIgjfxSwEShw7ecLXZyt6
GGcGSUvjwdhyxaGJx6aE/DgcjayIcmzuU5VXLU6X0EPDDKMJvU1uMAsyqzpoeaDxVLHBxuPBhrs1
BXHVak6RCQ6NISGIYPFDJxeSXigWyvchh+kKx1bfn4woP3rlhs97c9zk4FX6YCHTcoZ0Kq6HWXq7
wg364dsPWnhp+RySpwrPy0cCe7q6sveWIrkftqcKkY4CSezuglWSc5S4Mju0w3bx2IL1k31As9F2
tHSpIt9QPxinyGGJ5oPmSnM4GPe9CbuCu/8QFnutQzBXPnGoE3zJvUFj76BUCvChkRbFTHyw5IVG
7RVi8FLI+dUbQSYp8y2QJeNO81tUsh0fVyMhbYI0QRCgDL3qfLMSwIpj0gDOUNhcpREHebEQsssr
l6hm0Z8VwX1lzXGPgFE/811Qyy6HU/w77SPvHXxU+DMr+6axoxR583lvTLd6UHkuxF8sIUs5lRtw
gN1+RpChE71rcwsjQg6VyKmxVX8YV6BI1C/CfP1qq+fiASl2BsR2eSudVSwCX+pJsGW50rGGrTOy
SHwjqS3WgheJOXriIDqwq9hmMMe4gCiEMiyh6Oyb/t2Xt2vYLPLtk2tcOXr/UQkurIA0+z/Z04JW
d5+toWP0S2VQLJzTLdOEHO69WXWIs6iRJNPMmGgx6atwW9NpmkCZEYqdWe5QyveiwuekXxeHyhYu
T1r526TqkOcDngGpPhySsMAaA553QP2rAa8pR1YPrnz4j5D1G/K49zou4vE59c70dH1xJSlf3VmH
3aF/QTbg0f6Hr3JdURRG9ZT+nwcrmKNxmcuU3Zew7vgjXPlOGcnCgBPXeD8SrHUxZLAHA4TJgVwy
7Tgy4p+x2rOu0mXbizifbbEit4X4sHBtvwt452bShL/hWAEl7xq2u4rs5iTMNnalXjZDc8dl3HEC
QHNFKYOxmsoKIZW3p5lxsQLFpzg7McQkwnDrj8OTcMorcWjGSwg1oNBjyc6jO+93GLGGLNJvucI8
dpq/smXPoM2V6uH0stWOWjABdEQBwdPuhPgcw6R2RpwYGwrGVsG08MRL/5vKc9N7MZKZsUXTEwJ/
xZwu61b4x30zfNCusufSP5NC2n/nwfX4ECIxO5VUuhP1+t6C6b2qNWjBbmhq2TqkDMscDe+vQdl6
44KHnhEJhYgyUomI6BqLZRnShgBnZahMN8baAaMx/3Y/SSM9bpzseSWoAZQ2oFF6vAfsrARuG5P3
VCOEuF7i9nR9p6Ej+jwPM/sdXvi0LxfKbE4XEBs5C+lRWE7LkFr5++7Tl2F7nMWUSZ+dOPZZNDrl
t0bR4ywcKOY1y1ug+CzpBEvoHhOvJqSNrJ3I9Mtp+x1ALUsTFvUqQ1iguOK5zZiNed56kwWbCA24
J+dFCpk7L6two4M70sAO8S6qR1cGCxvU02Cim2R7RMONFpUws8tkPA448glBDrDfPaoyPWYu3h3D
wDZEcEvvOoSShjmNyAvI9lo+AYUcMlVJUngjGkZmODUTcbBixQIJ4RihFcaTImuPq91xcR8ckopU
Yv11yAUDSD55Xq5N1RAW29EriSJcxfI5Vxlr/3Qng2a2MYpGhtWe5x3jIo2/HS41OET3FM2DJkg7
6kgmIA635iACJp1oy6grNIrx5GdZ+OI/3ZSAM2bLrpasnPi3vK15HIYpmv6ZOJQEEhLkB+Klw7Mo
wFyv3OO8xlPjgF2WNVNgSHTg/tkYuC405/9aFy9NOvRFI/NWMuEf4XLtteUQ4RHCM4XD+I0VF/xq
fZsCJALR7qXP8WlUI60OBIMNledWtjU1yc/t35sMYWqQfL/hwbJs+FwHDNEnsI1JBM1SzMT0YJkv
4HJoSNHqt/YRTHxhrZaBYNZ1bmfJvttA2wkqZtB3BeN1/10VSEUlrFM019nG0ImPxr7esYlAjVC8
Y+zclxtWVRfPQhG0BfcxblYNIThloC0XPI1ek8ETNfggiIyO3rgrET0o1TPC0VLwnhPwaAWwo0YB
ybLsWhMcMyaWBlkRSDSrV1DAYZq5Q0DZ8Xba7IYK64VZAsRvSVIW7Jxodp85WyCAK9ElS58e0a4B
l0BId2G6rlRkZinWaZ2FEQutn3Xhi3g4BVWXmPwXXZ0dtJF8UGIHVp/U7Ih4v7C3TkSoHrLieS5c
y2ifGiuKAhzWqpCqNq/iVyiBg3Cw4lyFSvylnePToPQ77bgEuMDA3uAhN3LuAdW7dENkUMKOmdXn
QgGwlZrX+59Dh841QIqdduawsIzYaJCQToFzVQp+FDKk6Ok0unqHTOFLkxTnPJVvlL7zCrAH2WCR
Hp964RpaKdvkBTp+z0PCX52XPqtNr3HGFNmJnm1xl7zVTPVnW0SIRkYHtWga57x8yrW0BpN40qhY
sdqq4mfurQR+G/dQUPAinLLiL+eNMPRErNgQ0Pro0ZUQIfAnH+CC5CwKr+Q9n+7i1nEq0vjDDmn6
UJ2uBhoQMhrvvBl8eQvxaCNs/pCsgSXGz0sckyicTap5L3Fg4sqsgPYEA8RW9X9cUyGd5TJujtDp
5uI6nw5v67MZuitpZ85hGz2n1BbYm4pkOMYukHMNLLj2SUkWk94A4URYggZtN5mHizHkYXn46Kzk
nuRzMqSFAmzcKdt1xdBVRmOX8jCu5h80JhEwig9piCNY+bpNAGFKlZbv6s3VNIf1xLGMZpR/8QAB
oD+HhsisqFJB+N0QxnnShVkGcE5drwG270SkxJfCerSNTRSeQxTB6B+PYahG6dqNjOl7UdJIasv4
TZRUGHv2kq4bEIIDQ9ODmpxGOl1+wjLtBa8REbWavxQCiuh0ioyISSuQd90HqfjtaJ0pvZ5XAFTb
cvWZK6tDmAHn+3hSHqlwOYTrwF5Tklcz8KT2zHRWFPfpa8l1M3cJ9L6g0tO9Erub9Kt6W0Afi64k
RIRlEl+u2zuObb0SMdjiG7bqAoizAPXahemjzU9Bbji7jhZCoqP84QrFQQw0hkkiOwt11YIjtPYC
+gqKrdnlul+cc4XeB/qLQhvgQbJqYO64zDDAXYy0r1N0HtaB7y6CaQazPLGK13XtI/4gf4e/F+V7
AFWvHQTIB/2szoR4CJ6F8T8P9gtOfjMuy7BOfh6UO1KQ0urjtcPzVEPlNiCnYKD9hNX9Qq/hebS9
9NmhYbLHSdBQRXAMjcpClpv8IXfN6KNbHM3tJOpDja8R0WsLeRUXnhbrKEaS1ZlRbuqsUl/yQF/B
JT4CYchenMI/dDAkoiZ62YPNZ7MGkZQlXJW/kMYL+/d5Vh+tgm1ht2PQOcyY8NbNsv7yw0gzJkxk
lARsl+ZViIR3KWdzTC2WdsqD9GcVc2NPlxEZgJ+TnM/Xycbp1kyhgzsgROSTzk0D9gYUi8CqP1We
hUBictx047FaxsTYdotOhCZojeHzGJDqMX2Q7Zgy7MBDuIV2JVixCu69CQVw3ORrbCB7/gPnmDKw
f2BgwvrO6zx7WhbQPSAvu1xKh7oJORm41RV57VHr8eJoq+RcJjjQwthR/OOwAlL5mW9uJoKfSfaa
Oxpn+PzUqSADD6Kh4UfTugjrP9Ehltj8kzB7+ELyAJ5fQ1R9FxbSdBKlXPtBGJbEnUI0UjQXfguZ
eGq8ggcvnt16gOTIYY/vwhFqqNKGmaSdty7h/HIvDkpHePWE2n9cPBVwXs4ykjGDeM6Z0Po5JPVM
NwQNL2e6eKiteLLnusNnn/DUCCdV/GhkfKkn9j1A9jJXPEJMAA/OPkWSLpoh5H5BV5uRK+LL57rD
mhYXWOuOFTCxFjvoyefQ3othOFQk/RY7/DPojntRf4YsdeciPmLjRGqyGnSsz+jVpipEK0SgAa4H
K++OeVEAuQ4SJPaArVb1w8uHrUJ4ODzhej1I1GOV1QGL0AICSVgW5qQ4OjudASOFHoAhb0aeSbFO
stnAqom2GeecdFDO2UY+o3Nfkg0eZkT0jXt1dolmb2K2yld5Uvc0oiZaYIpakbE2lAd3T/gKCQw6
OQPBNSIJLpqHirwgECD/jDvIyETBUL6uZVvmWoBwtNfQA+8mIDlRk1DWHFJOWsmf7gGegeOJEbe+
ch1TVOofKZbNnyZqkHv9PN7vTTbsIQTBN4DDDbF55hej5raNVWcJCkPga8EoeXYHQMrhUvJrCkLU
IBTnmvrolyEZ3TmTSCJNOo82liQ3pSCdidkhzXxm4QTYI+B3Mu2/8R25KJsygWL2ViBzJK1ZmqSz
pCZ531+iZw4fXs0FyZLgSgPPiYTEOPivbmS8U1txrDf4UnbC/R88GltLkX8dDeCzcjveaL5ivmUC
8HIpjI7nJH/pcX5UuQgWwffesEZNGWZLm8Mel3rDStMkUZGBrwo9UXp7ryNKbnn6HuSP0MkQ3elx
umbgY3x45hHn5I12LT1/W6DcrkH9mOM/G+MvGuYTBwIjsLpIcvK2qsv04KwK6upqhXDFonS/0PUl
1Iuiz0EujyrAE0U1K45ygcE8PF9LkBAkDXTeArW7o0Db6JTWjougvQPVqOhG3CKtZmp53ZMOHC9p
8StFF87YoLJimtoi1g+Q8esWlJIh7trShPu390eA7gP07ljY1uwSnG+d1pGK+yzupU8hvjgtwmtk
+Q1li2L3c0BlpO63504oeFYKsaY1fjH4IFnuOqNgVEIOzSlZvUgCyKZ2Q599+n0xRBFvR86Y3cVt
Ufgh1mXy+f9mOhICcXowxhu1TuYjc0HWXiasQFFuA/+WoZ5HtxYP0MP7sIynjHxQHGswiLEVeNR4
NjLAjaqKmXyZYWe4UDpBVtnaVbjaTZOt+gJ2Yu4yewMt6pcB08eETJ43vHg8KtGefxkkZn/u8Inb
D0iJoGXBcfWnFrLTQT63i1MVgv1qx0ZKJiO2262m6wYsa7NQcaPjGfAcfugQqOOUuixv7uoBkSn0
vTqvI83iI7pBYV1ExnwdCO5eIoXzA81+vrrwXip5qHCxaXvQLUrskCum4tY7RGnf3784Q8TRp8KK
epZqGrNHTPqBiqKhtwwjbTKYrGOLiUl2N3pjJfCIg1p50ZVfotGKQShfA4dR3fvx/CjMH3V2oQcK
C0Evr+NC3qFyV0ql3hJHa4khfejLrCXnZgim93ikW6O5eiCTvU3SwbWl0ZRJb+OLHfzP/fcERFz4
LG1bF9hyQhmWnG17MD+Jc6KMjsOqsc3N60bX9bKl+TbJhyyoXq9VWwr5mj9fK+9Ry/AhSpjduAlC
xNR7QDOxWnNh2+4yUeyA31qP9ECezyFuL0qLA52WUBz44MZ6JI7v2GfrbaW0oVilLOxyDJPm5yjx
OWJy2LMXjbEqDhxE1eNZjkkGSVq9dOObC0/7aA1uv1EKc5zSPDosVUWjaZQF5gMxT0v6SUgFeibp
mnBly63zycSKXSbVB6BcGfy9MrFsbZJIz76dACXpjTbrx1M6zvT711V5a2R6nkgWXE5oVAE2u+VB
/QuRXiAFiZti95afRkHpukeW5suOZqcGcZsyKKi2nkPqKprBwKXovupxtwhfcubLWzU5BUKcyOXT
W6LTnl5Bfve4eAcfASU1oPb0J30VJWSogO1tn0a9DAOAEeSfoeJpvVOgGulrvPiTcmo0eQSn2+Hy
qXbma1D4fUrrJ/8ZWqLnEOzJPYkySueXAWaNmPIah2Cz+vMfvSHeF89maWOeFSen/VRHdT/dNo2J
iCV4isJQvI1M3ncxJIQHt/4XWu0PkvpEzGwlwgDTIWYV77+4E1R06S/q7uPfKtNBuMGN2ehFVYnF
GaLPXi07MYQQU5CxHt82ncd/gOaThhfWlbDsbwkRgmDFvsbUEvDYiKieh3TdD7ILvza6k3lXnvS0
ORpDGT5knOlTF1zFJwJLH2ISoP2L95jJmSTilIpBnm5I0qJ0VUhH/xyqrMghpCCT7/9nHhovBUzy
IDVkT5wQ+fbQOPKCXBthQU0qpuyydwBuU8zDk/i+kdjS/rJOvkM/7no74lGXoNImaftOZ2Y/LypU
Fx/dRZl0x0nlmJLOxpMGrabrVhkySVKix1Z/I17HARy0UQ4Hk+CTUQ9XpB3pAirtkqxtzGqvRfgn
2ehYtSQ1ypixfZ+MhNFGVAVBhmkUbfD5a4gmPiVkYCB9NEWOy4uhP8rrEXhp8nJumKzcZeIJlpff
gHEmPpRT1/G7Og/7udG9uOuu6BydH+KQeOQAfZh4CO4uLiTR13aDdbvi8tIc9Xt/deeC7oRlWEyg
gwXr3uLcCUPTLwezAbpqxRI18R+OPHfCYMDaKGR8bxv5zOAFC9URNzFUNLXVYUuB/B8TTqJqDrW2
MYSHuGRVcC4lis8UNVE0ekWbX+0oaeZ83jV2WtDqJn9q/DHG1jve7oiO6PkYNikXQ8phx9nF48WJ
D/BdFFIvBJPMMH/ahdN+ffuTcl5oNSHM2jSO64h8MdvFGlQUFSM85JAblYZwZhoCjvTotUOxQTyO
jTSfsmFFwI8As5jjOW8IMUld7qnr8O5g58AAKIuWgO9h8h0Ikq/V6FY7ivL+V4SWYEsHruYqR6S4
vsfAeCMnVdJsVEjWtcd8quNvlYaWDNBaIaxivRhe19l1sI48Sufx2a8sRPOpkYAZPslg2BtC5QcQ
hNnJNMoR7nh5OvgVKd9XIECkZB/XlL2B6w7i+PzJXS+EpFz8b5o/5kIDOEN6n2AEXNAalSEfUlkj
HKfcmAg2mz/qICZyZ+jmSiY1DtsJfoLh+xJ13ODegO6EyJ1qu5pOGeLM+dBjvVKwubZ7IYU3c6K0
95uOHnYWgoBm3I6m3+9Grxhh1xyfn9sVv/rKCklMsoYhXzNjoSBfSXUdaOAFYzpls+XQptLAyyMt
qlkLbY1NMPWCWLKal1Tkqqc7qMkU+ISpUJu2eWSoBBPYsubq621cqUK2ukO6QX3Zz/7RnEstF0Y3
NgxvN0rvUnaxtAbrlka37pqX5eXpYTJS07EBVmx3/dQj9zau+x/HAZo0vaFojnNcgkmsollh43Zk
RDuQxy+BpQPAFyCshHR3qVsOcQbWjhpmntkVIFCb8yqlNJyqynVv8OxCx9tg4hcilAjnHWDX9M7p
98IzEB6gLCyMIOptMfBtJM5nwR6iyxdLn9u4sIYIc778ZiWQeolVsJbSjxjyVsBmJ11VruSLUb3s
0QGn1ESXohvVffCc1qLZWNcPSrj/zINy0BJyOWGcDiv7vFdAEb5EOtCWMviK+NkFxGfX+oelB0gK
D/Kgc92JUUWqDDFRV4Au1QX1cfTMISRt96DnZvKQTINmBpPj509j5OHJZNouKmAdxQnKGxglZAWy
ifmXnAxmD0u8ZYI3o2mHseSEkXeLXSCO8R7dFnt9YL2o2zuQqCjvWWQLi8mKz+ISWObYLxFJnUYq
V0LDvc8a8deBuwp+GWCscToEtYs9+3E0KSlXDA6SrR08xVNN9/5pqbZOdmS4mS9KVIpGYHe2hze9
Tk7FIqyowS2cQ2EyNO9/p09Y1DdLGFF0x2V+aFusqBPnTjgwDNlrZrSgP90D5axlHSZhSE4ABzcg
5vZStMnTsi7lPJmKcYTqpu8X2TF84Oq9GaqMU7SWe39cdbEIvhD78X7QlQ57jibJVpALsiBQb0Iu
6mSuTTSoJ/hnIxtbO8Ph3lg8oteHnOAq9CCmk0OiNveao5brL6QaKVsARJrwQ4v6OUeWGd5I0PUv
REbaSPjqqBxOs5wvIaDiZ4zrqp+09zpEK6tqwpC0bM6qAzlR+GTDlaDHnjaPlGB3pgdBKId1Jq7u
pi5VxI7XL0XQF6cS/bE39+k9rAN9rJOiV1WG8ewhafhfCqKernCmEQoPtzPAYJResB6rCcsk2InG
lT75KFr8BQKrOpF1iOMy9YGHWKZ8KVh56J2tJ8qKa97FcUfpl3jVcOygXFQ6dhCP7g/ILVdY/4Mt
3C79ynJ3WR84ciKG0L0UpPXwLc7aF2rw/7TvIhl2Rlsi2cXsqLP+X7F0tQXfm8uFl0gjjA5P+LB3
ycEC/OITO2acmMEdDHkzLNSYihUGTFpHsvHyLHL8Fw4SEQa5kT/55YnMuNzHjqD59DAdVxq0S4LU
nsqrujCwr5BbCmiVfUGuXhFhDu5NcYXlRPdnZaGEfLjwIIqXXL2qeeC4bYBlXer5egrE2eq5CMER
nYiplvHQamziXuxg3Yhz5a4jgfp4wcsysgx5XUwrv7rmkArG5s6/IHPk5d7OHfRP8FTxX3czU/U2
3lblPNMRy37T4C3VsgMpfENNkvLu3SketNoWUZ+pZz0WgCwEcjeTiAMgMlnMVKial2wh9ESqeRQX
f5rI+H9vh8OegJnd58fmlz7aGa1TqYqY0Efp58mQ41E138fOydUVq5vo8URVPWV9he63VOkhJlLp
LaRrsZQ+EPzX9qukJonOTZ/Xqr6/0Vv1flflE0Rzu6E6RzrFZcqCxEecUat0Ix3waYt04LTXfzM3
PvchBiqfeZXHJZMyzNGSA6HvnOMX3/6Gn7DFY4f5wVDGvmP26Qmp8YE7wFR/JfOduCT/9ySGs38e
7qocz1Ay8OWzdM/NfULr8gI234+RB9sRJikk6lJ95616ZW+Hf9N1bciGELpcclvQcAgqNg2t66Nb
Q8Wvs99kKS/67w89EGy3rAC7ZzzQ26iE+PS/o1BDFv4KfbvPXxFiOCcSxkCggDMxzw7YxvFlSBTA
JE546B0hOVeLwIgO4ztsaKGnOF8x9uJMZ9EnWXAcwj4XuzPDUn6v2Em3y/EnE7gg61ujeyrXxbBF
0rkL+yOe/IRyF92w8A7lvRhvVU4nRW7Na8zZ0ctEcpg4a42HUQ/5M35YWztAWXhDZF83sACypxE4
7WmBPGYmYd6t8t6PVGwO9/a/cvsBK4hXlMf6EYVNvMBlB8DhJx+BlLmI4WcD5eQ2jCA1rtES5KCS
Imj/1QvrDnuG++tG1JPAQMaQFa/gECANRxzUVL5DFYpGY48KMEIXqVUANHHJ3wYFJ8ROai557CE9
PIM0nZaa5VNLSykojiY6GD4y2bDmSAUBjEDu7Jrmo+6+0XN95PpRTlhUfJCMjVRCQZdZDc3pLz2P
mWI8NOPXBEZAbKPUYl0Zrf95VsR6KNO0MotsYyLTJzv7BrCl4KHAvAcG1+dTnlqNPever8GhoEZv
f1tuNLCUyDGu1VULE1Ob+hft0u9QCzn1zFz3rhkg6Zkc8DNpFNzVpn2Uan4JqDkU1UqGA9TFEM3I
7bPzuaqXgG+ENvqIm9HN2CI2SdK1chMbqZjlpvelljXk514oUguzyj+B31HPX3g/33IGsaAqeOEn
RO7iT4yHTOWu91+Zt8OrMIwL0IfJMkusISO6OvuwUia8seydOMZqcr9v6ov6HwgnMYmlHmLUPbee
6/sBHV9Hxoz5VqbPIIc8XmW4tvpDGQCiHjofru/t+Uzw8vkzrogonco3beVb5w/RDLvhZ16NTltB
4J5H5Kbn2L8vOCQHCPvZVx1vND554DKOs8JLRLFwPxpMvUuXcHIOyoh91aj9NcofjIkQdU/j07pG
lQvD2BNy8ycU9uBTJhEwit9f6BvDFVDc/Jl7+QBxATt4fYYB+sjbF7c4my4HWE4vzFj+tnEv+piw
6k4LjFoJN9+7PWRxpScXR8P8+QTkUd7dJwoYCSTu/uHOhLNnXAzTXxwOGycQD8sbLzOMLgjotCfA
hCnh7LmOZYbtsPysFPElEh6rEWNVeIe0XQx49DnYLZfvNEuLpmuPVZ4b7ydvp3Wi/D4t8qQ8/ysD
3PYUR+iqHYWNJqALoK75yn7wosD7aiBZbuo3F7yZzSiIGz2Aqhc7vZhQspeibdPbaiQ7LOeVszd2
xJH/chplKj8lFkZYKXExb50UfDS/ARFLERWmSnWog1VnXXtdj52e0/vK+fYNt4500SEeNskqqnFF
RI01mNbse1R3/iXehE8nX0gNxH+TrkcNI9dCx7PAYTbKu5K7ci6nDR0iJ4hySqHQ/t3GlZFmmNHI
994iu0vcShGsDsQ12abGYHL6hXh7f2nlUDxYudyUgJOAxfflkjkqL/tqnwWrBkpLxwISZcw4m0dS
Z2CMz4KV+vGBlVxAudPjTd7QeLoOgyAhmzUY65lK+8296DugMpAL6jQt+16eow2UwA3LBz7hmYOn
vHwjGTD88ngWOb8RU2lP8b2lM4Fs5Ddro86r1fIqXrAi4FFH6h227tgqYkRmwzowjCJlSayIFEOh
wBs5OP6KbNQhDEFH4WWyaVFpPrRxJkTm4SJ6bYsan394SDDYzIEordTCTcKAjsTmzVtxifkLnfaf
KLPpcw/Zaz1bBVvqbkvVkKHHrcTsxJcPd8LRJgyISVEyk5XcDoqlat2gsvDgGEV48VcS6nA9Jpf/
eihyyngNTT2Dt+ooIWtdCzsuioGhBK0GS3gyGj7vPqikFQV8Zm8nUvgeif1z6eMYJ98VWrYf/ptX
0jw0OIItBoZ2yEJPJ91SaHmqqAsYUN8i1PT82U7CFJY951vi5zsOp1jE/XGrmEl+ZJmtZHekqfXE
cEJALhwjpeH+PnNR6NQykdVRORsoWjLM2NZTCat+yhWwKGFErzGBWpvgBl4sw0EyhW/p9KcuKlgq
/btBLMiwy9/SGxj6Qnp048B6SP5Byyd4y8TachEI4q11RJgyDn4vBM80x77DTAIgWLzjMfkNJI/0
ciy5Bp2aPLTsrAe5pJRAmvxpe0CNA0AHeGJbpj1oactFOTpA7EEQVa0wNyR0i0OwRzJ/nVdQvQWV
FJLNC/m1iIcEOOnC8ilT8Ebh5OgMAVmFWhAJOd5D9Wzpi7oQl3yDEsVr5QRVWbFPKetgtmukrvBx
PDw7K+8XTFL+Ri7qQf0MYageTX92+kBnUqQxD2DzoCfHITpkQGG9Hy02PFE+WuNNdRXQmmfY5tGl
U+yZNzs0+LqgaU7sO/kSUE7lHGU3j8soY1yNE6/H/pR1sUeyrPMhWmTLlTZ+itoOIs6UwoNMKSR6
eerwJE6FZrmkYJ4DiB2vMO+5rNaRBX7Kbio9yIqI9wDcc1a7KZhYLADsWjPKsED5b3wOas2EWuN3
bjBfjH53SBuJX3jLxeo/Pv4+revFsXlLvTb4u9ycoinfwOiR93CvX9KoHcuC7J0byDtIffdFjTR/
NWxn4JeRIZtAGdRP6Jb5AsKTseYZC1R40j+EEIiBowybn+yxy3Bu0NbL6stmu8+Gam9/65A9ghPu
I1NW1Xe86258qso2d1kMIFtjp1Kv4tqQ1CxhGmw9v/CSYybD1V2/2imSJiPOomieU0mSIVybSjhp
iOWeMqylloV7O/oyhqv/CD0con6WtCy330TdahxtrDmKd5JwWtPUFJWgQAsR16Czaozf0t+XANaZ
qIkrWjR4KrSZgJ8bMtdXPrOK6VdzLlNNUBu2qCHVWXOU9M52/luAa2MItN1O7rQVOfIibB0wUtPN
GfFxl4F3N0bZCYs8vAJGh9uw1oaJhL44rxKyNzL0rF7ELzM2nnFnaUfrazYrfk2BSMLBa21E3ELh
rBGA5U6wID8TRLpngYYazwofvEmaDpllZNG1HEgdSeGNYMa6Znp+0j8UlW/w6aFRb3Z7pT1CO3FQ
ruq8j4iDk/bZAGUIDbjnLVopge/71WbJ8M8lRHPZVSES1Z+Az6r+GnaEQPOD6eqCjm1b6WVq+39A
aJvLui1oEfrD5Cx/fYCcxPFQD84bvVtduYaK1VyJcjHYzoSnea5hmuFSjMaOb4qVGkeNswxBkxCx
rcKpqKIQlN6VFGzA8ow1FFBhFkvsdfs29i0Iv0m0HGrX64Oe81qjMplyGsv9d4w3iT1jjaqSSZbQ
ee5xg5vUx6kl8jgwQZsNUeeHY9+V9byBuP3wk9DK5jYEHhHV+KE+NdH65BlYrgKcsaVTIikEvq5J
WCS2kjGn+wR88wL6L8Cr4ryg0RQEJ/B43IJ08FUegHaRYQs6Y67IBLYymRdzFf+7IhUYMAB2WFlQ
0LQAp9JGizy79zGXFfgybAH9tdRzFcUt7+QzfF4T9nlGLu3bMIN6N//vz+rLkD+1SRrnRAii/i/3
f3pagDic2r3hJqEqfsiPF+cW7K27EKYQVrUuzyYnTG8XAL8el4QfunY1BtX0WMTT47RuhMs1S2gD
nKNIikVCXguxa1N5evAd4iQL2khIk3RnEQYnnfYES6p8qh0ngtmUd5zc2pGIXBZLRoOaPlaUzHce
be6FdiaVJ/jmzblww3VA4b1Ux58/I5PQdfsxvXCKiG6UcUBk61HrEGocstLscYnGqpKfDBfZ5RfG
PzI5y8cjEH6niJQlfEDp7EHaSZKGDPbHfb8tMHpgSrVTZD1h9xHihyGZuOFPeHq6qadWFLd8R2gP
FCKBz9d/5ZVM3XkQmbgJ9JWQK9AZNhPuEPuzRcXr0+eOQnyzXVQ8nhjLZ1Dg0wilOOWrEWBKKGvp
cxZAqUMYirsgYOJE/YI7MDy/gv2E7aGWOIds1nOsUK2UNv+PzeoyajX0xiwU0dFjsyjzJph4FN86
jot9jceiNXGYFqQLn/1TbtU3EloCNXi4Yf3Ka9trmx7NG+5jynFPOjh0MckEIKOryyFpOvWjBGtp
cZzLKMAmN+XpcorVAmXq7ze0FPm8spZH3+15s4UnMNeVZMRFgazL/Vajqtai0bsvZpuh+ULDs2Q5
SL5WTBworrC7XJrGFq2XRMfnL8fhckdV3GIS4Uy875E31xV4BuZB63wphN3gdRbXhSlLGkiz9UpZ
NN/pyAtH2pPDF+C2cWbRgef3/sCqU7tx8DmhUhwGba7Gmtvlrw7camHLvvj7iEMzWUnpDQIbDhJ4
MPFQIUsXutb3gmiP2MFAYjGwYtP5jHubPz/VPar08170rSDI1GHW3JwHcTgN2wMJ7Fk4g0KsIg5s
s37D3WZbiu/Ah8JyBwr62IK8I1IcE4hmRxXfgh/bHx8NBvJDcIaU398zfoxTjWzf0d1wtHsS6+sI
iAmFOHQQmsQOi4HRcAU+opl/VQNc5NT6h+RhBupugz+TbZf0YJh1MHQJVfRFx49GyzNSHyQf7Wz9
wtei29P5VgfTCFcBp6SVbHXLhOhU/nFMb0xROutxdL7LRbvBx2KZc4IDIDd14yUHAaHa5KL+EGxT
hZ3Tv22WbaSqJcJr4netX7Q4+4DkCxQI8NT2EXt89OqDUO6+mpciL4QTMIEjbx0wdp+hc2A3/YC5
ttwhLNQHReEwoLzlSaTaHR3hBES2DoU2DhN6IaRMRPorBH2cjAmtRRNsQ8nKeue+gR+xlrBeM5nd
6/6sBlGlTdRx66kBIfSszLceo4Mw2K8065HmiBn+5X5szjvByDlfP+pqGXAK+9zkLuonJklGwpQ8
ojH9qlfL8C5/43fMhI2zVatSDReWGfeV+SrzBMIs2exvQvbKPCZZBcE+kpbjG4Y2O+g1XWJfDFAm
nrSEmQIyUeOrvy0umQiF4GWkTkHxHTb3wzWyJJhi+9BQ63oVE9h2ccmM8eJSGu4kb7i/HMJExS9y
dWhe3CqOsng1mRQfDh11f60yYErQcN/ve6GTE/jA8DUanzO8mYsAQHvBDxOXNuOVaSD4iYqoC5RZ
vVxNzU0qKTF64fcNV/4PVZL2NuTEg8eoX1hYVVyA8xx4U8OrkyzKz1ciHUUvEnKHD+8FRNUteZZR
6pPIXGbcEJ3UYV/5PzhmSrmv3WSjNv94b1bQADa+u2n+u9eBn90sJ6eMu/2y5+PQGz7uV7nY/ikq
YZbVuomkoOUdK7ozQ5ZXl8Nykdaa7b/uKmxF1IPk4xyCNbIVPSP6F3g3Rn9taFprGsFS875NACKd
omoyxSNztbb7fq5+8+Ih6SA7aKGOxoqtC4TyqXYZaL8a8T1PwZGjLlK1N8Nv4LlOTBtDfmXctfxK
LWQNmILKjBDd6UnwTSYX51AMhxqVqN1lWcWYingtz+4pIbGhW9S41COQ7NCdBNnoecTztmIlenTF
aJTuaenhYZdwjrwROTS0C3uesgfY5/NG2WIssDRfNbQxZPl1QZitrCK/UTchL8NH1tmfLmv1lymk
stu+OeeyzN/UxOMOfd0ju2HVO5YyS0Hwyoy+QAQIADdOhONAcpHUbL5Hqm4FdI0J0DuZ30mbO2zT
VHmeIUPWCzpNs6eoA//i8tualDQBqAHDQuOJS4tLYckgWt4/NwhMOmiuB9ph8Lxoj5hBhUZ5ZnFB
1fBPONbumOvMPY680aUAexlyyfrQVphpJ1y7EU80DV/1PAXQLhrn6LDn/MgToJuiyZOAXvpi2CU9
hxuEfpQeWznd3K62yJmRgVmiu3ofok1/nVc4ziz5h2Hj6hBOc2g53/RE1whyLRFIN1zQiwf9X3F6
7LkGigSdFGoZnlCl0AXP9HwrJ0v8CeY8S+ic+XZOqf6tzVpn4yO0eX4M9lgVkHjQ5yrRtYEWjtZ8
wbie4r7u9HC7N7q6iO4s5BXiwLEeiCREzQwjwByJjLTizdpTyZpZ3x5oPtWA5ySq5EVuQzBxWPF3
8cy9vMHYkP0LzrhRy2vq5VC/DMsprIplt2mEMKDUhXTnt362LGoVtd1kqnYtT/yt43LxfTi8Kd/1
iOF40LsLeEEK/W77DT976z093AHMe0NRqTkaX8jMNMoPZau8H5YKlLB4v+F/FqXaqQyfBj/W/Ihc
m3HghtZLioc28WfDbHb5JP+/f2AwncUaUlGAQYH0zhnuNF7cJ/0Oz7k820U+YUSWKNN2zkHPiyWy
JH4lSrj5hUqwA6fzRcIfPCX710w/r8EY/hApfa202XFDtQnnq2lePY1YzuPGSPK8nlVJbJvPF9SK
xVV0xUUPwjPmwip1wBAy4Tfxt/YPg/GkWwfapRzAx6dm7K/6mcEIKxkEb5FXf5A5SCHe8f/9cAoL
PZ46kiEh0904lZfXV+IAg7kGX3/DZxwJYUBcW+bwBd3gGaT9cshGYssvG0u2KT75uevSSHBJoJ3w
k0z7DNICGpxv4gH5OW6V9sf6BxKMTKY9H5ykTHsDwXsoT8WfyXcsOqbot84raeStXl4qr6DPZ6sP
FnGi88vFT1mi2gPl+cPHWy4vIVrsBWe/97+9SyS7+fBkoOpofxv1qA83SeLRbfrqILddQMJ7IZhg
0Yw1FUZzEaSdRy2J6+hiY7iutJ6sCBAzYfpLXy2U71KxGn68GBt+yy9CjBsA5Glf5gEQJKo5q3t1
BwcmkBZ5/l+Fn4OfQmlFU2QQehGNRdfwI1Gc40b5OFh9lW0Vi+tcN6TcE2wMwrhU+Vmcy9jUNl+B
duAmG5SQ6yz6EA6zCIuJ6s1yIQqIW5r5uIxPV54UvDuoHOuUzw8N1VnGmbcWatzhLghKI9QTzFmu
JosHGW169kFdH7GWZx8UGfY3KA9LKiZLnBAk7mKqz3uSEhag/Km+6ynimi+4o4rS1WKrNVWrG+Wc
u9uGWjFbjeDS+Xz06Raw06xBXfIeZdI5rFah+jleuJHsMcjA8HM8bwmLFuo25udPQMGLoN+UYlrd
+Ys7EcaTw3Ypo0oFzZq1iVVy7GxGkKCYM/ulu/rX+s2qSP/S25OnU3aD7wcbTfRv9f6egeXnj8Et
ST8NMZHc+L81rnvWCV5sZlo5dinKE1xRTHUK6OXHggvypStRKdZ8Q+QgHUFxLSa3T+xh4NIcAHy4
f59deWU8qJboWYEY1PnLimZLsYDvE7GJhr1Git2lwPoHBzoOV4FKJyH57hvr+ke15RvIW1gnSFFR
hVWsqNp33453Y0XVoYVDoiJ7xvinRdQWjMt1CR+MKGw5y5smWc8wa3668JyJ47axFMZgPxWr4P2R
9JM+jCqohoziEiFXn0HE7yzdc4DAYxjg0ZmJqfbMOKjR8Cs5EYhLeUJvPg+XBwH3eFzJ7KjySmFP
kamxwB3JIlc4265YyyxEmpTdKtuK8h72MKvJgKWHKE+OwncWZ297yoG7A0mstq6dwycssgbmtn7d
xA87Ue87m58BVnMagfkoncIO57607KT74orh8qv5jrO1cO/GWLp6LqxEYChP0Nj725k9Z1QoeSNI
6nVdyqdu/4sCZXUOJBjQCmHU6Pe++Ts6D6PVFIOmR9Rf8VwzhyqB3i3yEJ0H/OZLbVhhMpxch+8e
MF1MNMWF9THhcnP9MJv5vQ+U/M1ZoZuIIcS4oRRBunzIX4/PMEFIs1SleLgK9JAAd3xebeqWbUB3
IiNKuuE1DhKG4/JUzFvd0qhV8RDgXR9wzzi/bXnuu018ng2QeH5+4K9RS3Xr6GAYXtFTudm2x0ME
zhBsV8kEXnQGHFpfg0ZJ41OxbDI5iyQLPFLJdH9FLuy0g9ZyQDhsAEqlDIHyGRwq62nyH8Wr2hXf
vS0rtgQuEXPNmI1qITinPWhzVw8p4DT24OQ22s91J26LcVNVwExhstYu0xlrw95N4DkW2u+XrZhe
esO8Se/lynNS+zvG+a4BYEm/Sx+3G6CfnLB2Lczbw0MiE9MBYRfjQHfgPgf48il0MnwFOOEPCrEW
5bF6q8/s3pFVn5wptD9yefvMdZKcD+bltHU0pVuyiV0o7vKdYZnrx8ZrKp78ay74L73Tp8xCAnq3
pHYxGiNy5/xFAyCrnWZUjNtgw6ALkUf8HIEIXJKKD3wtGTDjSQbkmY+7QQVoxkyso+MoZ6sJIUXV
kTImhdYUwNtq4IsSkmatULrVQyvEOl8T7Zx24PYNDeD73pm/5rN1k0NNv6qhEIW8NaD4vdDlzsHU
MpDHEtRILpmhveJ1M8dktz87Ik2onRQLu4AmZLjeWcox0PbkP9iqMBd4thCI7YQtpyUxZfpPo8a/
rTXT/6hN6qWcsRBa36thbbbP/IlkdXP4nT9I5PFEjBMKFd88c5ZTDdYZXuBIZnnLyZIKqEEsLDOc
X9TZPd3wRQsyqtknupSTrPwiZfmy9bbBHs9hbjtVuwRHc3emm021l/SFSsOxHUxQtrD8YMtQKhuq
+Oz0Bw28kuf+166hkr1dM68kK5uT7xFMrlsnXgvK7psIlXx3QN0XZ4wk9QMTdXAZENG9+GqNX87R
u00m2nwHgyxgQXzR7hpWWJ1kL/hWfe+c4p224PBirvxm3BD+HW5qb7ahKUDaIVtH26lXq9YPw0fa
LO02O/LJCoI/w95pHjdZNRHOKjLtSdoHfxWAWm5ybXY+VyvIAVD2FzWN/w9JI/9zPkCOkXmz/m0u
yrwRDXW+SYpr2B1kILQuVoqcOiClt305lWYSr6NTTCqy7k69EjU/bYjZfOh5JoQAhmtiAddfg19Y
/8Z87pAIjrXuNkX8QOALthL8PEjujb1Y9tdLVs+YW0ur1xvQ4Iw7/aB3EMneWY8VQm3mZ7NRB5IN
xuutusw0vL0V7Yht58GqwwiL7aoP0STH/6LIjRh7CmhRu4l4q//uDin+z/uo6q3ipj5YuuhADyc4
c3GmE4v5USjdTlolAJLgT98t+smbCv0rWcwfNh+5yiC8dODWrorgmIh/Z2koFsBVlTtzcHWcLR/7
4nzO4ibuzAKmfO/e1+asnv1vSXyPlwrgC8p/p+GTmi9ZyXw/l8pPPuIAZv7xHYPVZvC3Ivjn80QO
kkLIye3xA4WRk/7zY6Y9IXmZz7noI6zemlFev5XNIBAyION0LAdMDbgQyORW0iEr+Gd7p5U0ZCrr
KOHe8dMuiBcR/lp8QoudqzhYypekkd0/uWAO8VS/O0W5GKwIKEUHxGSeLS112Mbi6FZkaxjSA7DO
nDycBWC0gsrfWIs+B/IDwNxWpgc/qYOn9JmZNtDVkrQAiAq32Z5PBC+YVaJ5+cdRe7UcASII9jxm
PsK6swM5n8dnbwzhdTj/i7eAjKIHWkiuRaxV2EH4Eo9Y35B03gfY1eRtN4/sJAsov2iOae3NcJET
F/PMZzx+v9Y33b+uO4Bvg00dhd+aickB8L7CXXtjjJtiNtF1PfAs6hCTrRzjwlHnUFCIUkpnrGqB
ZV7j45PizEgRVnsr28If+x4LT+6xeyFIHG8P4elH071YSYlUGrEH3nf6QL7a8Nt1VHAvuBHsRM4X
RucBzl9YLf8rWPLkFWoTMeURH9mdyO4dkWi3WotZouXcBQsvAncru9ofLt0nKNwxx/PaxplcrTxB
2o3AeJL7l6xTYTotrwtj6x3PoI2AvUrvvERPr8IDwOZGqgUybzF89jne5Z3efuL5fwEE4Xo0maPW
XSjEfV38CF0AMSQbUqizk4RnMu9wqIXl5UCksS/fvITdj654SEv4lWqlIEgib80pryph6are5qBo
Pu2+qvwbUKmQ6X3wQamCveIQwuBmk3+lkHmFCQcXJ1aaZTbs6eJgMzAaRAQrbq+4Zg5DoY5WUvG3
PsGdFP8REQWVtBi6IE1Rp9VLdFk2JReAtjfKfVet7guemsli75m9L8RWnw5PHvDzrRB5Y0vW1bwd
jDmM+DzJszBP0GDzULyeYHw8dUwCbSiPqowM8mBlQUpYQosohqH4dRsFlqoDRPZBsdHOrboATpdL
2ggoye1HIWLlUltTIWYMfoAfRddy7g2duRynHBEsvN/3y9NUOdRbeIDSjpHHDE6/24g3mP9n/EOY
79WTZyzdsAt8jFv6Bt3dyURz7daxYxR1IPoJseTmM8wHTGwMfsystN7cACQVYZTXOlLc7DhfUvYl
TQFZHN108f1XBCXgJ3hGBvcJfvhALHZPWxs/QIDqr5iDFf7gvH2d3+fEJcNUZ/arI/xbM+ZqVSfc
2ZXhKUOJMpkUIgBtlp/5EUgBj7f+OvbdodnkoDeqXmg+WI7uGoAWPW8MzS/8y7qPWeH3uhkDSxE4
x+BrpKabQZYoTOP7VrwpZleBZ6bLNaNN8Z+p6k3QDQF8Gb47PwulrMCKHAswIePRUYJYAnIYDCWk
f+bSUJAqDS3z0daHjCHqpIJKBh2rznZjdue+SWCN6d2GPF1fygsEt2guLMye3lBRQSp+AYcU7gq6
QbNYqG0+Nh1DeK0fk3jfZmHFvXsoCOTnfz9+XJ6GINXuqEEaNDiIQE1vbW63c7OmRyH9Pj0t4qz5
Zj8DkaoXCIeCjr0X+p7EH478DM1PPeyW/bo4kY2DJvcMTVW8DqtdglSLvR5x7zDljXSq19FbcF84
5Xm9vHoJusp3csmREE6eOh7fz0yygQpxLrF8jhT+eowkY5hgdaDAx+URpIvU0EWdzaTh7FIKtq+i
i/9B6NyIaphC4XCvObf3xAx8DpH2/wdbQCqOUDYiz059icCsi2iiRVYZd+oarky3FnF4QaHcYmi7
S1KsKxtFDkq86142sl3NcVIdfTvR4klY9sDai9miN9ZAlDxOoJUVWorw3dvDSFCRj9JLo6q+JX/h
sFUj+xI0ywOSZqKmze3xJcqjgjniS3yQrdMNlQMqfUTMxZHR0Tbie6GIjZOiMjCPY+/nU+h5HbVh
90bvcTbigPTJzmwAF42rfBt9ybBBUM1a3MeZsVodcUgfU9yipQRFQYl6u4h1poPLLjFibnkiMBZ0
PbghciqttYNFO2DIgMfxYiGSpASa2+3YlwoVMOSG/mNqdZVdqzE30oLFcHd4uIzg3ErVdVWGNK68
rLNsh1c8QTNFYpGsaIYBE2hkdhEeIa/rj13pWQq04AgsQ2GaqOapdnZrU2fK8KuQMXXgyZGgD2xf
fbXDJ580XxtfC8vKBnC1vj317DLpnFomXmE6oPchSzRQD+nKr3zsaYE8CA4qzX3d6/epdRDc7nbB
xNhMkcyFIm5LYduxwLJVPEcj9CtfC0HQiZ6vkGrvUsl0MAbDBB55OkvWKSdkWA1ubCRLDJN5P787
itJ3BYCHa1LGPM4f33/U7op1nAcGkZsmGNAa015Ug/MQzX7AK4quYl1Mx0pELdiSoHYnC+Dd3UMN
HLF/IUPBZ6tQUU7mFZ12ddaqLSdiBGiS/R5hyIyaZpCzp1d7MJcNpsowOdUDaCf7rd8zVUutOWhz
zQDnF+4iSpln6HLAmlk0xeUiKv7CXZ1JqeXOb72MWbRY+JlZaI+Cd/6NewiAIq+JVUxo8iwzn4rE
UXJkApp2s2H+4d7m7xKvv3kVOTupdkLaucUA75Tw6XxMp58mATfEggedMa0rK93apvP7rZS65u5e
rdZ/Mf4Au4zPXZG2GNVJGYxncXhCR+AB8RHqkiYV/nB7mUdAcD1ApWr03tyjjUNBSezkpKVspE3U
gHFrXTGcoRauKHyQodLtqAG0H5YV9eRQV7Xt/ZxK9oj3wBBk+Armrp5+VBFBdVhTVzUj6RtKEGKb
zR1JolEyx9n2xV55WrtDIerIYBKA52Q0cbwPY8mZ20J7zZ6DtPPxn+BpcLNTVbiIc8Y2lmQ+V8j8
qGweS1DGfirpl1D0Fbditv2iu7z21RnZWGN24tyDJnR0JYoxeI8aNN5GccRErxQX4Zwj8Dbe7EJR
Lz3GpJA9WTKQQtsutW/QvoGGfIN7MaT5ZhKz+RxU4Tdv1qoKa5T0J4EbAz2xcgIAL+aeBH+eEEim
Nm2cRM/6LhCT68daXtz8vMe2/3QPtLGRRH3LO3RZVWyODjrrx1L+p7qjpNWvKvTSbBtREr45oKoS
BxVmN0Qwul9S/hL+dVBp/IhOYPS/jdXtFF8P9yIcxj9hCXR0HEMK1lIrNIh4sfiuj5kxG3N9lTOv
r1rxiqVi74aycntuZWOv1QkNdYxAtn8a6xTOCqyxM1WKN5V7ukBvepYnigyHzRwT2o9UPXZIzj84
K5LoFuvHgJPUJW4No6idjt3w3pXrAuny6l18ac0TJG9+pMz+YOSFyutvD0xCnqsc16E0O6LeVgNa
PpZIBFLhjeX6n+LBYoOUB5qLyWwH/Bn5JDWUYvRndpechEn2lRWHJW2YZfSGfuRLeiLZdvNuTiiz
evIj+/0Bcnnq/SwLCRCk4Nbjmzy+mVvGg+UGhqYyhdQl8r5daIPdu3WVCil/d+YcZt3l4kW09BWV
pz0FGyukYhO3xNKwoaDicha9sS1TyMLjWibkv8akUUiErhcgR2wAajSTC8x9stUJnEVQsGp2opTL
asGDsUHqPFuZ50IhEzj9w8UTPx79JzrJGPAbBZYz9bdfRIe1KtuldFBK85BAOYfHE7Tvnhp2JtDG
148zzCU1+2EreHXtR+I3YMJOYdXJuTuGaFMMTzHoJo+KTlXRu2s6snQY/3i1+ZB/k3GF2NOL7aY3
+sGmmZgHcc++GyYwrxgS+wA9/d/rPtbypLLvRPq1UJ9NolLBOlNOQ2Ivscq1E6gYac3XNdb/b9Qh
OdSYWtP++k23KWvivvlJRRI4j2KYBv2qb9QmIYvX6GnhasAwH1nj4lkeCjLf0d0/tKwcLflBYCTo
NRWwnOT0uG/hyaES4HnWvjstIkdiR7gyBvIaRPB0MgMLvL2IvMZ8OnxkFJw051OrEGUW2ib5ddve
jgbD2DnjY8xJTkfRz7TCSkOLsSqM5TfwCNciViM2P92ZW67Bwquq6AuNiyXC3NPX/VxNK9zQjLY3
a8Hy+RPlsTPlDEsltlV81lvXTcRYtSXi8MUnZmKgwG/g29J+IMLrptwXzhXQbQGccLFXpuzBBIQS
YZHZSHz7qUMeuFmaQUrQGAND2ZZncamTR3FVa64nnDy2p0yKf2qzRQ8yJfvbrEisn9aMyMldtxFN
i0Jv/oF4qRDVZkhOOOjCFoqjJ6vsK2Eg7lik9qmV2qfa2WNVmAA9CssE9xm+seEaLu8vBBKH4ten
khE/kuZC9fR2yrU8EgDguq6q4hlq58LrJXAR+N7N6FAUdX4d0Er6qNdnzyCqTz994KoETzWQsXRR
wEGrAwHvM4XxFw4erMwEPfD/nMhFbc6HZTdr6GqBtZAH4Oy+hlIOd495Cme0c50g0/8BId1DVMsn
oZG+DY2afF91Vgw3KrcVK4+yz95z/J4wFgsm7VqVkPHP6q1qu7mcfF54rmA/TiwOKmKQZfmrlr96
yt65Ldp5/5DTp4DD7nUERi7EedmGhUbqUKC8dSqUdSAYzv69Q+LI3PgcUWIqd55aLErgEKDmyPPE
Gc5DPQi1gdxeAr8kZ+VHypxr2BEHJVCKswWwNWSrx7GlWysYmZ5yhidDxhxtLKglEdqG+Vg7qQ6j
zuMuVd+xUCKCPMdpUzHeEHXXxAbyqH+xghbIlFXMDDonK+Td/qUg02dlyni9wkFwAW9f3KDDw4Ts
c9POsNWy7FrAZ2JsnaOyCiV44vIim+diCOR6BLCmyvt/mCePqLvIWaCEsuQgsrEJCPccVOTsFUnw
an/AbUgb1ARlxL1csT02vsnj8rkE1FryrQlVLCG0HkXW+xK+07BZjAkpPgvtc8N/m2TJFBnx4Kw2
0STbPethaJUBf6jsMxSRJ6kHhi9r5rTtNmS1Kx/6OU6voI7k2zcU6nvphOpd1peepv9IQ8jlJAaL
XufV8CKuWLmZTy3CK+bUan29nQf5LaoopQLfbvrX++/m/orMDRBwE5nhPEde9rlFsNz+zDLak6BW
drRSf+F6L1vc+erVO7U4tb/+p/ZLvyUs3Kns6OoAnBFlp4Va2LtLiEjxhHWa2sailhwR9uoWGIZt
elTPE1U8vkaoWjsYAM2FRvfIADiSgNzQMWrFfFoUWmi5Qr3EIghzMaqLYY4g7NZlTsF7Ww52SoOM
weH4j0xitIQB1iJ5H+gfJlpaTZLhvKrnQg6nDlsMZca0YpZntQbolLu270z2o7TF/6p217NwnooN
1RltWNn6n6g0EvkloeOBqm4RkW/FHxKGQSPrUwf/mrUmyossnSURz/0J2HRm4NWiWs6IWBbTB7nN
yuCUNxh5TczwvzhfLAXH8z1Dpos5ZJsGode571eH0Xt7XB+gr1KU6MlbdWHOLfh04a/pBCAQ/6Ga
R9n2G1eU9FYAmxva1qefy5T56IHbhyGEP9XPQOvEB0LbqnwMuMlkWSNgbJO9vaR4qqmL21+xpmnl
1Kxhb4IHmb8vIChq5AJkmlfULFJJmge6FUv+v3Qbu4/3rcTKqO/ORoo4lgUlfdDKRKXw8w/+5Mx+
8tahFq7WF9o6DFaqx4eLwf7JRTyYwnKi905yhXe0bWW8po/tTqvcgHCgTLIQR+dlxbuKIOJidJ1A
vAqs0Ut7rRZDmGv7w4WKtG0BerJgDB8gmM6nEkfAh47hfveYdKNuBZ7LzdTIy6ycBDQoXbtmH1Pf
sF6Yayk23f3xQzOiCNpDYoI0jhHzcUQqJxlnOG8Xob68pIB3358EgBHiLF2sJbe2SRgf713lbcaO
8pngoyTNOsAWqtgcnqMPdufT5+yEeTJQpjzmSbIZLsvIfvLuCCIM3g6yhrGtdTyiaYQ4KFbw71a+
SLZ2rTSlvHQvoSkwQQl9if0jBuC+PQA8Dqjg/GvFfw/MhbGtFcMLFIOjFQ2LU7YM+sIzmWrlXUoE
tK1QOvkcf/Nu1BXvoKzZLFJTZ3VfRxvpLCg4L1N6M0GQCnOxeGaJz+BHa1Ipemq9rPzWYjDy23ug
GfV4XeMte9Gc+jzLgBMbaxvE5/E7EUfA8b3pZr7eLyONwkiW1ZTNOx7m3t8Omd+ypkHVOMkjHOx6
dgx4Kq7CeV+/K6jDgLdUihBvicjYjlPOMIJKeUwjUaBViBu0bpYw7t3M42+SOpJ5KVGkQm989F2Q
5xIXCJVhU608LV9Bk3LrWW/zak88MKfIwgQHMftPSHR3zvKpQrKT1BvgEeIzx6v7xmgwgBJVi/hc
Y2EXkY+0tpr1lv2e8A42y46R+7xyTnmnwPejldnd2HuRh/ul/rq0ZdrsINl5ovvKm6rvwGtdm4/E
Xu3eCa/aiR6mAWmxfKsYB0db8f2xrwYkV/fctcvkcv2tp/T1/4SmvYxIfrmxxNKPuA2Yz936Z/y4
8/yEhTR0aX0vvd/NrszT7LOXeEt1m+IqF4HbTyxhUjf7ojO5xW+24Iu5MeDGPnezv/lnULjarSs9
zhBElZ8sHoQw4AdqSDMW/a04djzLE1jnf7KxpQHcptirBkWn2ElRexkDLDq/+9zJKnsHLEwV35rq
vxz8jUjzJ4zI5DClzKQHJbaUZZV3pOVTkZag84xVUyFc1Yye52NxNTaTE2gomUorazZXc/oElXC4
D13sZU3JGHyNGjTUV0SW7sRCUJYbCRTv2x8kFerBNh2S3LkzS6yjAkqhH0nn0li/Yks/uCVaHYDe
OM0oR1B0HiuN6nVdqJKzRKu9z+NO1manGqcNWAwKBgkw7loCMDekt3VJL+Kn7rRWQaQjq1uH12HK
stQUSr1+asmNlsEyXrKMNxw/kesKqQGPPrcPYSZtXdf1/PAjxpBk3xABvlnxssSRqoCbFWfUbfPz
R1j8UZv24NdbeIjeom0eVr+y5ctWW+Kd7S9Ss0b3MufuO+oKnz8wXrYQUOYOs9uatzYW3p53sjVT
RFQHVAelqRfRyH6S9rU7o2STydeEeDqBVBoo/e6VoS6jAEHdCNhiUExLNRL9a6LYjtHnmaumZ9pc
6VG0jzTG/3lGxmSGH70GPhbvME0AqLqSs1n7DehtAlsvTomONiYfhYepGrFa5pmdYXNcQP6A5HS6
yQm+g/HiwpLZ8BApbSarjZ1JbaYGTbhVKwX2xR+akT/3O+K9QQyoJMq1cmvYsW/iJ1tBZSxlgmeu
4FEgnBaYkJZfAPcHrDJt6aVjDpZ2p0I8eVqBHRNB4InEPZUfoirFCOn+3ny359T6+A7IVgPR6h8+
n5x8O8y4zN8Ov84HzaezHOgf51Z9wU4A8QLbpKOcMmK0kh5qm+9YruUGa8GlcO73HcPfBt9lXuGA
5hGrijqET0TPeykzxgSG6OvrTA6e2AmpjvLwFLil/Tdj9rPS8u6c2MO8PDp2gw9fxSgktvexJlFS
an7w2UWkYGKbk5bjysdtTZmHVLKUTeorJWxf1+gcllAV3wZ7hM9DNoAWBVyKVjFLJ1jHRlMZyK2M
iJNso3RN5eYkc1JF1awrsPUZOkZZ0rpuV0PpQ4D/qDs1nt0iXJOmDNMCxOMyiVZE9Ze53TEbiS7t
r6PhV2gZASzYWTzMFmpp/6W6cKqcchbuJdBn5ELQVlBhpTFBwLuB9O4OlO5V/9OKqQWr/mMSu34s
+D//xnXRm8c+BKXyLEUbijZHaMBydnUTmaItNRLYH5h8Jj1SWkfht9g1nydL8I2H4jYWbnY6ZvF2
IucZwyEPoTA/nJVfONDHpY+oInliobf79hj9UZRFPXHAt15eDbRC9fP3n5OmD6wzGt2YKAZo72nS
j6HFFFY52r8cWjio0+93KBjfQNaGRnVXAyRikhEu1NbaaCMcH5nvJFMmOh26rUfi1OfzFwYS5CW2
CdLQ6o2rWd6wpdMX/PcbbjvuIz1mYNrFZhC19/3qd95Eh+ZWR6ayCpKMpPRmigtC6iZqra6pc8k0
xTzr/hICAc1Nnv54G9cSnOqjWJ7pvhKpx5sI60Nb26jjv8ByvybVZfFjn86pXKTb5279bM5NiFDv
uf1eMzwNwAmld4khgu0r8jFIIeZPmy+1mjOn+Tt9Z/jlFPeJ/xb7tzZ8nhoap8b94IMCfxVJ9Z8a
dIz1dT0P+PNRFu1ugIZ8GY2euakf0RpNDSyt0aa5MKg0ze7zXrIntB2z896T3o2fp+f+/H7Vef54
Tch0pFecmrhAs06xPGeUqJzJT+FNLl/NtZ4JdllifVs5NVlNEi444NjrxyoFCO++jdT9C4Sl7KGg
nqgYSJbNDOoFXKcWbu4D1l8eXUI1d1ajZfm57a5u6kCX4MMAoE3Qj2+FoUdPxOIBMDB9wPAROkyB
NJxuPC3bxQZUxP5VStBU+jM7mSHnSbyE63CFeAzNYp8vAIBEsxeepOktHvBV5SWfgywc/oUUwKUd
T/fXEhYb+BYx6ReeHSn3SK6kUKGgTdw3T128pGairqS30BEWCIDBXQYqFAGThJPVdtO5huAc8M8s
Fmiq4P3MUw0fNM6p1fp2W12S70EGUp8BNJHF2POZMDDLWn8jv8Cs5eZ9M5YVovrRDpr2UTpfA9EP
qYcx+3yy2VJ1to0RHYFH5kbZJGEesuEIYvRTYKXqJzzBez/P1uihwR9wkdjmsTeRMYFZKLIEmnhv
3LFq0BnG/I6lU11kOypq9TgrukQvZs1FjIzoKb+y2w7qcfH70qlnLsSkRyG8tfdRScqtf2SUA3oX
lmq3/tWOsCI79AEGJnWr7T6BK1+Uu2Wju12XYCC3x6xmLPfP0V5Q07R8eMfndGwziRmAyctV9Q2m
pwXF8jJP5BBWPe2V5g3MEaPmhWOkI4FsYOp1JSDXbT7XHal82+rLwqnfLAkqXeowVY8OhB7YwqHC
N0SVSF0HUBagCX/F4AnJ4pHQCISGK6RWHLImmZiVOGpexkfC0MK7dWiYmRG4vbpgrwKoAtamAOMi
e3Od88nIaeuj/LXgMgpwD+ffh6gj649eY9iRVvMyHDqShjYRYsxbREsHB6IBKWP/bv8Sz4yykyWh
uIqR40pk9BNLpNZsuF8Uvv7G+uOUBXY6TJp2smNCYuuR+/ZlVaHJ4leIfHLDDO6Hi/6ngUrIxwDn
4WQiniDaU7DYf+yvDnEY/qIaQdfxNghvvwFORYOIJ/8z5knvvyYWsz33Ts/clTG2oqu3vuT/ocic
dWTFhXaUAXgg4soDOqgbNqCs7n9IQUc7a+Y+ye56hi4IDecZCSMFj1UGk+vu4dbOTT5oNUnd97EF
iugcxc6ujybjDCe+RqOzJw3/ULoTURsb2f6m6K2m8oW+QlU1Mpr+3mUDt0H8G9K26CuyEMRCVxEz
Zss5KtZZY6i+53Vhve3Ke1Cy4KBkCeKRIXTBvZZzHnx1+a01PVYObU0vd/4iCWYq9Ua/nU+67Hfz
2ur+IkrnBSSuxhXmQGy5xVrVa1uLZJPA6/tKtLp40I0NjIxq1VbL6ceugSB6TaUja6QjNEtDlZuV
3lGcYr+evS9ptwUNUEZFIU+vMRSxsHrr4scCoI6w7pZKXT2UMUg7cYF4LGF0sxRgjLKbWtQp8hMD
pgRncRCnavBiIlk3PWGSpi+z7RurhtPmh184Kw0Ymudl91tvuq9tknVVcpz5lnr44e4WRckbcJ61
7qkdWlUjRXfJjhOIJmqaluXZf2oXzK/5VomDJQ5U398XChMtsQtynpqUACRmkO/Oq15lKiGFdiH3
bZbhC20yaB4EnBjSJC/9DL8W0RBnmhcZildfqobo+lPBR5kPLxYA7bLbMy+hIGFJk6XGt8BQf3MC
aT2pxgG1Vv91yZOOVCRDVR/IGU/jPaeck1feEv/HuvUQH/yQZmO3hXSvGdCrJIN21+QBCQO/fhJ5
otfHYlQIrkTynAnPz4hbzJCSrCvqKxjBeErFBkCGf06TRf9WcTQOo0fILXZ3UMRQsC0grYmf7xCI
NuW8ovzrH3tQwY7g8jCb1d2k5rv42qkEHPAWuqa9lavxH2RaWKQw2nfyfBQrdFBpKUsH2Aw+yOkD
6OFBzUpZVmsKk65ktjtmGD09mUnB+y1mDUtUAx6Q5+Jg8WHArjhWLZfsBEHM0IX7xYV0z/6GIwYA
hoK3Yf8yjiWKyThVrJL6KbfBZ5dpk4s6nD0XnLJ8lgNpWrspjCnY4cNYr9OMovGeiNNEw88dkzZh
4SpVb8GU8gGe63dXQtoIskeSUoFyjaGXaZhEf7fwetNNGer9AMOWfe5UUWiaOh0ecfCPtZImnfmQ
/4/m0UPydwCVCZHSCfOrVo4lkPrZeUYwOHT86tiItqaPfhHO6x21l55Yd+bITZSuQY7bWbTUqoiA
uB1QeRL4IN7ba1EHswk/dDsvsL7NUNU51MqYCrL27ATd6Q9wnmT8M7F0asFfsiuu4njiYDNlTqXJ
zB+yUXoi2GHviRfeUjl4jk+7JicbAM19wO4Yjp6Fu9Uk1YfH3OiQXg4igriuyh7henkALaPdDXxq
M5hLavXs8DZgShjdqEhcz9OJHfVqe33hvNGQbeL3CZWyANd10mmJT6M5S3qSig5xatzjfDfx9qys
anKUWsqfGKHSTd50Yk7MxQeqjZoqin0E23efeZqHskqklad0b2xqPcqJAyRMEJpWjS6eZhxL66Ol
teg5AmsBz9CaCs06lhOj1Tab/OEuWB7oMQ7hnuhk4aIBkVurUNEPvf0CNPnumHqiG3SPdnOSDuvB
lqmKOebVsjSGW3TDtnjVJ3eif5gUzLeQsTzAukZvEqsMfeBamRsSQXKG4OI2E5xTyOghdZ6AN4MO
6Upktb/fZ6oRfzFN3Wpd7VMBUsHnK6N9hSwyPWk8KVirhW5VkwqvxJ3HkkytYiLLtsONRyl1ZX6w
ER33cJw98Dr1g20R2xsewpPEIEYXGLxj0Sm9DSYweHRnCvhfGmJ4aT93palH1vEnwopOrcqd+AX5
9546T4E8XwQSptFBEV+QCczbd98HZCrZZKsiJHkX6zc8TEsS8Ngs+S5y8hgpzuJ7tJ/ZtdY/q1Q7
CHrw4iSzRrWUyIl6XNdm/GYeC6rKWQVOfkEutuPULezNbbswyAMJ+nwZy164LBzGYJJGzel4eg+g
DASQ41CGwQQ594v5xlWszLjaaJcc9PBOoOxeSUAhvHj/nBCTt/ii4hcCcW2FeUVIoDeZ16a5KvKN
TsD/pmQ4lRIl7n+21l65mfBrbw79kodq60ZAZBPhP6ntRJgCY3HxMPCaiiNeGuynnTTHOOj8CSse
ItdHW+a/wpldknuPAsa8H0PFibdWUxR1lzVW//t/o/Hw/7UZhr0nkRVghv2t1/lRIBBZsgaXJ98X
T0GH54xunXocqUv1M1mXJ6IPLi9LYCMUGUDoBkOdbaC9ZyRl00LUQy1g7sDVPnyaf09vBR7o9Zbb
sSfapmtwW0ZcBKtPR2ksYRDUPFSZfla1b/p0uU9K/XWfgYYPD1woMFCdUBqM3MYCiu9QuA3zk2Av
RezbfDSLkwe+BxyeC7AmbL6yEkKOn13xKYwjttTVD1dsnjO0R5nyF3M4x3Fnl0VaS+18ib7dPP8X
Qrbs9Fr3574T6POSqNKwpP+KubJ7Nj1C6r5BskbF6o71kLhHE4cNDzyApv4ATJnlpPlhCdngUKRx
C1GmIlDYlPMxirEIZV4sAur6OpQikfxZOeBAHfIAGvXcJ9h9GqLYrUsaUu+SdxttMyF+AF7XY5Wa
HXaGPZGf9SCBt5+c7mZ18+L7B1WAjrFMQ+BEtjJa/9PgmilLW7KRcP8S3ugHsLzDgGGiK4r9vdcB
/cLIu8GBtfu2GeYj6l6aOoj9Uax1NO4lccKN1lYFWzTIiHTemzl9fU6otSdpaY0Wp1+s/np6KIA+
ptR4J5r38SyCOR3EkczX/ebN0U1Ojh7ZUU1tYQ3BsdQRPldtrdihbGgcOARjiQUgih+tZsf8QYEU
i1Eht/yqTH31skh0t0T6CpH9mZqfouaQwBj2u3LKiG/tEDUWTjFAue5oYoYoVM7MjNnPafntV+cn
UXpXVmU6ZnFtCv3S7Tf4wOTo1IOM8f/Dy/kGxhUJjoj56GsEAo3NfrS0Ohq0c+Two5h3OFZ7Xecy
Pp9KER6x/FqqBGkrPe4wfBURZWmJTHEVTGWDvLmYmKTh8Js+72aQHZ0CaE5OlxAMZ1o+oeRaZRqH
U/hdS1ggi8mLGphHKRfnjiNHGekimZDZDVcM2Z8OD1K7ls26gfcMqxxV8mGlXtChDlvEtoGTZZXO
4flKRWzkXwsqCDZji1eV/v8dRCB2sElH5Fg34tsTiPrbiBLwbbebc8PVqM1ENQ2DlD0lfKauINz1
HeQsvqf2S9/jUuZfmM9LyyOusmZdHsDx7P7kfVoBUz3vpzOp9ppHWqa7boNK2qLJcIxw8h/omjh7
lDlFs8FW91f2jpC2KWcnfevPUsgJ88x86bbqWlOpXxBk98wZXcEqf9n4iJFV8JQwoWtTYhyHj1S4
Pga/jeWZw0rrEmKtDa9q7CLOh49y+c+CQFf6MaX0sFW5FBtZzpTcS621F+mLAXVg3n4+Q7c1/5RC
fUc+EhDXaoto6S1sTqKU3tJzemw7127iKXRQ5B9aehj6yWBTihx8YniJPY1mikef1ZKNY9gDaCwN
H+zhWk6GFt9zoNvqwIoLKJAX6SFf7x7wStP8aGlQSXnw1SYlysObNnanfvgVjKPS206EWCFe7ZFt
QwN8hHUv0tKUvyMqCzKAximaFA8RKyAM49kmQr6mhpG4W4zLDA2HYCjiMiqPqzn64bqSa9AQJyQJ
OW9FPekXVTGqREqmz/9coijE+bpTpfd8iRPX2FjSU6xU/9loS3Nqh5Hck1nlrTBYXOMt+vYtevL2
AzHBDuxwDvvoGCOvVR1CscojNmoicz1Kqkg16hxAi2CwcRZ+HRBEGICdHWj08WfVvHOCwVkOXbJb
+RHLuFjxxz/aJFyDuwGObWSGSa9EzvV8e/SE4d1iSgWIVkw81piAc/BWK4xB1oxOnaFCh91O01Ut
a4ZCt08kojaAWMHw3BMOFncUHwuDc00t2/bCWcscyygB1JHdUzMxNbQEntcvWU1UPox2SW/6/YD8
5qjwWR3nY1k536ZmSXKc8zpt2K5VgH4wvIvtXRfeqHmdwUEDLQOvyIpduYf9M1Girh2fTNhxroXT
yal7WWP2sd8aHpztG6DcVa+Q6IN0UAE38OvGDHDNBVaB8AMj4xxfDCwehyJ02X5H1xUGODMs1FkC
TJU4AxAhlGi1HmsQA1D8JKCxJ/YLGC9+tmomsDR/TSe3yy17AXQSW4jX5QLccUNFCgVFsSNvc5cW
tVwJ7ne63Q+f8e3nTPQqQ8S106/3d4STuJiPW3q5vboEd3s8CPLvIcCvO1wHol2jk0lNHY4KbamP
Cc/JX5ptXEWBA8LgKvbn2tmNgMfhldf7MP/ONMdOYKJTMJi9S6X0ZJN2ThHyl8pHrPNFetJI1Mr4
+F1GaQ2dmNG7bJz1G0Il0+bcqY7DT4I5/RM4etr71BYZnxG50RbiW8+ht+y+WGXNRi00U6qRJFpg
lWkY9I7oGpH7aLsk7wGOWUy7F7HhpQhPxXDmwTGssFWIPg8N+IB/QSkkA+28aIMHT8ifys59tfC3
XpM2i/YNlsdJEI8CxY/CkiLBGjPSP+swtNhhSCwCpVExjM4IwXrIDsAKEcUXdqqiI/PQDquVXhPZ
V5mSgMLYIwZ/nJz+54h+v5PgMVAg6TyfFgisbj8QSdk2KYJ7ukeOuCyxfYNCviMq/lSStrXudi9J
jyDsZEShxP/iT027fOrrWNssDksugLAYotS0pZJGDkAUyfZ2Q8kTh+4zRRcdtKaHi/KVn0vOmtpm
5eHWQbAfFj6YBDwOkwY3TUMyBZ/rE4+yb2tmvrDG8sSO6+JJ5fQGCBRE9CfbNAvEFPGsldN+gr+A
fRKE2jXtSmI/4lt+oz+aY3V1hXUs3lyFk5hegyEnQznCftKvL6KnDodiz1NgxTENtQvVVFtjgOh6
OuI95bq+XAInmjHO/dx1oW7z5lgfmeM+eC7tEXY2S/vqPj5mbW3tqpkTvXQGe6pO/8Zy9KhDYP1h
UV1F8b/qznwW8nI6qsZmNLfbovV22aRXPfcDfe9m8cGSZyQI9UsnhXzins0/mX3f2AzpyBq2p75G
SoBY0FVic2DF7hZF8HOcvbDwzax7vnam2aIl9aJnUhwGyO4cEna6FaJV/QkGxD4jLNabL4hb40cr
To/xBDVI2ndLmjoYpkJEdAXwv6J/6UUqI56qnJPvEmPuJQoqoiib5tITEURaPeM8U+RAhpUKaeYy
xrXeMGQ6QaPb8G055TKT1mquL7aAZG5lHh7Cwt2IsFcKZg7/h0DvpzRCCoyCKxKqXlNQxEWCOAZ/
qTBPNPMz3RZe/EHc5HnHMKGrBJer3cYjIPU420+rcEd0gh4apQuM8yimWFCWpJkUgYoM4yisWxmq
nlgnzfgwqxMVXnGTixJLBz4Y7AIDALodbmZ80n7MyrnHIipQUbQ1ASZVrmZfkMn+yHgfy1NNWIH8
1Dpydwgo9NYGsMn+qr+mxES61wlZB1C7BVRETlaBEzEbm/fhVppCjvpDyzmfu019k0ouSC3S5hgW
VPgroPUH6oJljYuSuqJz5mhCTwPYTv+kRHWQsvL1nZVXvBD5EJ93fi2Og1v+jIsFDa7AIjXDThVA
PX9ULt2MpN0CJbJXkzaAhGbIsuOUYdwgaBr31WHNrhDbXPiFC83qC5ne7+yNd1iRz/P2UCgc5u14
BZXqWXc6Et55LSGm+De/yArdTvveKYTaUaysj6ASROAt+Htgh6oIzpkhh9f4+20yMvF+WSzNIVGW
gKCUpt8cu7VzSiktW+5Ndqoy/sRxKKsWKrsi2xZueVgrnqtLjvw9iXMCZTklb2ovHonzNBZhQIey
t5Q6pMTCYYYMwmAdkDBKGS+9SOxW1K0UOIjmObJEQpm8kne+Ve5Pa7qYiIU1VYfaJCuusmIsArsw
trQyQ+yii0CVqcZMCS5+vquLqb8FsNB18nTCpcZkeAzbC0fiXCuGO2LSTEpW95SNAtGmKSukGkGM
jPT2MZ1S+OTzzxZNSn9K54lGskuHCqylssNhbW5BaHyhGK58ce7ecLQioqiasV4dFKjRVDk0fknD
FgFgnTpVVsaL6c0403Nz595QtXhsujfeN2I3Trsj+c8V2kNwakSUZrYG/Cgm8ZpltCqtA3og96Wr
RoX5IAbBNV899KS9BhPp8pV6CoIHh/UYCDQG1QnO/qd5iA5vrnP0Nt+psBhJzr12fAFpuBQJZ7LY
yAwNiGGuUq8bNvPyvByuTN7pjN3iN7Rgy5IqyzSkFTulWjOEc0rdYCJ6QxBuKotPb3jcze+gtcyZ
TipzMCaJbphIQmRq/e8HvANCX52x6MasC9vBMo+BHiHJYzzPhUwH7S1ifRJj0NeNz3AXj/sK2FaQ
Sd8MCloyH+R3EOlW1DdbjujTvzC6j+AEk7moK2abmcsvfUy9H1q2tFUB7tAMQtd+2SZfhzUvyUBj
zi90f3iDvlDOYoQ4OBbpgi5kmuydo5OhXpNPD8pluYAYi0jm31CPaCQEUpiO0FkDhJ1tqc9/o9uy
RlJXsqZMaILElB+7OnsRhfhFwEnw+eOuEX+79TOSBwHLzCs+5TilHAKXJ0UTmX19i8PqcBo4BWsI
oXxChWJiVQDZez79fj8QNeHch+v2xduaR5mH59vOjSJhjGnNTZ0rnK6pUi7biim9GBSxb26YNhZ7
GHsC2eixmCUWj+blPfCdpJ4w54bm4ox3JQS08SEhQJ20WvZAcFrhvw36tdPw298luU3HrtpNPGsq
aoXmogqzxTEM+Pr+h1gqsyN7uSW0cxM0AfGMbcUwl+jW4W15jq/QQMSIFIZf94QFGFqvWI6EtU1m
08waIVhfs/+Npmf146GbJLCLim9whuXXRBC0Ea2CV/BVoJ6LoxqKw7WuEEdatsA6MPldXFa0mwZ9
eFjO1TFI1v+auqFLX8C9r4PEdE1YJyXWC9gw93N2nCrSAihyR5edxT/zMj9hNtZwNb/LKTvL/nOV
+o09D8lLPzlQzHQq9MT/8MVFjOrpkEqPXBtK9Uijmj1FFGZj7mOVl5eSNM6XcwzInCCrHyYKIIMl
qJYQYLO+7aPSobN7B1Sl/ibdVBZxnEaL3W1zm1X++yxxItoTPWzO+GuQkSypXhArklf3k7I+ogYy
+qc2ZQRRxHQLqf39je/ljEBAALts6TJzltq5kOD9/ECyAaUZX5/LgKY6T5YWaRRhItB0R+YNYg3s
BFxeM4754J4/peRash23KtwC4Zw7H8B3S3z8OudLo/JO4CZfTD18/nZZR1s8Hba5p4HSn36KrZwo
MHeSC9nntZgo8mec0+tiDTxmaekNV4qNfHW3BOfXERcp7RtmXJlJCilxkCbyOZj8qGk88Tk4MhOU
ogsWmz/xhVxUUdTIcXMKDhMf4UOOnW8O/g0s6WPbzU7YaetDZ8971uK/axK7gRxe5FTsfb+6kpCB
7zeaCM5vDjmPiM8LmYG7Yxj2VC8o9MfCKkPuEB8Dzv1+ojOlc15ReBGnM5VrSU23tRetE+GZp5w+
dLgVqif6ddShogcLyFvRF6UqKOhLkhcXpOCLX/5G0t3vkdWxB+2nB08Nq23+RBTqYDqcWqZYVPUX
B1lcVcWHmTNfHz8GsKoAJlRBhomnuM8I8IGudZv9zcsF9C35Xs5VY2e8UPwv4lW7P9T6Bx52N5Bn
auTEuljGBr8FG1VTG5qE3Yg4AOxiUXV4/FwMA1FOHNRcRd90bMOBFE48hl0KayHff5d6tRWM3ypJ
yZX5TZqwmXokD6X+ORzaNVS1MejooZmxPtQe0wyqmSery0TPSv/xE7hLMSgkPrrg7rxOf/rH3iZE
mr7lILDZzpi6JOewntuHyh2WmCmBk3ora0ESEY5ollpu89CXGZCY3Y/0l88vW82UEqPYuixmwrO7
/ewaNQJfg1C384TA91MCniJWKE6ooYLaf5p91WK0B+m3vKVfU6yg+BmmXjcf2lpt5KdTHBkgUxRR
IhvkX2WRvKnI+LDKxxhsHkxXkVmj3Cb9EyaDCAuPu+ERM96rCgpggv8rJ9qbkCDYY5Cy10jE3cNt
1isXiCX7nO1yvU4WT8OMfg5vR4PriKQ90aCwfSGzdHVeyKp1FF/JC7Rjevmtox6/YfCO/XjFeRwt
qF2fqp1AwWdGCMmkJjxXXWDRPkJBuQ0h+p9ky1PTcDH5bU5DoLINH2f2B3NrzovpgqYEFjG/yTqK
+OOX6OeZAGWWEMnbqwJuijqVVA5loPODiUssSg8VOoNjgkKqmE0+einC927qOMNzLHHoyYxq3Iw6
kTBkmd8ZOZqKUfE2dX3xSC0dgO3r9MjaSBPoX8LbOvqVb+FyDliJ6BLVWys9l0a92tS9p2De32kx
vZaxCli8A4DWRzcZ+KEZ50QWEBT7lfFrLwK+U+63KsLoIxDW5evoubUhSURjex3G2hLAPmD7XDac
y/ctvC+WIIN34zyLNfxcjt95GbtDVXxAVopVztqqyrUU7G0ZR6fOASKoN0LIT5PmcEqIjgWW+WmI
p1c6XHiCWNzw6JWtHxSdVmprmAMtsMFLD3HGH1RQZny34cvsCKoQ7/KQbwcgmRPpieXcjUARUlH3
036zipr6TEQy1ZI7EmNRgHLvPJLMW0S2GB53VwHw2lnyVIP2feXY3y2wt6ZLSbK3kQ2PhtuoYN3T
Z8kBWwjZTNdHzcLiowPp9c4WpPil2exiJhTwWrXmVCUuRrXqTkDlfZ/bOdVG7p+JOz74jFrGdH/u
c3Ci44DIsIS58N/vxngdP98dIwWgdiodhqv9+kzOHFtRKJrdECCcC4w9daakAg3dWNGNUh1b9NyB
vag38Vf6OULTy3yI6zRLWhiWR7RLqOpMwzOMv5lDwgGAv7eNjQxifKZWtsR9aumr11OcHIfsGuC1
/EPI5ddhmKdbQXbvAxPZvZGPUbAG5Jy8hBgbbZ0+eoBa6Vh0ZeUsFj5pbB9Eku2aWZYwoXRyCU8K
+onDvPFHyQXwcBxfGN8L0lMuj3OLLMb8jSOCSBNzvUqer8AZ7EzV0tNDKynPDfN+DN6eWi/U+YfQ
iAJgNpx3WnUWwoyHvxaU+qTrFd8vDbZCy7dz5RxrgYGjJYmplSRCq7131i/JZiC/8eh7/ZcHI7jo
W1rQxqcmerqe6Eihw9vkC+6TmG2fq/PC/yet4YMaGB6+owXvKB0bFrDc9HkU+8jwZ4ys2PTIfdES
ug9ozq1jVWu4i3afoX2pd8kbCUhFV1YU4QFpaatfLMvbFLCZQTQU++dYxw+483DpKS/LKA6rKWl6
j/nK0Im6+QZ+nY0cmo9qd1TjYSekOBRuA5WXXU6iC2fcfRD5f8veJclgms6upFI4PDHu8EjCq4O4
VqgF5I2DlU/2XpWhq8Ib5dkDSG1+gYZI2z/aSH+buabj+9ACt4Bg1pa7YAgDfFWkS3nMwBgXpfkG
xoUd8KbW5ja+1kXtOeJ+OytMJZ+SgCBBilWOwNC2mwqkyIvwx2gdzkmHLTvUpS4kwE/xk3QGOK8x
QMGxT/T1FWn4SyBFCyH6/CrIv5+9TqwS7w1g0gdIKkxoX6V24MpXbisL6nfkSTmJuflRljawxR6D
MIJUQxcEIFKee8D2l8Z6t7uFNk+a7OQYQd1Ts2oWq4B4er4YVC6qWyb7rZKixepbcCqChytsF5Zw
mq2kZh+7XsdGcIJU6GswBCZbF/pfKjBev4tFc9ykWGmHlxrAjP4FuqHDnHKsDS0YgCthZSrzUeLA
Av8crCf3KesBJMDZ0/T7ulSlnny3y5XwYUFZ1kzEJKlJBWGGDR4Ot5jnjo3ODzC9M3NnKz+YGVG1
g7wnxXJ4TVpdPfau/B7+RVyIEJCH2lqwKVALiGbAKG42y2+RPyYVU50I+D/M+t2eVFOkY0kp9vFw
0uNbjFlZrXedkIktFQeEXIm+ZqfGR9dYoduIS1XiV4SI/FU/qnPfw43V8zjKeY4kEMZMCRss+viD
r5sQOBjWMNASdwdfz0rBxJsIXVLeTtLDUG5KtVZyczE5iFEFV0fCZocKithVDPJqGXyRJehczHh3
bzcAN9I1mQZakhNov6e6o2AtSqxLn7KuRuL3XLbqmqqWZyZDVle8lliE+wwAsSxGQWzm/fFTZGDS
RmqhJ8hokdxG2UjPxost92IwcfIkO5sMj8hKTZnnvHTHY6EXGxalc+CsyqiIgFd0GF+IdXRiwkZB
5UVGwItw6I4AlSr6M91/xSiac9GihruI7kDsdk1eFBJirZFfujzqIxg7bTOLaDGDpzehnOsQe/oH
wOKZybnRv0el3MbHiTVQgO3K40dwStgxXX2QcBBPjKiXj0D3Ndz1gid65yQ+PdAgjjcQTExSMr/G
ZI73po7GEcXymqIDHGcvIRZa+h7UWzueAQU9V7MWAWFExpXnBex3bIVgKaGDsk7ekdxLlt6AoTlK
umczoKLJDynn1Bg5B0a1ajWkV4QVGgmCZ2wXSIzOv+bL0oDXo1HCT2vK5gyewXkiB3r2gmfDLQtA
vP57fM5RmNyZBuKQZSI61rgT5vwAw9f3PSZ2tyzAfJ3N2YAPRJwpsEaVeg+67IYF9uPPi170p4+2
4uy/jZy4zJB1PueqwWs98hDWfAQ4yvlZ093TwxbVsQIasmTZvHuJrRzXtQBk3FTYIXOtAAQJj5KC
RnBjbAtwY9LSaZTDE7zALuUgMzy8x32tzfwVwLMohADYKStgex1Uk0Djigl6wAPURRp3KvAIjqvn
ZPX2i6m/lJZNIp2N6fpy2+fYs/CWGz5+pqKrO8EI+o1gYUgsIC9LN1w6TCADxZ+ZjyJoujxyPCSw
nBWB7r3j5RKgOOQGeM0byp54un4BULts8mG6NVvHrn8aS4KIf29oqjHNgIiTkTGYP28xcx5XQIsJ
BHEH+dklJdHqPJ2Rq/ZcGtWH4VK/nWRySkDs7zOMMHaF/X+5y+9MeZwGHCja5vjKuEgommCLoyJ3
sSN62eY+VklJK+eThYaY2eZhKhMpZAZdfb5vCMNyv3NJv5OITbFsM1eZbDqvHz9qUHXvh286SrL9
PXNyW7sH2I2jbfRPFauYmnyfxmO+sWAQYcy0OzZhno6r7spJNgZjwLCL05qOaBoGxhm3Lfn7iILu
yvqDZDrs4ZcQaxHlFDp7Dg6cLP3jafvXvrHmJ+RJsZM5ML7d4VMnSwVPDmYLl62AXBz6n7qQESnN
dqGWCOlG4JiZYN/qY+WG7ffPPl/r4WoFP9DUg5VB5I+h67MXz7fJIBFWxESNHJMrI3jnC89mXPKQ
zyx8XncYdxZel2RBBx7CJ3NYBd7emSbb79ieb/kEuuzVxpZQwu8rm0Ioi1oSbzX47ONKD11Naok1
9gm4pG3RsajOzmtuWlQ505Ql2x2krjqWo+usx6SqTh2yzIL+pl//Fv/J9/CnikLR4NtUlkwi0nNl
PW9szinZYWwWck1fgVYwOzNFHioo27BQh/G6QeyqK4lnPaceqchz5UYv+zUuLo4EcTCYsqoY76QE
EX8/Ise9Be+oKXFdz/Vom/q9fC7zgrSg8s5/m2L1CXo7NCAOdi9AamxGq+ePrarSNC+1wf+diw2v
Md/knGPFY40/g0h1b+aikz+ZOhXHlwNqe7S/AZUktu/HRD2EpumGXVmRLQuxt8cEoDVhOGsVj0K/
ku90CMWPZk4RMZQe3ToaejidJgUma66+tL24RHTaNafz0xMwCqF3zvfPqLccTTBgqbSyD6xD+SD6
xoP0VW/mEGVFAloYMlcA6cEDaWy7Fy395V+8Xz594mvAPZzi7wmlSiDI/sgXA8srJrheJ78+CHo5
/oXkIx79B3Nu6VmBKahpAu0NI50dk3E0dij3JAntSDwzvlwKoKEM1nY6IP2p7jqaNYF4aHDjNyt2
ASr/apar50INdo6MjOzpG8bE0Zkr0QXauAMe3GmqQPDcpWDM6pz9rEup4MbBO6l4KJ0MVAGWgcsM
asiM9Ngba2eOlFKbX/D9uaoywhoyBZfo/W8UWjlUgDN7dpp87gVFLiTtXF91j0a3DdVuY3jQjb8h
rGpvpTqd0yA1sXkgWiKFEq3tWrx79I+MwdxiX2ulfNGJ4bmoh07N7e79M+1D/OMsUCEn+DDYz8JV
eMXi5VLulfkgZuTUnYyyqvDjOfksCey2gn3wWn4iOe3vBl3vrbuZhdxzwY335xnotm+w3zNbTFey
1VU3uRN0lpmNi4XTJCMYYOo0JXGOMYfGXohlcKn9s4tWuYFFphr3cvGuFxEXdQlNh86wdqEHcAMQ
TMctGzMrmBhkIBQ8WDJoyD45kwvEUxoqYooLQgM6oYVHisHer8b1paocfl59j504v7dOV0YY7gw3
CqCh+2zabi6hLe8gZiKFAY3zVx/m5IUAMSjLiZVDklJiss8sIyXsB34cXg/+DXsx+aKPGWJnQaHp
NYldyxgFDJgUR6iqKs5ihmB60/4Y9T6tlcjzaCJ021BFqKNG5uT20LLoo4Kgz2m5omA1SXhYYBAz
OiKsiRD86kLkuf9HP0ypds2NZ4n5k3KJCzNWorI//I+cB/EfobPeV4sdtzP8XDxTCArRpvYtINyc
mfQS9d+Hx7dlkUQHtT/hExZOpiwaSh2j5K+fm02nvky6f1sleiQJZDvq1PE72Dv8wFguAoJcCjPM
z4TFF2n7FADsRvlw9bpPliHc6aFU7wMvsr2octgSMZQDHneeChya7jhxoh7AFXwmvE+BrYPptYEA
TNsVwHKGap+7kB8tnpHjNmCgRLmAGsyscHszOKEnoeo0es18ZSdCIhElHPpKDWDgSkUyNBu/xWVF
9WbEoYZ0pA913OyiaXC0zHfFs3A2zrDy1PV0gRtRXFa7D/PqHWXi4hVNeGHoJ5FhgFmElOtec2VQ
rLmxcn6c+TLxLLfa5+dkLE35PFGx52EHRA5LUkQUKGgwwHCX47mvedhzX3lbZYi+9xsU2nIykp2V
0BHKMiVriqKeiVnhD9LxBbNjRsqopHRw0ajGGfg8AT5BioPejHjXAFvqhEUg+tTLUyuHGbfRf9hd
719Kst18Rsxss8Cwzj+H/byqcIcgTFDVuKQ2B74t+XJd/PwcAXX/TJXAClUFCo9n7p+o67ONXHPB
/kihTquseQhfe9IP7T3Oq8c7yn2a4YFy+dtFma0vL/Vaz8aFbYOsi4WZK0B2w+w0Udtb+J6lv1+O
5PYpr/h5IoW7cuD4mboONRHtrdsLzXa2g1DGQnZS957WZ30H/kJBm7BS42rK/wnxNoSkWCONZ2ru
qF3oUkbxgBnYbluY+VBhLX+/hqzZo17ktNmuQyzFkFQG3cDTI2VQxL7RkxroAolsFHm+xoDGnx+I
5tYEdJy90/M+3GnBNr0mtzFROzBKjhyEy1GtW5zsjNwFALjjnhZ85KrnXEcKtY8cpcRi6RpvOkSe
WNY6nem+Bl/ysSgsVAHAGXE6+m1w2wp31iJW5c/tIkXhSrwJOZiU2J99KvVV+ITEiKlkKMlH19dF
xHKEIGWB0rBlVel+oRRJxn8wbqLA55UFieXFPQGh9o/S5gP8zAkrGki7EiTExjvcCZPDWSccfw3h
rmPdVyLXNswa71UwiM4HiS/ttBjgT6PNwGOGmFJ7SISJFtc5utIlIGZk/rWERvaD0KCa4nN5m/qw
WueC0GI2wBi2YJaY5/6/zNecL2j+rfiHeC75eZ2XUTub0I+txzINN2hB7/3S69Z7LHQrOXoClQGH
+L0MxSzNIGQ8jlpeKJUvECSu4UhqkoKVgodnSpDGovKDafwwJOLXkFrihae/AVYVmvuj/G/VsW0V
ytAJSiuoBtk+CkPapQFdCW5ZJkbtBFNbvH7l2qUW5yLEmri4T1OLYevuZXtR0SPJUSLPX3UAMyvF
7078AxC5BLgtU6P78UQpDlK8zK5FiBUtMCPEurVyjZd5lienjdZ9K1IyJxDxDHOvMzk2XhIDO56N
2LWtjeONFD9k2K4vByce/f12BkrJALQVa+tHGr05wFa99imdXKDYVUtUb995zgglVt+KrWYDEjKi
GdTlb+pjV24vRyxqHCXIJodd0tEBrVV36HtVdcpn/PVSAKdURUz/X5hONxaeBqwOCX07PhOvCLge
BdiQrF1DalyuCjMnVWk38RiWSzZJVONTztxgeLiX2ynF2S+V2Zb6PeXlVhsG9lmU/Bcn1kczLpJ6
HCfuvn/T82UETMrBtcSsGzJeHFCcDTCoSQgJ4wmcjD/B+YbyjzshDKp9RU5t8jvYFuSxgzscGo0E
JfBMJurb4X2wvSfNUyjP1+P8zVCZhDjYvcB9JZuyJeSO7NWeTMB451+zPRs8ie2F2OjWo78wyYyn
TmQZjx9soYCETjzAep7Vj3Jd9CvbGhrlJQ5XiEsm01Q+tCJ/Ye4GmuwmeuE0SOV4YwHsrm1AKjmq
7SpgDclKatEt7jZsO/wAx23GIj/KvYu9JMIV8NNqo1YznOefHHInCsFzS4Jfhql8iHgJArOaFYRd
MAHbxjd9Y6eEAwsWcAg6jbkQssG9UDEpHQ927sjwJhpmaxW5mV/EWW3T1mbDXumeQjnvljMNhGf7
145E3f9+NCyMQBqWnUwoiRzwmBGHrqwr9I9G3NKngBVCSEj28PTplArpBWQOmYrn+yhFs8/LV0eQ
YAm62Jdtqw2YSu3fai499tI98mQcIhY8MFBMYzyfxHXfUNjfnV9W+8e+ptMHy5gWAPrpRUmfK8CM
8GMgxDJISoNFL1pBaoGBoYT9SC79n7BrhAfx26haahycjTsyhREw86wTt4tWTCy/lgeDO3X+23s0
J1BXgT0AzDexu8+mb2rp9yHr6GOmuvyHEQrkktuF6+iXmwRrD7lEOjIQruEkTbzAWui4Hwv/CG2q
cM3dBdjVTiDWLWUV+Hk/qXN3TZevTK4LVnWd4IgRXaeNpmd7GHVZgI1EgqgDGUAc/NzTvT0Vtmrx
KksIHWUpZPa4SM6IGg+VedLtazNpkCGFpHCiYAEWCAw+mLYyqu0/yaLGi4pT3tuwSaZtDKdBI8vW
9toGLHR6fwwnh8kXZL3kUzuir9w4H5NkjbmFKXhjfKLhOc4FurAOMvIF+aPiRh3jkP4e7qnlUCM4
Q3MCst9CqnLtCP21/h8LV3IvO9/G+t6Y7pzlTgqAVomNcV4F19/eVlg82+9gx62P1GAjjvcdng1f
XdXYxG9qXt7b7BpUa0GALsENJ5PUE/cdXB33JcAia8u6j1z9tFAvXx7SNplEhZl+2oXshObn5zn+
ovIydmLunuZFVF5yw/jfPS0ogDDj+Deb2+eRQy/fR4HzjyQBhKcKwy+H6lICAWrPmR7ps0kATFR8
TKqtTlQHKz9FAd3LUsFrvQklYOMNWsq78A4UFPDuP4GWypEi3goQqV7ATHIhHAERSQR9GapmTZbL
NDIei85a5sfeoSTAkY7RxPsMa1JkOaurhLbs5u+pl2TGXbHjSzgawzL6y0wHypA11QqlV3XnIeoa
KFbOcV+nX4CXvdTXrAj+cGLpX/YLvkACSZFK3Al17vvNZJCo7Al5FcnSM+8RhqZnpaduMdVzmzwM
x7dXq6mCkYYQqSTRg3jECiuBefUTdbrzUxGsSM1kaKaoTf0roj1aYRB9x2iXIGLHq1CdmdMb4YQu
sa09no+chNmjkNFIR3XvyIpsc1S/d1ouj+Nz84gFr/6F8siRT5rhFNmIYYCHPBzV+l++RqKzMLaT
EiGs62L6N+Ku2fKAXQkjJe6ZRnmMb+7xpveUzlFMYVZGagycmYv6Hayi2DksTwwh5GG/TBlpN7lU
4OClElDrclMzFg9Dv7EFqljbhyANJ7g6sSkqJcNaTtlbZPmvYbUJF8ZpD98c3npHqKN1Ul839XGU
S1zTccBPE+8TMENrHY+JmFr6eNuSdAyXSUazyknXaFnVxCMiWkqU1NjqHvjSHo0+obXSkJJMFkuz
fXLMAbZtEPUJygij6lmcMOtKvA5JUzYwGggv/SEYvK2mnBYaLWL754KVepksbX7LEF1aCsIoG0Qe
YM/mZc+e5KG0JA34yrO9W80SaabcxtJrgknbR/+l3SIGmG4JJP9YUOPYRuED8zzj6WUAeP3sALsN
gWinrkKDU5K13heMG+AgnwI+GXvzW3oxM0qLnD++9z0ehA4aYPbuEFaX7rCyPX02Q3yF974eBvoJ
w5flLxC0rTG5aTopg31rjY5Mw6XoDW2Rg3WxRKt1Y7XdGcCzs/7/zvnGOR8rRVV/GGNKLhdUOi95
jDtTXQQLWu1pv21sNhFTpCFANDI2Jw21qMk7BEak5J+fRigRTcGdWXzsIH2CxhbpGj6yTP1fYcG0
1vzIuxF0h3Hdrc/Pu5OYzG2qslXmy61caTbbv6GNEDoHDPBcO1zq/Zy1Nl9Q0vQ8jLrRnyxqOHHt
jaZyKLzKo8JWRAa8JuScK82Ij1oxaJjm7GSmcUOXLZ8lcXLTgOU1Cd59ArQHtbBTyGiCbcQ5t1Yp
2gGKDJcfaNmqI/hacE9AJRSI0OpM3Oj1TPndzdIIJtZULTKQbhVlfRonW8JA93VgN493swdpWVWb
OIo0VdfCCRiToLFM8V0qwaYqFdsVkKF4MVl5HEogHcf9CbRLeRS0KOpP/rdajeJoftB5alMztQor
pcGqB98YgDsDDqLasnOImfG+rDpKxmsEYJs9gB+EBgS/hflrqwYbnVUn5nPUDY2+hqRGzN5w6zS/
4q7mZ4rk8lYNqgDRNaa0oAeKbTARAlP8PEnTdq9rZaYpEdaGIx3WktfKgD3UQzfsIUQi9a8ir+dZ
N/bP3x53sdDGrla4rmQbjvpqilLHNym/aLHa1+eODC1ukY9ukwLEStFvvOLJ/6ufs55pApn0kSH7
twb9JcnDRV4du+pOfWi0W8/1KORwT/tul27iHzJxHa36pOrb2ZqFV3PxgPZdmFxoUG0rKBO+Rppv
owDzkasp3TBFeibl+cUUJCI4Ie29TlrdBDTN7dSx3XX9QzplWdpXoxjYiEpjaPeYqLBSTUMoTp7Z
CdbOD93MtSbqz0PAmzQUmrWGV3GvXK6cpsoF59PBGuVUn0F3XPvUFHT927WjJ0hIRe8dGWcG0yFn
bLIkQ6JKDqiOE+772k15Bhk+5sYW+nLIMy+SQjZC/8vlxp4+wN3GqtW1oz0nxhzyG/PRGrBBffqc
zXulz6hQ6D39Nlg9iSGH0SA34WUiUutZjlc1Kd4qTKaKIcRVblU1lE1F8x6Ga3/Gb02enlKs3Y91
Dv92BGxbshtCRpICNegzS7/zSC2CMFNNpeu5t5WHlgLtwZDPEwd5xjwuz6wMYnYghDs6QCwXNoCq
DyiG4Q09Ou+hoAuWm9rrBagDP+Nsln3li84wo0KMuJH9u4mftiuG3VmQf3DDksiw/aY0t+XLGib3
6fLFASr/12WAFHIJ7buSajuL0FEztBONp5TeTj/0R20dBpoPcYTnRklDesOd/+gyYvgcFR95Zvk6
AgwgxM3Iw/ubzTwCciKtSAUKZhxCrD8gz+n50meXn/4yJAt/efVNrTEkREMkX4tBLafEWFeUCUj9
xwgx1lYtj/9a3oyyQKJaY2h7t6Vl2sTAvYzWHFL8GwROzpz/HRrn+HFwZvSU10oJibTCp7TMZPk/
2CIbFhiE0m2VnGmERo1zCqAtcLscAD1fJSKyF9GfslqATdCPHY1O2WqNzu8Va71JJokbVqi6XSYu
I05oMgTKHEPgvvqog4Z0509uGr2zxEgo8Pomg2BPi5BM0JaC4IlCVQbTayGxdSAcHsvyUJzuwmWn
YM4K4sQDcW9DAOv54mV1Vk+22eQH3REwgNZrAlN+DMhkG8nBcxfhLMMPWaujXkSE1uFg8mXxnpxU
8gz5BoA2Jr7h02AlwRGvfOvhEhqq5mNjaQSPjPUdSFJF06aZu4QpPXqVtXffD+Gr0ydlnJkmQUAS
Hq4Y4ayczXtxK2LfReId01YyNsUjGuwMvIhrPJKqimP8SULLXYKSpw8QvwNDu2U87W9RHKe6xpwS
Pz81juo6VexGMV6GiF8PbB1LfL5ky9qyavU2o4Sj4O3CZ9fDfWnkkPuouS57Dwhc3FRPL6jOhaNc
ggO6kX9Uad//b8qQHfC5bTayASalpSsnzwkmWPHT0tw4pDnCadI8ls5YpZ9zQhvG5881uctr4TBj
HKA6wnGaohjUBCrpT52//0Xgz7j2BmCfulRyS2/rlABRo5FYuhn8JF0Xlpd9AD5kqvy2oBzV7+dQ
x6f+IRD2d7SWofvwXRDfBbALgfsnBvs5wY4UOGOz/1xIQP3hvlPh2SNuoOuGljTxW0QDCYZt25Pi
MHsBq6OgAXViPHgHqUrxz9WjqfYToHAG/ksqvu52plzeor+kKamjZSKqF2eNi9aLE9aryPqgr12i
s3ilcrim6wVMrY2RRa0kvMbbFtSGGRPovmDjNvmJ0zAPr49NsZl/0BUnaICbDq75mSWbv41Q5XiM
0ESKLVcwNK0dqtMVpxmIT8MDhqf2YLty1k5N0yBTJFsuHjnKkwXEEtsopb9MpTm1efNns03WkaRG
v47rApjPyd0059ygoE0xzTU1w4bbRPeClkZvRJ4XBJU7V67KW8i3Pi30yLpnEujA6FL6o28r50lB
N0tL4kSOxgZeWs6JEQdcqafHEk+rKtQhsTG2KO8ORc2LzApb80IAQ5UVKqMOCmQeSYEA6h0XQMXT
KI9ALGj0FXJD/+uc00ScfR29n3ZUuiBs4KRyyH6ZLLzRFBDRAw1o3DHjBHrTeWu/eGEeadbUOs2k
1UNubfBmjSzOZpZr9rG1WR8EJ1Wdv1MbgqEhgjzgyb2xrjA8uk94+Oi1nycKkKizHx1feUxHji6/
9yrYP1SaGpQhMgvU2Z+Xxj/hgLp1rAfptSMvgEVh3QJkOLPiSSndiTYJ9+47TnKqmaimpgvCaqZR
rgqwAcpYNCnKV41xikhCXEH/tar1K/TakLHhBMEitM5CAH8M99u+hqH1t06kRTOv9OeqJJ6xQakp
IynD8a24/KXAUSWjF5CyG9tGFX+gEqbPHO2ysKD2u7XrBkaqtap/eh4i4+n1zZYPT9ISjlUfExUW
9IyfTHS7Jc50ELbXorx1SEIbN5M9cAGpt3GP64xT87py1YKMoHKSGCsQS7tLSLjgJtUdAZJxeNtI
gSL/1RK3VaZMiYg9NMsl1yeHmgpHsNFmlg2aZVqg017QcSHNK7BGG52QqLZljtmp5wAis+mZRFhD
kX67R8BmgDNVdg+tPVRO1+nSa0KESqZ5MMhp2L0/d70V6HnKLiJRIcuTnb5BrWQFLaecNr65Q5Ul
klFs30UvJ6LgTyvPtC8oKMCWhqQ6/y4sKPJie+zEIG2MqittzrhrfshHTSJ5eb9+Cr/YGzO1nSfn
MosR6lnSD02gE64QViOdme/NoHKawk5gV62qcvfrJfqHMUTmqCVu3Xs7UQ/9UDdo31syfNKpqE+V
dZFHZuBbcvNO/yLI0EXN2+PYlDqpphRubSyYDdUgU4NkQI0Ix/rIoUm7N3BaJm8TSC4ki+qapQkD
ENYqCATqOL3FfLJ4lw3I755NjvAqlmRe0+rnL+ayFSZpU8K4fdj9OTmz4JUMA5q2lOweO2tihiSz
Loby4BttGjJBIar/vSmanbuWP63C9dBmW7IIOSG3nU6emJ2IO7azNbl0fYexcqbQOsIwdB6T9Okm
VK8kTr7Y66PgiH1l3CQ2pURR0qnGDc4JNj+M684OquR5ZutuhQghaai2bRqXTfOwwnXNCA4+rDzA
2UBXniHliqnpijiwqg+KLkAU+45kgBWI47DrkrII57QZwj29fjo6h2Wz3ySK1e35NzJaw6Awmx6K
udLqeLzOc8IOTmXBQddajTL6UkNHIQIE2vWGAHvt0773KBfcRIoincoq3QSVYCJpN8CwkZ+JCtCO
IuDsnUrN9ruev6yYhmbIX3453FQs985BnEdjeA280BeLPW3G8lMDDt6FY/BbROWgDZqzKKh0wny5
RUgHRCpb7DXqcerGZGI2hQQminH1tAkqk2cethuXPtNtPwqFgapo93FSHA/rlD4rBV5GZo8h6cch
ob6VLIS1hQjDRNudbvtKhf7/uFGF3O29TtkQHpEcCRn+eAxrVvkE9uc19T8NGNk8hwvzl4JUM1f6
etef+n00ELBo4eBRsNABtweFlCzUIcZpztvvGMdQNCW9IKPg0IYpoL06Ki5vtBA38GcR8lgvHfq4
HzyJa2lB4ODkzu1ueCMgjx9IVz5SsHL33pMFWXeCvKT5Z8AFwabpg2NbE9+IzKz4Vqlv2XDvoTXE
wSjTW0Efsmcvd1mWIU4m326I6orBsO1v11A65W9kcjtFRNybBx+Nkro+s6DSDaUwnDzsVEpsyolh
rzNVDpE3j44Yl0jD7AmrvROY33YR5XeaDMQ6n3FP+cxbAYl4DW6nkTzk23rkShHCS0sxegBpCn8p
bEGuuxpxv35aE5/0viZxh4CaIakQSKX9cY5wWoYHIEf8PZASX7VpyBb/jAwTv1Pss52/kTs91PMd
6wAWD6B/07/MumVAIc6Ut145P0SkK+AY9AhboQYiDH62jVqufYaGNv0pjLnJ/fTjy33tNO24eTn7
nqz/140zyAO/PnSNT+lyoQ19wvGOmsPSVlKXl+I6O3nH3/rtHShgiYXfruPO9L5tfppWrx5RyM3H
H+gdAz7D47LIegVHaGQOiHbnx7gRL0u6OhyUJ2EUx9rqBNJ3k2TS6U9yLEjUceyYt54bA9rcVQI+
1/xt4YUbc6fPzZCmuF6LdX/G4qAHK8K4PMKoPjblaaY5FCprg2pMtmtvfzsqpoym4DjEzlDCYk5d
cM06L4CCQHoNmbeX4Q4+c8MoGa14hSlkZynfYiMjl3XoBKIzsN63Bmbf98kO3SFxP0Uek9t9L2cT
PQibNfyTeijlifSfVD6ObOssndq6I5cxNqyLfIs7QaTrffmWrjUOEgOhSr3PtVA70DDSfXAADAB8
VEwr+NpBMIlYzgFdLS3ZeaJdujTQPtZ0B8XqF0b8dDtxxTUnNKTVtNnp6YJJgGBR2AEII1n4lgYp
4dmy814W4k3rLSkPJ6xqacJWhcJLsfpmcoB+LlHAGGr0C62QBVeAt8alktICP7r5bYYx5EFiVKoO
rZR5rxXbzPp+CT5Iyj4SXNjymb0qjW+SYwN6pqgKu/TugfU5vbvxni89B5TsIvu5REhzuoA6aPSw
Ux0Qr+J5ZPW8CocHyiIhELLqwamCw4kDDq1wsQGPOoDeEqOnUf3Hmk/LxyMYSNlPBGZEYSu0pPmV
btWGn6HVkOGcaaEWJugnoPmgAEcPaEKxL3jY/rgiNgeVNYR4wCzt73uxOGhtIV8A07HaVjMrT8B3
A7ndT45MBFkkfbFw6MS9L8hNTsm+ghhhYVl98pVyjUdDkZqg8PiX9MBAEFigjEk+JtvIEE2JiFfs
HihLEAym005wZXivR5Iv9LqjnA1xvVIgrV3U5mTMeT2pF7EFNwGICoIGEm9Hx9hH2FhS/PqG0XRZ
rCnK0C9Y9Ol6F0Cxo2+EhQtvat2Kr2aEXxErmPa8IppkET5nqfUNRD4rdGdg0RYR7sGwU9vbC9YE
VdW0gZQlmJ+0gazDw4OH1rnUWW4LzZjG9MoeqKvu9QuOPvFdxfSHgDzKR+Be3bVeA3dKrkSCK9pI
Ph7MWWsWbHFiyBFIR3O35Cx3T3kW278dPTzhrVZGD51+3DKqYndq6Bv5jSI3m4hqMqZ4fB8su4gh
mIQLJ/Q5HYd013i0hq0Hy17Z5KLWkw69u5zmmINkiUM8ffG6RYDQwkIVdWG+Vk8kz9OkJaKpOrET
sPrPXILGBzJrXMUWVHv3DOvTL9SttAotvJ5BRVHdb0ssw6kg/iwqd8wJEI8DCrSoLlVW3pRuUt/s
DNqGjhOBhr7Cd6ZRNLqXuBrFV6OBg7uZOxHSYw2SHfzs+Y4bLwrodn6gAPa9AS/NJz9IJebKYc/m
U7tEe2VacWCeyXTl6MRkXemxebNsFf7fz6lhzFOIGZ8jDP5QgQIjAu+5ZX3qzTF59fLKY9V/1fNw
TAsp3vv7KsZEE1pw+ZyYFwkY79OxyDrqmZ14ZLETRTaqNvdcN5nyBIgkrn78qiSTJqO4UH5LbTp6
8tDCUxKFSCwmLp7Gcm7XjSy/ysvtw5gSoofqIhPhOBJYaVU22eXSTJlmQKpnEiu65cVj6hFfN67Y
fcoG2LMavw4gKjGhvrd4zyvQZpKtP60wmAyxDvZRDsMBTKL9tvuMfJo8W3tLm/PDlqTjmzZgYfM1
uNhClOvtX7AX9ApZPpCnaYlrHvgWhcscbZHpx6crAFgXErYQGLgqxnsmsJpsunSUb+bsNq5KaDFb
erhaeabC4jAEZLWaZa4WK1iQWAtEIKdzEVgwRsYWQOGdEYqJEuE7S6J2dGlrHmVUpmBaoML5uWX8
fh0mdWRBLTUC92dZjXAkQwnmtpow1LOO9qWho9S51ukxSKn1iFzJZ8kmZMO21zX4Hwz2QCFLL1zq
x6Ihxh7ViBx60qCdU0qIbC8hzZbIn0WChmJNmohpRvKxxXwTByq4dgBB/M/tIQdI2MxJuLmBs97R
QWAvxj+SFMFAO9gLmClVeiO7HtiKxPCCGX6YxGRaF0IficmCpEx1UFsuoRqRDlg/bWm9OZbMgBqL
v/+cOGKJvtxaBzz1N7ajNXWWFyty9catlDdPGr/8iQz81DWSR/XihYZu2Z01snirHWe1RBqrwWLB
AhaktQR5mzB2jZ8n5qh6wUUWvbcTXlWpFX+7h5MS7LhL0ilY8l62AoXgyRw5PLh2CliQtrK8n1mF
1sCNBXowYOt9yqKdg+PiBUQeahDkwcWrCdfWsmAWfiZCCVis9YIJj5KeKP8kuZcFvo/3sawsGyLd
fB8W5ycugMUoNaGX6hGKpPI0H1y6xbwkK8PFP6DshAF1pb4fWxTHNc1+CiEMYl7K1fie4Ze0Xsm6
uOQKLFLUnPObbI181pDgwWkQjZiVe95T6w94Nmhu6W9JgrFa6lXZ4mKmzTESkqhlJ2cKx6c4zKQM
ZLw25gNqTMVsG/6PQYUQsoa8uopFOFd0+HpfjGQ8skgB3d68/r39Ar78jeqW7ChkVCRF9s8fssd0
yP5IDJwZ5gAavMoQXuv0d2ttWKlRRaby8u4Z3uPd552NeUoAy1s7LtfPj0FV4dU5OgdxD3sIJTQ/
5+i3ivQp6XtlqUj0P/BlvVyvn11ePrwVgJLXZ/JuhlbsugddJTxQV+Yr/pk/7pgrJkYxQ5vQ8i0j
cM/9NLmNdi+sHd53eO+2sUnfnFnAK82XZztOo4Y8dNVNyHgf8YENsebtVaiqKNc4l1p7YKX2GYNC
h/37viksqTGPe3V62kXrQeBxcf1RQlqb7+41BgFUyeU9G4qq7KJsMdJYe3vSqi44fdpF4tur/oaq
Vv2ldkKwaUX3kPRf8xMaLCKo1jcak9espUYEXAOp19g2P0XKkP8y6IkcAQI8VJ2EAq8CqQMQifKk
780hEmQPCHUKRjPGE2/xChS9ZQ7zlF8WAzfLMk1Q+dAn2Gh44e4btMJu4ATYjdYaX8a2nDIQjQlf
Iu6+nQcm9O+yhJEhxEa8gMG9ev5dpCHf6zUbKehgr0fGwPeVl3xNNrRQ9TYXCiP5A0ba9hd0+oTd
i2s/KeA89U2dYPtyEZRCcIvCu2YuX8ZMZpFkoshYYuzl0bDpAk9Cw0Kg40fyUChKQz7YGCOeNmnt
wZ5loOqnenTkVv+jnOSsu17q0UteynatFZTOQdsA5P9qQG2rAxQlW7sXEsT0ItPYqhC6CfiTvP4p
wNDOK0RUMIiGN3eWeBVbI59guOQIMEvcvFjhKkFGF67B3jdGg69IvsMB0kpoADMkyv4PJ/b5WWJT
ZQCZvH6YjFdt6CU6UiBm1t6773dMXR7WDorQRA752o6OWi5A7HOwRPuJ8gUdERWZeNih5UCi13/Q
UB2zxedFvj7EcGN/oYlMDDB23sZ0qhBHnQu94exfGddr+dIxL+LtjQRUzRN5v8TtSrJq9uQpb+Yd
bi3jJlufOtAhOUTD++yEIv7vzaTQOiyJbsy3vUWXyGum8jA1DAosW/AQrdiBJc9Xw7AyNqP7j7Yn
SN9MkGWDMyw0Oh30APMi6gqA8Ix8lEW+lGxMPh8ISF9i6WyHjveO30n8iuHh66fw+ZEocLXgAzfx
3lk9RDkq1ijr+s60AuK26iLlU8iPV51sN4SxaOGAtQCewfRmDdIRL1pC2m5R9V5v4t66i3oudt9v
T07qYSUdFrVCPjdIVicWs+YEk91fVPxnYA9TDYmna/wTQyVCiF9CqzZlwNwfieaLbl0dK1cuqRVX
OGCN7NJT+0P0ulGD0hwH+n6uvv0iA+AB5tsJU09ofuPxD7ookfaHl+tNpqj0xGtDYd1Kq9gfDz12
tc9JTBwucLP5VJrZ+5zRXn5DboUpttQcNJvM9Idi62p9l2mtpRnEnuO3tGMUwHOXKEhzakncSiHR
q8OW1Ng6G1IU+sEbKAeGYTAqr6cRh59YqwKpfNXhqOPhEI2yHJB/OZiEiO8fVyEwgWjVgrpYhYvp
LlGInnrrs6cMXIz1uyM7yCFE9w0Aw0rJ9npThoBmC5mkBnaZieiBrcHRUdxXanPa/Rh3o/5fJ3kM
oR7tT76wnp65te+1dd0aS9BKSW15pVSUjaKlRZeBanNvY9iHD+oUQEsLnsqfco6EiSPjkyG9wCYl
6csSN3Uw27yNMQbYpXlIiEB/nRWihs6Tl1/FXJfh4kZnkjSHFYXi48k67PGJVqnIammP04Y1hv0N
VTHn5p/LSCthViP792/lQfIzLzGf4DwcOcvvYmXap9MqjBMnp7ln1i3+zHr2dcirZBiJs6BzT1KH
+p/JAUWWJDx/aSHVqTHUlf8uPzjEdqigI9E56RD//AupaDSmd3s7w01AvlKbtxqyT3RCtu6kkygg
UnW+1dn/zV2wP2jo1RaGjtlZ/i2nkq17U/zk05AUg0KpTkpojXcsWREeUgQ60VLUVmwojogztrF8
icTCvNcNNE00JcRd9QCMfWupV69O9wNTaCo5tWBkHiMTY/GgIez3Ewe+DQnlaOaUe7GRqxxcr/14
6wRyG10ke82IluVNoW4RjGI+h0icikCRxnxKhcjz4VISLNWn/9PSfVPdNbYkVwszPq8T6yHm3KG9
yA8jiS00UvWfMwjAc2wOe1MyKfsK+ifOCWtrSx4oLQuPLFSacpSykZ0rKiU6zNDuHHFA0hl7S3h8
dm5Au9rP9rYaVOUhUWUELmFeJXBeeX/wZw7tDEYe1erU9Hr6krUYc25iLT4QoLP0jO2nSGtkeQDh
oItql6tP2erVQE90/j9Q2gSRPB43K1gj14tbpyNdGCM9eEKxD0Gin36bjAiPW++2Y+ZNCHofdJIl
ERKmo/+1O8E2honviTrDcbZeZvWcJQ2LaVz+daSYYWJR0QoU4pUJQT9RsY1ZEm3W4Cu5Hg5flwMR
ETc3LXsBN2WSP7wlwd0UYcqwuB08V48rcAtDpM6qY+Q7UZdIOpVYK7cgcyF10H61T2x2HBi45iox
y69PypbZGrvICXId+8w/vjgVVebOGsWqbAiT8TfQ0p7of42hBxA2MdTZCgdZ1WewtjPEA4+GfD+0
7aO0YYCKAY5L/rTaRWtRJNxk97z2JeBoyYdrHeb3dbqBG8M8drHFHwhyLssV+Nd0Whtj3oWVu3NW
CoNRC6x8PhXPaFNsaTPvtLCDP8J5zgDPY3+yPK3xGyYimPMU3pHtY4RHcFmTlGj2p+/FIx9AQW1E
eHC/IBvHi9oS04DAz+LczD0bC2I31Z6i3TzrIKhIUjFVgRBwVhiFX0RTT4J+dmGVlQUtiS19ajup
jxO35nfkxFPkENflyRaCwKGTSlM2QPjsqOyeYdtsm1ld9wXEmeHfDFt6xwlm6wGv3CfkXzMV+a77
VUeE8NMk6atk5OgIDIPIG0nNFK4PJeW3wa3/YlzMfrkRORip1eEMOWLJchIcEOoQvXpMwmVEgoVl
igH9JV2n2HGZ2j/R1KTg39IRdE7wjSViVp9O2eop0ZrpwCBFe9ua4sQvtTsdkPx9DRNMmfutfgO/
X+aWf3rov00vClJ3KdC7EGpJ1WnLLrFeCer72b+YioDj+ZgQo3aKrkxi+E5tXAhIkXRiuDHzi/y2
NYs90ln6P/51XA0TLiIdUWdx6WmFMC8QwVEmj4eIVZ0FIydusQS9gfcOoP35m1d/8+sG8lENwEXP
vOF3NkBIOY6BM+HLqJuSCRmFesYF6CqjfsDoqab/kFv1mija+CDHUkz7qDD1S7wGFmXu72LEN0ED
cfn3MWNezsWhD9MJT4un8Y8ynZa0ksNdm9V69DW6HYBqdNts/R6CBenm9Ewyg7fg5BHb8wtuMPqd
zztabWbwqT7E/+aaq/2QafWf6x+dsYSnJlSh9etJ+pap/Whysyil3C2o+W3nJPZ1XVrK4uI3D6mu
qt12KVJVs0Pa1SzOYammwo7kzj7Bus2NtH9+lkbT5MC2l5Uy/XzZQyqJJp6Ybf7ON0/DvRoqe2/I
yimsNkFPSOmONcnZD3nnVvQnUNF+wBIrQY7perLxIn1g3HhCAsLJuJmYuhq8btAa1kQ00LhM7D8u
mAuGp2ZRvtnbNiAmI0Z/VyRidBiqYUqj4myyf1ry7y55w6je3EAXoW+l40hj7mC4/eANdRt5sGZh
juNOl4IJwe8GAqwsbElMqMiaDiTSrc/83FlBivDVYZlMU8V1CDPSZc+jzrvluJtpAljKsWJnJQP8
Vv2g8dN8Fq+0Zk3Xsckxi0UaPoD7M5WQNs9d7CFG0SD/AQ7PGHAd4bStMvqLravQNDj4McRAauxN
GpbMOswrizIxD/hplQY/8SjcgN8nuPIx5IFiXhhfbRj9hD12AsS1yFJ0HLausbVb8Czg5OZC1h8y
XyUuy76WqaCw2fbovZUqEt2pvLLOondIgDWZvEaG3LkOiO5brsDJcp2GHNJ2udDF4SmowxxOGhOn
j/OTLk17k5cNaNtghS0hagwJqdlGJvgf8+hPR1r/sGZU0R2IJpzktbSWOQQ/dL5Fxm6MZ2FpNlv9
NpwcOzB06jTg55JLPXhuZpNFNTywnejbEvbvPhHZP4stvRwHEqJVjmlArWM6LI1VkqDNrstacOju
OHdXw2yVWQY4tYaQ58omwTVMVW3dvLkFCbrH5O41FDqGBiG26/XGFlTVZFuFnT0IpPrrQZIx/hHf
UvRuDo+NJJY3/KLdD6z843gVoz557AMj8zz+t0jvaQSg61MQIIGuaDrzUAvLXwDsEzdCRMjmFLsM
ITQZm5dsSiL6l4Lj/o7VFP07YEkoZcHEjo9XAqF34VfKuPLb3svTxIqJIYNMZeQs6YcbCLHDskqS
7YkvmuRrPwekoeQVJUEiu1HuNPDIITUievFXegta7/8EiXqxwyV99VCDi13qFYMK7jgz2gdhjWEZ
U32AAE/yRgAJweyDppaoUo0PfoVxHL3Fsj4opepZVQdM/oWQQZhxF6JQwFUCXmGECehmbDwBdg3G
QXvC5jrLgh5xX/VHZ/Ap1PG0xilGNb39gKSiZtwaMC3cI/1Rn4fCDhFVPwOvgyWExpmIUq7fWCKG
BYS7C3y1vDHxVR9+9MriLcjmmuKgxwdL5rc17632azK2VWwgMiM3VxZJet0KX+ytc+2QemqNKh2k
eaLS2DRr/1sOJnBXrXZ66AK/GHKRH49vAp1A+vGVHW4aJFPMq5LWqM4ff0cT36dUX6S/ZPs+v3Ml
NS2jKmfcI2CE6NftL2KmY7w7jJ0NYfmL6LBetqPGZxhCcVtZvj/50PrG0L2sP87/njxm5MXuzgz2
vERiiYWyMaD641RWcBCrqMZYPsBAnSn4L6F7UJq4pyi/wuBOvz84FK+b1qZZZRdGdfxRSgN8tLwY
7Gt7EeI+4nxqH86lGA79eN5KS3s5vpfpU32s6MkT/xtjATBriz6Y75SM3N+ULPaC7ig6Vu8Y+zxj
Q20vLStSX3LpyKQr2LSCVIUJy+eO5hci/s0MgI/CgHJExnktJN6KAH/u4ZdThtlrI/B3lgkIjcXw
QysLbGyhn8fC3bu14WCsbUCWNTQhcWlHIZlQ0VF8yOPkh9DbdtI9pr/49A5rBMMJuRT644PSMoro
5we3zqAbH26PR2+ponpcJwRYU2hJiDmfwC0WeHaBTC3psOj7/sxYesVCkutEBkqvZhcMSGZN3su2
TRwNsi20l+uGSLdY4jrEAhDqw9+Oqw+sf0ZxzHeN2MPSiPnONnGNVs9G4ChvBB62N9vF3kUq/lbO
SqLK5yd0IskbjBl/8vm4L9B5S4ftl4veVH6BdStPxbbdbv/126vB5CUVG1QkqEabIOmcqZ4oOwym
ubnxwFYxQcyMq/klwmRU2AHdHQ+QRLvPHcN7YmhNg3isC6dR7L9ET78fqH3VSZYzCAWvx5AMUecY
p4QVpk+v0NsuIPk5iRg2h7tcfFzV+ZliSzikT1M1evSSR2N0zut+xyo+V+znBMw5JZoiRUZgmunn
3jJyqVwMdUn8GQ2QF1WL5Cc1RVYRjXOjK+d74Oxqo1wddMyoauSg5EB91oDVU39ITy5HwHa1tLwR
h7+YwKzi4b9NRwwKCIw/Od1l4qjF4OVjO3tp3iURphCS20zrjPyd9FSXX8brIce/97MahayyueoG
tpmT26OI3H076llG8o6T7N8pcZ6WInLf+gAHs9FUzEDQiH+CaIXckLopl1bOEuA64u1dwv+KEpZ7
hLVMpJ+lxuDu7yxxCU8YEYePkODerHUyscZIQm8q+Om9vgQz/EZgEMEYdFgxj9pMPoqTmN596BYg
H2SNpJA5AvmlDhmvshk+a3KWb6sMYe0lLeT5PWz4EJ75gkDETBRO5PWAdVvQ17FAzHC6fy6PrhWC
RoTYlzwrWuc9xJf0a9WIE2V/W/NAccCFiOS27Xx9++eOygYDyB7vvreAFhPCrrQBhEwII2/nXR3T
azs0oDsG140q9pvvv8asGeSzkswBLCzh0zOj7USTxv94wnJq0zF420tQn6N8vXbG5QSIDcAlMbMy
EhIF/WQRXlWLesifc0Iw3THpEPzxDkvCaN1nudP/t2W2cPu1U7oA5D1YPth6o1L6XBu5jqIl0RqY
GYmeJjw4vSnEKwsK92YmIL+ZrN4CuvqlpM7iVhEJlTMkrVvGw2uN6n8P9ID8pH4YygYJM1g1Zojk
I6zHaupRrlwlswITheBqXXASylYfnKuwkgttfYjxbYPIbXPtSkg4YKhtJGVwFkQx6DgGvurt5KZv
5LmpEbDN58ZSDbUw7XFW4DuWK+1ZEv5eijBb3C95A8xwtMPLonOJLFzmAaOc3YxeLzHbGV7VNJcY
BfaPfTbbHyM/fVIjGKo1TwiSFBGZlyI5vBFPei3YKDXZYaAjNorkJMk9ThFvU1CJhoQPND9frvNH
ENP96SYdkfGEnmN0jI03py0zLYYpcYAz3c2O+giNV/ZBdZmxr/AbrmsMy0v9YhvEqxTc8FWJNbWQ
sVCyVTsL74WcEIOyZZgY5GLNPA516kOj7YhYo5e/yxJUb66cfW82EZQi/+livEGyGN4vCUzjj655
uQN8iQ3aJnIa7qSsscYAHfsT+/OjHBmGMBXl4nKWB6bHleu4STQMOx+O1cBgaBtQ8TUHgQ3dkd0t
6jDXvA9fVZajVBXjT5WMWeuEI7v4Y+uPTa2K3aeQI7KUFY9LXfQnW3CnVYtCRpzuZLCfx/L5Dlg7
VJkMsNnAgVBWq/Nsa89xcoHUQkFVAyMk4WUWSjK6i2eo8i2/tCMwTFXcKBCmq/tSqA7W3YhMBADP
zkYcGm4wfxng6nT2l4AViBgPkOxoajuc/8ev70l3O0T7UC8ydEXc+LDoKOQIsow8dfDIzJ1D49mU
32UEbb4n5m5y1U8Utd7VUyix/265OwumV/ugOfoI9o21/1sxPtW5cgbsV2VZlPRboJJHyK9UHzx1
QvzHkgom7OrBrPTu44ndVZY7WhkWmqvGnh5aW/tQCnU4/Br+2xGRb2EvY2pc6iDd7e433NfIiVr0
r1B5X85U5oKJ0NFmDk0yFp2TqPUzigr3J3qt6is4cxPE7ApcxDBqWihlUuSgoY4vHzbSmrjYpbQt
I2eJQqpGJyWQNuBeTThgm68yxrMtrigDJbXEW1jRZpzY7RQmE3HVwsvOQLlmELsXO/IvVU2MVKwP
5hHMy8Cc5QS6js29x1T6o6St1iCS5KkirmDcbKIGXAHLNZEbE/GDgpig4EqUUxndYgSD6wYgi5Vs
T6dzjvWCAgYblKvhhgJ0/3/4oX7JqtpBFrksReAN/gGeh26aWK9MUHak7aDkdkh6oWQy2NPDmGTW
OyuVItTvpyI+/hp9DL6a3hGfEtWACjIRkBFFtvK1GaBmVRkUw34o4/DbJ5jsb9cmZbf73EDKSnGt
EnJHeVniVyFdK1O/pn2W2Vs+94jQUqnoclIXL6pn6aFIOEtcM1GvuBSlHsul3Ql7tZxhspMVp/AT
9PsTG779H7WA6cznD8px76yOL1Dd6L0F9xSqOWyXTqMi6pbQ1eboUcfLxlIodvNrjvmNd7tg1Sy0
nhAuwJ8Ul5iZY6SbwaTcRRpfXxbaiRjraJdAvK2whKpN4iz1t8DAz1iCnB8FUQaLxEm+nwnGWAVi
GfJcgmjuAKQmQXoYssWafdP0dHkvG+6xEm9x8PLjtosBxfPRCzZShbkGjeGzFhRWLWlK6UuqtQMt
Tfz/uFkfrteEUHi/8OE6Q9A2bvEFYIXVMwpjoOvsEzE0FiA2YtknZCdpMhSdYV3zR3cQFMPcLwaJ
3mG3yjSokViXlEmfvSFSJogYH+F4YaDNvFl5Sz6zjvnCeO3nq88TPyBd2EhCSC+IbX+rqqXc9Xbt
Yt0Bg/5AutWRlyZPENgnkNc0mPlm9tFdhX7kIO3oJoERo4HxK1tFMjtl+XW9pPkYZ9ilwxfy9cDl
gBGL3EQDU6Zm1u7i9la/JxFi35m80KJbyL4kXByq80+xATa9HYQ6bZMczjzvdbpRqI0DDOJWuVq3
BD3C8elojgAzaUDYHIt40VApcLnQ5qJPKfAy0hSm0lTj7vJAXY2ibF/Nwbw3mOozMWF3qq+UVyy2
2Nqi0p+QmQ57K1KGkctMw2N+6Kp5mifQP+AxtytfGCtVm7lE/UW2kBom/x1qM5fV+dXCTT+0Ymxt
SLbjtN948MLPSSNhX9vBLGseXdnjDYFQGs60yFhY6fC7zMJdMnnVO0xybVfSV35gq2kFE+YlqOOc
VWjqqNd3GPYX2dtJCDaR628urTE8AWSPw7qiDYy5HZe70N4ykJyOrYNQuNB9+9yQVEHBE3/tcaO5
0Fx2I3cirLKZDyVn6vHNW0wVlskhBvIHaybM256YSpGuAYPhFm/bJx6fPnv021RCTv5+Pn9LAuGH
jJBNswVOBgmIIlPcyvjpyXPM7nhItPvDIPJTBa8OwWzha9EK/NM1/6IoWniqqZL4Xani5517GRpg
0umc7QMCfrXHovxvf3NVL7JnOtno3QcSI5AWGsX3/INqRyjTh9yUBRUSHDTmgHWpROOgkyS4ojHv
+p9pAKLF9JoJg7NBOP/4f0t4IE3wVImYEYpwwxTcHZTNzeuOq5MhRVafG/bbz9etrlwvwezB9ePK
GQAuQmPd9I0S8jWmAtrVoxeienT65/WJDOTc+Pq1ZnEzn1mtOmMhh3J3Q3jU6eMaTuUlzgPpH0wo
pFT4X3Hg+QbQHwgtiuswt/1OA4LvNWJ+MkGqsLyEdCbDLyAwc9tt5OIfkzs632yZIOxUj3Zu8J+x
TDn+F3WxXPYcjUgYhv7IfyAM+oejfD0GwEwCGzlQ754qPFgVkf9fNe9a4zOs+jSnSKi2YsDQxzoz
BZkVQ1lEA937fP4FtlMDXDt+LLhYDBBW5R8eL8Zbm9hfEqJrdzf88lMyo/EMqGmtz7TLxhWqGPCO
tM+nxytjyBpzyCvobIDPw5FLEv08mb2s4UM/fra4ooUufSy+G50RfSVLb6Mzr64ZFQ/SQyl0ukxG
+a7cPHAMajRSp6WotX6GmBTkMbfdn8ZXSmdGliptc0UcQyiZhtccOOwM8ECw08WVIPKDYIQQsWd0
3VsRej4KIsVx5KOYKXV6GYMczP5c4uolamlJHWncsjkqVTWY8sHNRe7shAQSnbCDgu6E7RYFWgff
en1AJIzUTiDcH6OSFvCqtEOM9Ou95qkFT3UklEiUsG0XtFSIColwrNi4ES4+adpH33AamRyhqhXn
thm6Ose6BcGefSXOSe1/O2q/BddSYOdYdKZAM80A8etSM8MKaI3e3kCy7QUVyYom7570uQNWRNrR
XiMCXe4yfrqaOIXn4vws+7naR7JpKhIoef1xjYaKaVRI2mXwbHFSsT+2VZ8xiQzkuSl0OGFtVnWK
nsNKbLb++QiPjGVC+RJO+3yGQnt4g9YoNehZqoPpH1fG5I5I36Z5e3WHvTW3Ml3TxoBqHZYj8k0w
PfbquKR6fz37FnTI1BXAGzN7cz0wb7Qpxyurf2yzmBxhZViGQsAZjgKyQj8/Mq/Env4Xc3dSztUs
CnDjzGBbr0VZLbedyzmLQfXkW055MYCKWHe7EGlNNloa6BDbVYFNrvuRsoPLIFn7YyEe9B4IrFiy
puIXZWA6djwEEf01drRfwTcNeDaSgGiiFquBbqIb/tBjc8BYEjrBjLFZ02W2dQ+m/S9jwwgBKqx4
519Q+slp6WaODTqSvcJE1ltXNwtuHBf/1jqOQlcubYyy3qN9kF7voYuKowOsVKtBS63DkEm5ldKN
0SF2RXHMjgqP4ccXQ0Aqo8LCy+pTOKG8s2dRsN3PnMTlUx7BJB7XwrsZ64TFiVJpCel5TJOZluk9
Da84fM6a9BW9OBDB4VSPcLXdBTcM60llTpVsSfEI0RuGc0nr4aBPNYgjmgFE8VwE79yAaByM+GSi
Otl1DlUy2DsInrLRO/zo0uitCiDWQsAJGW9Q7AnVA0dNGOpvochQit4cc3ThU9bSnHIVQK0txHo5
9AQO70Lnk/4ENYSeWck5BwoCmozABke8qztBeRkkSNCn8nUz/s48m87RSxAL4JM6MVmMjHXbCLXz
ngX2WMsV5CAZqvkQwTfmehU04KExcaUJDIe130zY/34RRSB9bx6+7Rs0WCVNHUUNML25ywefxRRF
JbjDD9UszCuOSQHrzBq/aIBoejh4bBvf2w4PZjxFC0OYXRhOuL/uzZ0L/B7QIiwIL6UR4li3NpY3
+ICo647jfomUiseueCvcoA1FpjFKqSxXilKrhPWSuQ/S6cuosTh/ervZ63d5Oyxn+/ph0KEVvy1I
wkLowA7Ax+6768l6mwqZ9fQcXe9Gpp1EUgIQCCR6tHj0RJeF2ebw2TaSmQZY4DASifgOTyQk6UxQ
ZUJbhchbAz5Ihy5Bfix3Cq3uAPTtE9M5dF7mMYMtokGVfA3HZtKeNjywO80HqPxytkN7LIThSLub
zYPDFpmYEd1GnTBQwGJb9zM3sE8GgSl/qpeaamwBqg5MzaEfP2iPICxEcEkourOseHS4cD8l4k6U
J+wNWCV94A2cHy0RVRn57gWj8orQPK6B3eY/dOrXZEVvufgtnjBnAca3GqqMSWlKWE56qqiIsq3Y
AButIVuzx1okZwK0Y9eoJx6rvnYUQN/bAg411gXfE1e8NbXy8hbEL9LPkBnylQhIRIama8tJAKu1
1WjlN9RrVIB2XspbLf6fKj0s3feiwBoqAksdElUgfdRogXN9sDQkXI7UjGDiKQLByo8OyIUArdry
UHNbt45wirm0HCzPd6LWd5SZfcuUQV/JOJewOxlhhTSjlUdm8Ry4seHEkNk9EBc+8ToyN3+OJYId
sQuIb1uqy3QgcdrhuDX8u6I169GFRCBiqg12Fglkq/V8jaYEDcbOqQtuZZqmUM/EvSmCKKDMyWRF
ZUDEkoS8b3xFVa3A25Rtf8iP+yNJ0cfoznGNNIc/zkk5NUvCFNolC9xsBtw65mSBCwSR9opfb3+E
gAxtzHUWIL68x8emti/WDqqP354OB48GgzI2Zjoco4B7JnOo+zAkmc3H19rddo6wjycFhVm1aCAR
jIgoQNkdKFy7OizjD3ZLgoCOz1hMzwsUZ2rHPVoj7tvOez7E/DHLHrFtwC8hMxtAc8lpr9W/kdcJ
l8uCWEsk04jYKzXlaqwB/6IgWrPrkzshK5KX7xSryPWMOM32qBCpnBa3QrCLF9MTcUYSWCz+c0wo
TR+L4pmVj45jEaLHJDWppwn/2qPDGsZhqYMOw3kip6uIkND9mDi5VT0zrlv4isEcLBkpybUkpUcQ
/Mw0XpK+BDX+AbtbGXs+H/nZ8qw3hRlUmk4CEfE/CF2CNXyH9M56yTDCMSCZUYyjD2SmD5F2gJRv
GNO8OCirbM/lWbMX/FoKSMQOEHDq82OK50AD68NrcOFokYKPv+++vilC6dU5tSV87QkoJjp8GdeB
yFRQRW8JZJVGvLjd3xKRnRB2qN56jElTuUBgB8Xym2KWd0uw7EIvAzeYtiedQHNuKAGpTzvry1Aw
Y6pRtkfoXJMJC2YktXXBPaJci5rH7dc8OcRtzrQK3UeNV13R5GS4I+zWgDXJ1c3aMl+7wYe6k4ez
AvM4D1Bw5W9uRh2B1rALkQdz5SGSGAFKRVlUuzq2mMSKzXFVgtIcxWlmeaqZR/BIwvYUP1UU9tUS
nVxdCd5a9vndWdpHUMAMRlZEi3Ls92XzR/PLNxfyyn7GyEe+w6grP8MCEiQUd35JSMYn2x1UBFdp
w8SyIZvx3MsdB9AwVnkp9bzMe1oUd8Q+4zeCAHlXuVN7Q4O59H+wTB0rI5dQtKZzUzZnTqWiRivD
q4R5GMcUMhiLhcOWsS/eevCOn7UHs+hGIAPikgvM4GqCp1XgQ5A2WH1DkEmZZrgZe84iYaJQBh8p
BsSLA1Rm3kOUc7mkgH1qxSyRy4TcdFhmGKpNMbT3HzOahdWBUYMN6qDVxoCX4dqcgDQe7WD4nUS4
8A/qQ/CtUNbqEnY7L7VoNjofn8UUQGgk4wDVVKh1HmXjr6LSBGsihDOMN3u8DatKBhBRHyE1NPYJ
JueuOYHh2xPs6TkXa9QrObjtf5OsjIP1DOBNQUPrB2tPWAuLNBI6I9lWpMfmpyE1/BU3ZE6Lm8BS
nJX42e4O92spJ6mlns/LsCTcjrY+0oCPH4QNEb3lEyEa3GrRAfb/ygdmQ2rLb/fYhIJ/KimJZr48
5x0DbIfkzwv1HqMpDQOohy8NX8jrMuJaL+fIMdVvl0V/k4XTs53n9gb2ehuSqqz5lPcAiz8eBs5x
Q0qgGWtl99uzlDX+VsvD1jeNSPB3ZIsQY+vhveXLag7+gSZAY8PTM1aRH58qkCup/MWmAOKbgIjn
rbUrU876PTo15uapXJm+sANjCtKsm4qh7Yb8mhY2RQn9nLh2X0H0HxlPA8L8AYakJo8xgwA404W1
XEGIknWl/UOWGYrwnHHCPe8gbFzbCzH/d5mweTI8rHXhUh1+/IYyKva4+zS4AWB7wLX5f+XU+C2a
VkXSuHc7juFwAyzGfMjJN+oL5trbl1KnAVEiO/m1LdLvVVC6qj6MFlFRbxaprem+das3xYZJzYtx
fJb9WD2tk0LyvDsDin1F9kyhXgAo1e5LuUmv2cp4P3gLdjkO6ch/tacXAh9ukg3MrSIwTa34mf6j
/bizRgu9YNhRHWenlJxTl78sdemwUspHTKtqvFwb+7aEVH/Fa+My2MLi7DW3IqmecCexlE9V0pB1
nUBHL7/eguCb3uZK5dw9M+NFRybVJQKAJ3rvjlbKq0mDDiIGGMtUatmGNGxqD94LM5EGysjo+f4s
Pg3sBjfcrtCMUTqRE8V8zl+CD18P1dWDt+0joq5U4WD245rUuGD/TGdsblFQuoRi5omB/TxvSgTC
OjUj7XqSQKof5QGrqPdG9WxQvzsayh8AlF5azoqynyDzC3XwfMd/r0uwvtFQFxgbcJpx3U+MhMHR
zTNG1Jm4rqJHionRJJ3/ws4jtVHcqOX4ZE3FoX54orTAo6GWO/+DndrfvemhPFsQqndowOzMu9mt
HlUHB+xTXIhFi6boXuP/hNzvwnk1XpVnq7y11uGL0ZNdx64JX7aSD/fj6VsKmVB1lMRELtydYvn+
4zIU6Z1TIsjg4iB9A8YD7Y+hSMI2MH67RQFbr2AtjMzIWFGUtPsQbRkt+FB7dMVG647R5dVjWQOc
9zu355zA+dHm7iOwD2n8O9ZK4IjNjLJH82y4TqCpAURKBbYMYxmCFNqOUspJK2gbQcZB5fHjGvLf
M4V5BX0oV3NfKzneDhVVrQBE0VqsIhvUydyr+NAV0g9Pd0KYSy9/8cGDlBgax64pubqRruZW/581
/ZDaEqiCmzeBd/sCjLkvBvdNQX/Oy5Obf0IhOKXoyagNYrnuqm6TtCWTIGD4hE4h/PQc0oBeDLwB
NYAA0yp53V+8ZX/HJxEJhLO9FAx+Ty/0aYPl/Sj8tM9AAYIuZ8bvjwk2jKxkefb98C6XWgPAN7Qm
rvg1QfhgdFhc7YAK6EqCeHScl6RDmZ1onN9jFSuWy8C+eXz08+tDJn2dVqq8N/QTa+7CbuFQvW5J
WlqFhoT5UYVcFA3j2aWw6zhzN0YHcqjmsHolzCSbNNpW/icg5ze/lFDwOQ7RuwJvzdCKc5kIvwwE
7UCMcOcnI/DoDcqf5WTtfoW4ZM70lnB2fswghP3u7RMu31js6hjvMYBaVZ6+aKV6uIdxdd/Y1+J5
HjvRij5jKBPzK3CK7Eb1+JhQak/xDJ6hAYAeNtF6BZSeHKj1vr1xdDzMyCMYV2oXJVVwh74HIDmI
R/AOwDOmP2urK/dONvnyDpTJWqcnRk1YrMm5+cv3qKVIf0vwUUJ/34BBaqsm+GuODhnFhravpd75
CuYI2d8li36OCQB41HE7U08dz6TShx9asHfu7o3kbe5f2VX95NIu5UZ+3PEKTKv71G/ucO4cOEcD
0ErUdWB6ts07uZboRaWElFnusIH67GDsXeSCJBYfEuZqL24QiDxwh+QUV1CDZyOsnFcOV7DpuZlq
mDY4hB4IDpnxbwW5D2siHzPu4yV6AX464uRYWJaW+3if2A9fjCU1uPo86A9yBINhoGQhDMSYq+xI
IzAHO7ErSe+MEtxcoC10kMBE7Zntr4eLaSS39CnLo3BTMwRxeQ4Ep/yfRiYtgXZni9hPzIraHw3N
ods0Vtl2I4pR+Rkt5S7cxyyAMYCyelI8A8/ijJEnOjcq/0ZOhP2wS330jMHRZOJ3qOZ4rK+NHVdn
gZh4wrVsXL37/KQzg3u+RJr+oOmONM06Fr4hTJWQ2gGTt/DEN0riMCcnJduHkCxd2xeLvxF9y+IT
DUUNmDMHAzPCY63vNlUTr6TkZ2KCesgMB4/jQ/pj/+BIAusSB9Uw8VoLKGV8PwE9rjY2IGZasknY
nDR0ZETn9Iah7K1+ankpEj0yy0URUuCZ1yafuTvsLYHXD/S58jyS3JpCt3z879+6mGjfW6ZjOU09
XDR0kpecVCO4NEYq+AEGFgohzAQrfOA5icPbYzr37stjEN9Wgn3CiUofNsAIKV5bMu0nk+eSgtGk
0yqkqUiikEJ8t/0Sb8PrpPql2i5kEV52ZNj34fN25+Z39nmmQ4J1nsLTLMupG3DxVp1lRxuIaNRh
ajKhOtD3KoUJBrPriB1B8nS5aegl+kNjFiqUoKr2WQs9UZRnUSgil3SBKPW+TIaqRie3/daGxEYF
GQzPLWPX0k+jH5MnsN+UMBXzB9aHMRkUiw/hh1luVSpWD+GY2QaYqr2mxAA/Ik2p9ROVkUNyEsUp
rDyGWsnwRTLrw99wLSWnOBYrohx0gIyqBvOOeORHz43ABgpzK8wnTdnPAUi8xA7rh0rGCKn5hQMo
1n7dgBdKwGbbZmEha0sFGZrxdg0NFazW1t9Lrt5WSogLWoT+ZK+GLmvkldWTOry8d0pU7dA2gUIo
fyjflaQ3iSeZEcF9zJGeuxJRKN6PumWAcsGKBwtsK6rtlJpFVTuY6WY1QDaxeSfDEtZHgNMGT+RM
vY6kileqmemELWWX8mRpb0cK5ITd83wdRoSDVaBh7YonwYjra1/km4pjTbdf3P0QXHSGejtXV7ks
A75yVTM7pNrO64RgLDSR1cFLdX/J39U0+OG3+jcx0vn/nOpHFPjIuQjVp/+v/93bwff3jJr2RKCP
dotSEKxVL3PiUpRds0rGZF4MrvSVwPW2VrIZkSqu58bbsu8mV8GiiHULCYnrv6NWYq4JzLOHNJh4
cqn4X0YZAhghxXszNyfX7XzwOdmRVjErkUEjAehUteaR9hKhgm68pZSnPzeby8UxDsOIIDSK67PY
ogkFdGPpNTLcUCuz+Y1ELlVOQFOv33CIXvTBXoa7cavYiHGyN8BZc+/UmldNOviHcZbIW+z6lZDL
JyN+l6UNN1VxalRTa1LuOmJ+RHm4OCnFPxJ9mmnt1s5foihz0Mul8USlJpcGFNutjTMFQ17Z/EAA
nz5ADmUWFoZ/1oh6CBuf/m5aWftCfT2nZXo0rm2IWplwcvo/qQGi8rlg0WnF8GHrCAQvhpHF9F7N
7/CVIpheOcMMOShh90CMy1F9YvsI6jR8NVYfhuKvHzkTvnwJ9OUyWktYP5lRfJTcShGKZNOecOUn
3FThvTudm5x54HvY+MaTIoZTbSgk5u7f8IbiN9uz0npSZxcCoPkU36DEBokeQOfb5U3JvmJAbLxH
Ev3gTgBEsm6YD89U47yRxrBopEiiF8qUt5Yg+s7S7VpJln5A3TJFSNC7C2ggoZ8QTN9w50gRtsXf
USFUzhWyxXI90NGlpeKnVmTETW1g3jHoE5q+lHLKPT3RC3OA9vn2ahLmRc+yAGQaYtLnyK+2tqwA
wwx1L99/tck+EnW+4m1w1pe5268+wOca4/fEgRXbXguLCKC8kRrEcGKEVeFFXszUB1cOOwvltT36
PKrQ2kpsbNgxSD5NGDCM76D0zlHQVbKmfkg1nA5KAHUV9uU5dP6rP4q4/Lsco9lcMp/JxMVgw7Ip
hdcqtLiI5rpgXYXIxy1/XPg+f2WAft4B2oKCBOvzSO0QSZ2jgpa1un6+9YITbCa36VkM0c5I9zW7
MohmegTJDXEGDhHaqROQIr/I4QNlRM2GoH/uUagxzQC1w16d5QvG6P3qf95dAogrU4+71lVLFHRu
434Kj6zmH6TpU3vNJ40v17h6kqKE+Anz05mgVbhPqqhgaRnT6n2Lu19IH7xUDKkennH/6G8isqI1
LK2wv2UWVrXrC/smDc2otwbxv5/RmStRYcqYP9IC0OCdJJHDIyIZ2Mbz0O6O9UfA6fc0KnBQu42E
avFgkm2fg3Cyo/QtkTWOxMsxm9EGv4hH59uS38VC96ZHQ0AnAAmkKcrHWBwrDvQSJhr6eAZW84ad
qzsvXQwdT228V7zaTAivaXR0vMWMA36jO5ARSpCCDeMkpBtCDtPS0C1y0xHSWT6/+DfgEFYm9HOY
oDo4dcV6zncD1Lk1YaiqYDwU+t6KGgBzZXRCnbRugCGQZ9HJDDT8vaf4JlmNsWyKwm8fgv3fABde
tO25hpjYPo3LJopNsNUF7GFArOlg6V4mHV37iHJSNeuf9IpsRZ1kyJ4RQljqZKwi28B9VVSXowtK
16SltsAu6T8V/kKJ/WWG0kascZ1+jVnDvuyIYreKAU56j1R22GTBJKOzZszEMMG1PuBy1cnyfFcM
B7g7LoDrVe7JkY4/hcAunEa/ZKTqzEfR5PG1HzLflglJr263S9sy62+xRS/tIYLjmdgYKUrGS7My
M+9jcRM2UqMm57sgGG9GvYC+E/RRrktYQPKRjRfdSGReYYLFHDf67PC3mxgckFZx/beGzMIDJmSm
e+sJ8q2B1hrTWI9ayS+segNkTMRE2H3BtOg4LUXnZrT6Yc2j2ZK5kmWeKvLj1U+O7KVDGA8v+Wl0
0Jynq8s9lMCF2XUAeFuYpKOd83juPXUUuEaoYIVIVVZJl9UcEDyLcpoBmW21uNhKKBQzZfL+TNf2
R96g4ek0Yq+uOal4fC60tlRjftV1ZVWn3tuwLaEIvBZD+O+s8+Cmu/Mz4c37g0eWqUvWRQu4smEX
3FLtbrPYxebgty1JTAXO7yQhvSVXVLN4J+yxU2/A/KN653nOvUcLjLHXNQYd7/v9nR1ytwxpWeR1
zmOcqPorDTaFoyPKwytmPnFFkOa93jd889JZPCwfciwue7Rio4coVuaIgCQnmJyaobrmfbDiMTZ1
GYjHPo2lnmjjdw/ad5dQXUCwsklveGrTxCeJCbk1tXsgpVWueddCp1J0XHUdZ9/mI2YK9Jr9/cPP
Bned3S7mlkx+LKUV/erVCvcgwDGm0QE9UuPncdkWV6eu8rwT6eJcHVQHEsCRHt2C0UWjF337v0CX
7oPcW1lXhEH76+vsPPEpT/VaU7zxiz8ZCB3/QY2wkICNnmCIseIMGmkaS0H4NUv7WbRdBJza6Iks
QgqjR9WjtgimR6zf2LggS9JBWCfuFiEDoWZKMmHRi5PgyZB+TDw3ywxy5u0XPnFfqOCOqEB1Mzpd
a45m8r/F5/h248J95ubqoEgEZ9RXwDcdPW7s/8lCAX8JIvH/KmT5cGX1ABN1yffaaA5yFWmeOvfp
8TCQuH2ZhibkqHey4BRcMQONpR79/QzkhSHoj5hRpa5khf+lGqZwA1C0FWer/5dCUk/LVQn/kl2+
i4JQBVEnvwXIUSiAnyqv52udEMsbqhPM0AnRTpi/zC1iDMaOHdSg4563zkxakJjCBs2KbnuGfiKQ
xiBwptJexU90NouX0KDLz+5/qmQp4b7D0zqh2QqoxqDgMxj3lMC2x5DQ2L8Xsd4pcagdPsiwk/v1
hZcasty6MLO7eX1ehP6YWVLm1q9gnO5OZK+JsZkwtXhML6OHoa66p8LKJNXLlf5DBoVQEa3cfKe0
jC1s1+MkJm1QtTQawGymO2SAip/VdGa7niS2qjECzxQnBlnN8WXF8/wtyyjWJp2wwuaaseaL3fPp
4QWhKA06IhGMpj5DVQRjitV3MhX31XApxM2QV6Yd7/m8Z1DfANv39NPwKVIPlGgZ1zEfBiHIwvwA
UjWfG6muine+PtBpWxIyOXoyZXjiAykTmvsYZ6CqkKc+4RWnHbuMouW2AphFp0urtan8G8InXX3O
Qr0WBi8wxUS2eprMQj2mZnFeieh1AmKBOhSIsVQtK3nBm2KM/fIc0Cytg6jpBIMYjjuzcKE+yt/y
VzIghnrW5ufFeDKVR29wBUquVf1hQ9soYy9XiLz4tA03zwkXW+x/H58kb3FcGU9aYicjSFMhtPHe
cZI4xUbNnZLuXKP6dCtZjOO6ebL/tiR8U1NyfzMbZuGxTnJsKJ+gsPj1os3OoED/3nRV0wsL0Xhf
FA6dh7cGGl1oC0uD22yitx/g/ymz8ifHR7ktIPmJTuuD5+RBqWiy6Op4bgaIOXDPAAp5rNIhCE2G
xbnI6fw3J9goRNeIMufD4i9goo8uLQ5APifTti/hp5OAx0b/aZJHhkhrq4WNMsE5uPeTw2wST+YL
jY4SokZhTfWg0h1rdnvGExiytZgy6BGGPT37nsxFLcbLWdT6Rh5Msqd5SG1vJGueEFLNzo3HkZIF
ImiQ2LhYhZ7HuwIdDjSmaF29zjFCCu8sFCmMHraQ4cVDRx6yMgRULMcaYgIiE9NFAuE3Zpxw9fAG
Rqem+UPvzzHhSHjY/MupuY3BquoAaTLoJE8sYmnL/1Me6YWmP6MaxeBTaYWd2hd0RlhSM8X3bEIj
l28QYYGTlPafKhConcKvLKLqNhGeC9oZSDGRq3FpwToa6Jb41J3beTk0K8ubg3D3tj/vjwcQ/pkR
R3HpXlXReyL79Mrkym1RRSMantn2KQQI695FuCFGrXV+MHX0JVwcfqAi9mS6MnNiXWhKZhnps2Qx
I37Q2bxw7iyViz+mDfYV/Unv3qqIhaVuKH6RuuNW19tWJd2hkYnfvm+rgj34mHqy8gE6Hp3FpyBw
xDvsxQaoffMACG36+2Uw9vZ29yYls+uEySsxJTWO4Tp1U/CVPG2Q/beAg2p6lQwMB3wKryaPDe8h
v2z4kVEJ9Cya6NivKJleMiHIMfJvu6q5xL4zOKjFhLmE34oinUDAanubc0DrzH766wwzsqKnuZTO
z49/qt2rv+PUofnOVtQOeFvJ2fCpSbl6o+NaCzl/9j2cD90UHKW8KcwNTGk7Qv9A2ZCZmixjnCgZ
zvBhO0XUkobtObWiwLybITYvOgh6pxfRzi+4mL1BNck1PKl3s4R5STmIHgLww9R6Hd3txogGZqW8
aTx6egyNfrRg0TO0hep2DxrvDZC+AKidOJAxPDR3hX3804F4+ysHwftftMBmcbLRkuM3dZFtCPwH
Hqq6gF3LftUnZu/ekL2xA11pcRs5peJdRTNMowQrKgKOPEY8dX8foXE8Lu9ProA1g0osAG/7qrWg
S8YkN8LEIbt5LIBP10dfnzjI7TTyxmnAnuAqsSwy4x+plqkXAJf8fFcx1u4wZvU/UHx6s9ptZ32Y
8rscICOdvYULGZOya8DLsTDsJ3e5WDd/5uaKhKCxKd1eGghm5v36CtQNMv0uDH9mv4iXYs0UN/K8
adEruT6z9aNVs9Ei+721FexenuIyAifn0+mP76eRJ0xRYq2ulB/BmQoQHqWUVwZxg/scGR1HJZXQ
xiYnTP8U9PQ6M0U6uY8p5cj5ot/YaLl/lOJFdn7nzpDHpnLe1GFERFiIYodgdjFZD9FCj+H/ZBPN
S5dQ9XP7uJ7iaT7+bANsZmv5KNKpk5e/JamiYM6SfZ9+5hmyDh20IVwbrQHsrglvu8uwroz+sbqI
cou6IpLihnN+kEFjRRyVL7oxS5le04f7Lx5lq+smhv4praj2ZWN71EnDX2RdebcpV/vS20VoHM/w
6K1q1cLBGSlXEfpCERTktIXcEE0k4F1e+G4UMCG9QyPNiSFlF58+F5oxnoL/XtVKWoX+i3XS9nih
2HIshEeslZeJID0TusdpmdnGx76Wsst19TV7I0WZMC7kD1Bfdckas6aFpVqboYSMkloWEWDABQ+F
GLjJaXZ1d4uIadmVPqv/NTZht8gYNSBlSSbVuX0RG3URzp7vkgMGkEgctpWAlYZZaDnNCUyTZzZf
IDP8FCZIQdvN5el8tvhgv9GhskCA+c6I8znIKH9tBYYCtkWQHBSbKyoNsnRSo3eGbahWB15rUARG
7qx14DN1ZbaCwnHuRY57wK+nKU4o5YeLG8WPXWtfZ+6B56xpNDKaY1X+qedpMS415WBCoVzY7lZ0
sTpmZo4hmNbBHQ+gu/BuHh3XBkZ/StOl2WzPR1WoVhWPdkpZob0yUqSExcRz8T2cRpVLoTwIeHh7
FDrYcGX1pgtgVJIstHbwMPjFZBzqKvkPoTjBxOanmVHDz9IIUgh9UiM2Gz1qu8Os4777r8U2FCLR
AuDGqiI1wbMwxAieDrNV0Z5qYgrdLEhFi2rZcjHeOCFCKGHMMZzs0+7T/0nX6gAK0OkeYfkqwe4H
msY9qnYS2AK4//MyzuHJno70WhVhvrZmiAcE8gRVGpjh6Mb/yrXIKnRb9RpdprKPGiA9+I+ZQ1XG
9OqqFc7bN+s0OVBVh6pEb28bHtLjvvBDPegUM8e5TnW4nowpPASuGhVzcnmspa31f36TguLrELdq
7Ks/bIsdwnL9AjY23EJZ14tIsnUuZx56+B6RWHR5BFLEcsu2Fkwv0KdKScc9YjaluD8SWRSdRrxJ
S/AuPnbIvcuCTk+7v2jdgFYihyRnC2T9umMAWOkuIZhv0uvcPydqZBkMNVCqkLpfNiCiR2GxwdiD
Tgy4lTEfMr1MCRX8TbbgSSRumIHujcWALIbOthgAOoUqi+WfpxvBa7bM5EYCLZGxfoQuC5V99PMt
lg8SCOf0wlJ2WJ+zgrKZoCgCjyEpEHESRkhPGfKnj6OCLdLmsU9OFncptMnluumwXY/zHKM+SZNi
YTsFxJSfuvC8VbC7QmI5AFoEIEFObBsanDk8EVQCoZNBW9N7w5ZOHLm5wPp5TZbqDts29ru78yON
AH82YdzKaykCg+bVehVSoq3XgEG6CzwtdreIBpUa8iTxpa4YHtGwTpq9VRv3hDWp7o4AIIL3qM4m
OSTgepjt0Uvuusm9zp96LcBvMX5fzA69YKwBRB4wL1Ceh03qggUA67LLTIu9Zr3MLYe2XtIwuV1l
yFOnCTOtAEqH6DbADGOdJdCxN59csm7hLlpaA2l80O8maT9FD6d1Jx4FczelEUjOQloFSHzhaknu
JVGpnqI/UqtFx4KzABOLIRmkqVAoCRqaQPbr5duLiAx+jphTdOHYA/7edJlIxwzACoouUPJWUyXm
NXaE6jGTK+okLB6McT8/nPWxOhoxd0vykNURDWVPy71hMQ9deMLx2HVdJtOD2gpIQ1zPUccfDkEw
ti7UuWXJdEgOucWEna4vhTvMi0OtoEy6ZE9f94Xal8j+H8rwmMP2lssM9/JkRBRc/XLz3zke9c2C
0M5ybmSqboES/eHsdbJPSZEtW3ejhtEyYwJoJeMdYBTDQgMhuaKovOgBNbbp+bMHvrFtu7G8mOxm
Fkd8/Q0z2PSyqgjSyzGRBjtsTwfwZxk8X53jcu8dovgIhhYZc3ajyM1rhVaas4D5RpdM2HTFywMw
wZG8d8h9q9vK+MHpLmN74+QPYIsX+dqqcWKGHExd/dYlAO6CU4CvWFIquEMYcr0bsDwnJwSH7NwC
mhnC24TOZwNnf0QYs3y0QezKqlEHiBgi0WzopGr5ymEmX6oqdBB3z1pZM8wJ1htOYPmSJSJ6Agpq
7uI8NXxSF2RtpTixMYaSeQaHDQeR1gY43SBSMEIbR8OiKn3pMY0G+ueysI9WpbdXho3J+3K458y3
bgyiCSrtxyL0aPOeyHq+bvHhlWDEsNDPKKO7NOfNt0I82sKZjvkm0xBGIjHmci8bCUVGMweNbhEG
pPGIjbSgGICXuw9tMFfl/qhIOAh65P/cmjsbVS0qhrWkEyZ3ErASiihZAu3Hj/3Ryb6VE6knBk7e
c9C38rnGm0PRndi2IKIEU3PoQ9nO6J3pRyjGlaPWmURSAUZdDgHPTkQ6fnPBulm8KGga7Fm4hXIM
KE35AWOr2aVNj8rViXsgw31G9omi7DrKcEJMeXiAf8AUKx+nv3+1fVJCtIQlb6peyD0k8VEdLeID
O38EIxm8JsaiDLEzPEyXy++gymTkSOp8aXSvaR4GeseyAqSQcVebMEkkIWjBE4I3cehnKWUnhLcp
fx+YrrAu+NirTdd0EPpNNV7WbcViLPNJFkfZvIevon4dQddYmtxsTyJSMHcpOpURx/Z5FuTRE6nT
r4dUyKMjlp4h79scfq8XCBrOACBDJDWQ3WfPTV5hAtu6ZUArRfA6V1KBqtwT53KDLBFiw+PqqMAW
b6wCeJIrfuGGwul+TEqVQwXw7W9VZv/dNT1vsOu9+DIVYBh+5/3vXXSr91JTHyvW7zVALEd0zx+j
ZBjxbjs4SLisnZYqrT7SS3PiBVAK+5Zwe9fOiAL55eeDDrDMA7459ylKsQmwRLEMXQ8bstOIvtqm
gtHQfSp/Itjf8By8Sxl+BYBePH697pImiYCC0KDCKfRZKHe93tEDNza/yjWG/B58Vt6TdONbvn8T
B+PCb6iivV6RHjA2IXpHlbRSNTr0CB8GBoH9KQU1nCU7YCL/2HW27BpeL/DaQCGCScbZIlIBPQuq
JSOh4pW7db9jsUXqswyldNWCV/VT2mRtsRDNHJ9XicsiEd24TepABjMlo+MYhktFjNFjr7f6GY1/
VC8tPSRMcfRCEDMmsCyhmq+gUyP5o2aK+leE8X+PQzbvxqXogYfmwc1hmEKl7MOIWxcofZ6hgvik
LN5OM5ekbivTuwgXFmLHZWl/I+0hb8xzl6DgiJ44JfwzU/d0AMh+6AjIH1lkL/qq1gQGE1j6Mehx
t4g/Wj1O2LOOPr8fGlvzprAwyrZGoB5eW8VsZG4wcV995IFQh3bwN4QgqllTzuptAjl0RRQ7ghZm
Cs/BkHvAS4vgFWo3kkirnoA60FyZfzWBzzD6EY0bvFNQa+dUdBBLSSDaSBFQq+9mX+/vwdTdZe1h
NZ12XIwfr8mwUEnSBdJ7uHC9Ry5YRUGeNS3dkMmvgdxpAxTvtmCKS9DZxfIVfKi8c3W2j0iF5MMh
j3Uyp8pojDOZam5aFP/Fp3Awa5yIj+H54foliT/aoNqPbf1sa8k2YSFMfbo14ZmYkZ0iH3K7tBvR
LqZQ6DdLZwIpGLNczwqLkinVDMm8+8m6HWaevSizxZFSpYW3ZHZM9LYCTyrHyoQAmcenQuDdUpLW
LH1SLFaze4pWFFfk32Iu1nIE9+CAeAWPCX9vXyHZkTrNgbtuNMRnrulMpnL3/b+R+8MJ0VghP59Q
EDqgonAIurxrBqDsf5aN88ePKiR1xcakX1tgWM3LuGeATYPLZEDBd3NyyNwqOQNpThU0sGCc0Nko
P6hi5+WAptJCUqCzK/ep7QGgX4I9MSh8mKmnw3deHqYqD9h8udNtco+7hHiWJgogREW+7dHgKyzr
eBbGrOVwyHw9wJOZC46B/14O9dv8yqvhPCrdKcy6nW//jFSk35Cef9GmJExMJa0XlXJAzxjaOhG+
Xd0JQCtMgC4IzQXWey6qtpt8Y6PHKHhW0EEG072w3CYgbx3FKI9GxH9cdnxw0CYvS3mei9vV/sfo
iP3wFPcEDwEkyHzYJPlTYMQTWCBdbpgVGw6lbFhF6Gwc1x2L5NfXvzFZsdvcuCn3Z3lP1zjWs6hM
UTSjRqiMs0/qPw0AA8StIbmDop5DjiWCvsF/2PIjRBEBXBRA7+Z8ENzrXVnEBbkU5dQuRfRJvxWO
5i3FbYSL7c5GLuc60n8v6Cfm3IArdUZcKneMCZNJEW6Tt1/66zzb8FM/UA4lBCQiPWslLCPlntSj
QpA3UAzZPA8Bi69orDtbc4CZOQxruAYpWFCljQ8ESMKakA/JHqeoGfoj/Y+W4A41B5dy+xORIbHE
hQgkhj8z5GcztHMUIvN50peBtlWQJ+Kxf7OPWGbyYrE3MYeCfStdGKP0x3fMtB52oX7aTIWS0kme
3Fqii67wCiXAAWzq1Pt9SgYxpTW8reQqbSlPxvSoy6B/xzUY6/WjfxCkcXeTJHeQQxyaKWvuXrFj
24QW+uuJ1bOYPk4isiHx+6WVAOKIpwbeQzi7Mypg5BH7DE6ErqGQ5aVc9uWzqYvC33HcTTqifUU9
x9kxqa2tVmLgDLxcWQsDuAG7gmuTzLWzA8dT0YVf6meZ+WAmYuokWQhrRqXEkSgJdWVpJ1k8TKco
8XiIvrewNfJGsNVlWfbAgxPHUoDfQEoLuITrJ5QtxR+sSEdQoPuxeVlQ0HIIqozngaRcl6BEBeDM
UbwAF0D54p0HW2xu4F3BxOzvqzJ7ZmfdlQzNAPLSu1kDf0jR9ovB30WmYoIKSJ5KCV5Vu0lKpnHP
6s4TVNG+bYBdayvrG26EM0dVX/tNLIVGq6c+qFLlT3DJjVT1dwhCle1Mel/hgBRmiaSlfUghwM5r
e56SCQmbKaHoNJCefgtCr4ynhYsV7yHED/JhjBoBq2RTwuP3urvWAy0KMb5245COkldt/q0aSVpK
LZYJdTTQ0bPCxz0tPPTuGJGKpgFjYV+kSydMU+Uwq9+uytehZR9wtHn+X+tgysMyoJdWPyy86WXz
oPyy9xyZFgcaPw9eAuSYKnHZJVLbVfeW+bBMJH3JfQ5e+uxRxtATlbg6M8wzQR5atU2+I4b+h/7o
latPr7YUKJ3UV6FkOe1IEKkQGX159jTwpniyxdIB4UZZwDUxQVa6RVcpoGNXGzBXDsoyBIgIdYt4
fsET46Ce1SpMwxC1K32HSvqo/vttzAOEmzyVvfop4oYxbwu56vvErEpOsTYwZDSTyoftBMpBSgUN
iQJOT67Vc5pNMxBALDgnqO0UDNSRr+7KpaA6DgALcR64GaZzXPXGopOESNK+fYDyI9tpEuzrK3kZ
1IIDn0PAO8vFbQTzk91YOtftqfiHpSo84E0r6FkL4oxMDwoOhK1cyK9jiViE1jVxJqbcRVxbeqSs
NqSn7/ItvjS7AJZ2AhbYQ2HsyIceY8YA909Q4lladuMP2IdvB+9gkYx2KjOjwz2KS+BesSZTW9iX
4Qbnwnav9bEttFJlK20RLgtrVRGaiuMmDqTOwg94Zde3xPcnjpyk0nXYsabyQ44bv3f2edLl9Z3/
VKfsWDHUYaxfQVaUuOmxAP3yKbUJkZ8AUWZTW4UE6sDfM89LPBIk2KFKAIpY1OFmH3TXfzJSlA8D
tvIcdbaK0lg2HR1oyqVJcyuAhmka27gzUH0rp8a5AG4ZR2p0NShJBdbs1HY8Z5jx0TURwtGqOLRf
g/JbpRnOMhBntevKxk2hpVc4zgMqOrEjlg91d3RVVXX0/TLOPCMqoyxUJFn6/Zoc0jshHw0BJJwD
wn80qlmqdJsUZByLBfZG7Nxaw+i+olI2ZhMptIU7mcE5T4YzHEHrug8D+t3Vfd03/teYq61vmPlG
eQPLD4/86CNqJ4JAlNHyP2DIM4Nxn/alaqgylvHFSSjMb0IH078CgRVmoUEC3dc+aBY3pG5A0j5d
VCFEbiMVT3SmgpZpiTOhNZ0jENZIxUog72RD9Om9y7JS4WM1dj9pUS5MNIET9fN4pZq0EeaZOVe9
0yNKlbviyp8aWHjqxay4F9xOb8A3XYy1AKDtMLkiySQ+ki927I126Q8rf5ZmCMQdF9CB7VyasSNi
UPzzT53KHhklOpacT/V6Ws+GRjcMoGXs1r2aLRU0Wh01XwDIN/kh2uwm0YsVjf03d72K3rFngeNI
JV9t2gDOv1DPKDN88woBH3k+lQ0ms/5ep3CIjrbmbvb3V9jr6rzP6tXqCdemUggNp43D5XR5/aLK
C72sy9+zoh5WHY5B7/jxx90+kDfOHstljNlGmic4CavS4jcXtzG86VlLD4Zb+bdEmKeNQNwx+S0e
Y9DcrajEGHUMhtE8iI9Mf3yaUDOocmSlBlU7RV00peIv+ksiBaCSi5z3euPW9KWfId8AB96LCpta
4f3WgkCQBCZsICykBMx5DoA1s6oChDCpceEZ5WBfDA8g1wDrq9Io08Z9Mjwd20KD9Nr/L+kjT9uX
JOf/KSMY5AAZwXOmOMkvm7PAJdh+FFQ4slpwNS/sgd4YYMi5iVV2d52VuHUNCdAY4fUadzk7HEOd
NecX3Dp6QDTRX6tKkS6hz3pgNzx+RaDq1b68Tlv5DMkxJ778ER/4+GiDnJnz5QksOM+FY0wJ8XUl
YRmqtCMX+rGEAaOLStuqAi+LagcLZT0L4Rpcp847UW5upW4GuyjefxJ9atiCwjR19wKjoqLWVl+k
0XiO3wnqzO9WHwTqOhEuOWKZF355nQ/F6nAdMAP32WzN2m1Ic79glC2n5ZULXfrsWfJ+TVP6zntQ
VgFkucF+Ckyo1C4Cwj3yh/9GbgkdubAf+w1Q1Lz14kdEd7pPaGNr4uILEM8+36pRZWaD3wseS7ug
VqvG3uLIjvg06c8EM1FsOiFIpkeaC9yi/PuuOjmzcmi8DejS5iHa/UC9if+VFx/ZwmaVCusnHQD+
SUvKg2EnsRhPIB+DA5DpVWfojcui6ufkNLnQWm0/Q7pkbDKFOyYARGk0xv4N9TEnBcEFmKK7/nGj
6fHHkhxaYJaocTJoQvJYmBJGn3lyWGf7kzfNOnyowaa2sObZlOzDno/jB6+B5w5+rAT9yxDRJ6oo
fxEKuupz/yYEBZJhikVCNUTL3BEb+csoQKBVAFCGu4tR02OcTvrLEQnVANLn7rYhi84yVBzAJUTM
znKxz5bcy5c7DCHNMM1cQ5kyGHx064aBYtyjFucjpkyxtBU0MOwXP+Q5oPPRBRlbOfRX3ubyjpbZ
OeT0wUXdvRXTOEnzDjARXJHkM7ImMJHXzKCdILCV1MMjld2SbJ+VtMYRWWDzeg932J3RPNCdiTyc
eX8UH64P7N/rRlLSmIYQuk96XxgIsNw8ro3U9StxBpsBjE/A9xC16wLbuPmvUL8TH8TXLrXdeNMM
J/uaMjZMd+jK53jzOELeGS7O/dbg9ULIGC9Zzm1CANp+LVKv/lpje/EB0No8LoL01T7bcHJJTfpb
UT1WYGLPG9HsIyd/9Xb9EKI8abXIqsf/XCoEZDSXT/3D53z/COEV0C3H71xuzlMj7LQ/OEQ95KWP
cIKrjcn2AVMTXWzBaCCkblSvtq82k+0Zfy1kaKAsWsdBUHhqjyOAc+NxvquVceJxfbWjqeodbwMX
qDvWM/T2QmHPLFmibuxY6ypTvaIa9q/AKnvF+git3xauPckIW35Dw3N378FVHStc+P18weOWfi/q
/pz87sc3bjtKV0P0Mt4+PdjJBLLoakBhx0ld+BDkW+N8cM234nifo43jiAOGffzYe4jGjaRxJIdI
PDo2u6QnDUIKiBEoOIS3FOIBoJZMbc2qzMP3UpbIYlqm8n64caYckAWAM/lgOYq47ZIKl0UKx47k
xs29SbUJteiR4q8RUD2f4YE0tGCpAvmhuysnrEloFebnnpT21kqbaNo902cvvCVzYvvG3DiYqHlr
tiE/CrMtalA+rzlgH6JF42FicAjKSs7WbeZOHxPVtZ/ooqWJS2LS6nkGYe8Kjrl38nODqxzDdb79
/W6iijs15bs0Z7uXjiVR946CtD0ZFsMmmRzWik3KGXBrtdi97e7qdwKvTtRdXgKYNqglM7cGU78s
FuYxr5yELL3ZUfyHyT2/YTa4CAmFaQ5kShlqQ+H+JycaKLsdrKuL1M4T/FWnZNKT+3hXs43vFUn/
uphlw3FxmXrVY5pYp/EbJI0EiVfbr6hOPgsp1qGXuIBm7lskx3lLS2oeHoB+wGXOiwhVqUD4fLg/
FkOvHhMhJjzmfM5TieuWUWfuuym5iI+VmHCs2N4cOm/uiDCdBL/RwNu5chfhx+JvFEtROkgLPaqu
kbZglqleAcNABTKYbJNi2OBNDShnCRXMojSBblZi3T5ABUe407G92j5Y66RPb3UtV8Vj2tJf8D35
JbIMqDZoTPUmVlX7yeCpz5LK/E274XrOD1sUHXo5M4B795YHttn1RdG90hYXnic64BbVMMM5iR2j
xQv7MBK/A7OmqoeAjPwgEvNfc1kY0Y7r/DGKAbgXPGwKcoJ336spf/1dvgKQIE9feaysG7L3Z7Tv
Treazm+5ZYqVEZewsYI7IKOTNmbuEY5D7WEgpLThCIsYbw0t17tw+3oSCJPv4nA50mGI0wMov6wD
nEx/WZ/L9LTuk8Q7m3x13e6gnf9CtMq1AEjYstryWrSsDrbqC+W1VzuIZwZFclGmSwmryS1qYyPr
/ibqxFJbRgGJWoQ57bEEHd10lC14ehEdhWhg8k6CZIp8QEeujX99yHLB8HszyaOSfUS6T+XYfa5y
0hLIS5fZtXmozK8HkRxvmY7hMF1E/1Lh/T4IWmz5395s1jBQIWVjT1zBfVX+QuknWWxmza7bLtXw
wkGcaFww1MxLnchzvVPNdV32F1VQLpH9sPkATVO2JfpaptL7QdWzgUtDJLjfQjpO4JS0SyjrFjRt
UT1PuDF7rXZS/tbnQCX9FZInETHBCf8Po2I1tSiFceQf4ndkM68cXPfp7qUOF4irWLI+Q+dQyXZ3
S3SSqwSmqAk/hcnoFkSur/0JDg8cQR5QWjaiW088qERiwTmSnBD+6bPfWqH52Yf1K31IqNJ22BTx
Myc7zm7QsYDf/2QdNzjNQf0Dp+pv33tjuV6r4d9y0DX+/rOBnWFrRUY7vXNWl08EnRvnCUjSqsON
OIfnHm4m9IVCna3f9YiXkNejT1gkyxpyHu+wLOP+8d5mLQDdiJIyrz2eswRfUkl6dinX703o89y2
LDPa/xUOA8kwizxoOKeOYSzl7nUiP9YN2Na9pRd+Ohv551uHq4SQqsVYTkkHTkZZPhXkmL4f3ziy
cPpJTCKKKmrZl2CX9SLHV2EEZzMqfx6bKpHJa647ekBVwjak6wAMA6NueONmVrH+9BWN+xbG9SbX
KwhWeI8DNmieQMJgrddZbbSHX8Y+aDzRXtQL1hndkOgZxVKWbiWrDEmlqmUY2s59p/obP/M6sYU1
BbDDK4LA59iJAlSlGrlZhR3UxpQvQqo1cNiLXzl5i+RwkIHQ6d3NWSglNfJccBiIrsB1ZqCXsV/f
3pXkDluUQg4Xmk+746Krvj9IGAh+qkM6TLx+O5xpQYkuCviEPWJ2Ss9JZwpgGZqQPWxT5V/kiGAz
LI3mhP22+DHp/qYkzn2bOANTdShiyMQD2I4RkJGaxdztCeldeTHjwxblQTvg7rphdlnmYx19+bhc
1sPbgOykJScAT3+Z3//htAF2Vgrp/C+ZLWPAfxMCEuzBVfFbzSnnkXVuSjK/yZ+l+8UpLGnE3Dgg
//Q5cSYuQO3C/xjlEMVn4DbFCmcORYPq0SJwAecG3QEPW8RN8MhsmFaWSTquQzZYsEWKxacl6aLP
HneWq1SJLLYAckzgXmFbmlbtDYOOdlTfpceq0UwbLiHPk+rDA3+2oCXXsQ+Kgm4zRDzE8kfbRgCQ
osF5bCCn8e26NDxkL3z5hDqUKBTo51m1RO8StxX39v0k/N94e2Nm2K8kD/s3/w30p03ubQoOgi9f
6AqFScBbimh9eCFSLqBbl5BuyLhhRthWii/5GYmb0ZTx06MZbJ1cmtkSMy5L1UGqOKyxjdz2uyXu
ycs37oDwwKJ/d+S4gNmoP+V50HKs+dnM56yTmbgWt/WigO9zEvkVemcQe9LgQIubl3B8jnQMk98i
iw3DcAfynuTs9sfNmp4XElNjnF4t6vJqUmoiqUhLc73j8SEoUcRYEK4ySQvUh0zsY1chEHKX8wKN
J6ZbHxP8IIAekYTvRy8PkhKVUjxpsLV417FUN2Ogcwbdx54XTPo5u8k1UVgWH3YxRHsAAUxulony
ZqY59hLejmNd0QGVfIqpf0B2j9ArGQ72eD9lvbm8ERvKe0ceGAXENTSYZdRc5RLzC7tSmZBciD1j
mBvipXi4oip/J9C460Xqvfvt4p2rGVbR/aMkzUhu4gPETCPYlGswTd+f22S//AWnQPBPvEs8CbX6
tzYTyC2/Zbo0uASwMF7UIYR7g0u0j7hlLVUA/tF+RqDOf9naun3LhNQwLcI7xBEoyEW5oKWDVbH4
tFJWjgsaZoyEEiShYy36dOoUE/AbPoCz+hZKqSKdy+DPJm6dsr9U55gDtAVv5eJpOqLCqnhBEJiw
dLuELvPwaJLqBW0btT3xqOTeeDw34MXq7JN8EWFlfI6SFqb9qH7/qAR6um81gEacXYmnmm7075gT
UwGdc0tq+37CUkXMAkF7J2mrTyj+7u2skVeR9Pxtqa5gL9IQ1zPzmgOpRgtpqG8+rhHlCKT5a4NQ
PKJKY/ESmaklpt7+eAiGb0AyzYIkoLZhElRr4/CdYA+CgbAEIbCo5OX2HpJKjxeypcpSkDbTrG/P
syRbxIHueqm+IFyBhKrkxwrT8Abnh9FZL1mqDDZvSo9RXxVQuLz+naqKWhAR9EOpgZWyCMnt3Nag
R7hod2Er8lWGztx4Iejx5vlXUKz/1dGN14HJ8mgHaUJmps3P6C6RbIBuh2pTUIRTD/bhBbEKzh8X
IgidZRhrl/T9BTV6b8WklMDdiB7qsKfGSPiQ7eg7i4tq5J2ymNb0yZ8yUyyQbGI9MS+fbjVJOw4l
KOAGdRUOR3JwAThEnQBgJHE/Gb0gbcM6aJdDxF1gDOWZ3jngpzGkzUUcMg7JFzFlHpjoC21DPioG
CrX1bkV6wdicLu4wz9bWeY5U468BntYGnnNpLd8taxOHjZ2jaGivMUEfYhoVlk2xNnhsp16+P0f7
fUjvlAGAmPA0oOqw6zM19CskIdYw/dQ8STVBEg18R3jaZeafMVAyqu8I0TGY54GMiVtGUOBTPBf/
i84GZqhQHILpjq29OaCH5ZyioznoiaU1le1bo8R/U15ZVLW4yjyNc+LtuC+K3pBPqOeaZk53tWM9
NJxjaQ4AtPV8DdDqt4AWrWJ96dAxs71sLVSgvvqgeY0/5qKMgm5JuaQgeNGn1QzAXxtQXeZgzsUH
Hytx12XA7+dJw2PqZo8CC4WmIXiGQo6Wq7qTmVJJhw8F3ATNcYxOwlrWXyjMCzZnnWOwpdcowVjo
zH8ZLse9B/L8yoU/MFwtSEqiuAz6b0m6XFZJ+EV6A8T3rWuvK9T6NmHSVkLUeAuhC9BSN1lu01bE
kC9Q3rECNKV4kDGvM4A5OfbhAhhrIV6BoLddfQq/6jmDh4DmXxLfvZ6AwzhjY3v+yncMGagzYD/u
OKATqVVPJFQk6nlLqbvp6OeQ2TH1A6bd7SPsyL0Yu3zwRpWbeQYhZQY3y/w+PhMAHjYzQI+9gEvg
lTyoBlpYLj7WXu4v0kYMIMPeYAV7jlJ+Amvc697JKNEy5LymkI0U3mmvF0oD0LC9GRnVHDNtoYzK
tEUA+z4kgMrD8QBF6r1MU4m8+efUE7mYmwRDZrrOsPyHKQILxfFeXnupT25SJ9oreJjGD/apG1YV
pDyuQ46mRBqAFVfX8lWtdxDj7FqA6tPiWN2NirggKh+PMmHkNMe6MBX+VoCkMto8kwg6hbn2iUbl
7YOyl9jHh1bDEWrNnt79jJd1UjUhowGPyoLnJkFo/LhI8lIiOy6JtMJgf5ZFaZY53m9hwchbWmFN
Z1LqB7HZHuUXnU3MnoAvn9GIF/QOzUsovbPjyC8w7/78gZx5u+cuU3zgn7LJ1HfSRilbutXCbt4S
J/VPOfoEo1RTqT3garvCRY6IA+ZcddQaaZpcw/u8rFaQ3PlQr7kvyVMelG0eHe9YorIKAc9pgdKa
+sqrHWRuj9eBgLy8w90/plJd8VW0WSom/EJekNFUsX3T1pXWLndyY2EfNRMlQK6sQuGIDotKatDE
fHlVrn7w3cn6jZVXl5VZaHFHWOScinX3NeNTE7mMo0XRLGfaqJAvDMW15qWPUgZSONbCAAPY1HQn
FF/qcg+Fwx8Fk4ssHOTqqnnuQWdsIAd3GsZGucDpexZpHtn/c3O/4cfp8R+rUFv7oEJn9DsrznYc
HJffLtLEHxnGbaZBf6eAw+0lIljkJDFs+ZliKHQymwtUZiNOIE0BToINbu7ck+BbUBj0hN+STdRY
aQwZm83TNoOWH1HkHBgu59WjFaAlt5vFun0TEAp1pY6zRRgeWk95jOVcgWn8r2b72x0qLFfXgLsl
eFfTd3Wt8KnKFjHoIAgIjxq73lMJqPLHtYmEXAQULu5i4xcKoTpdqIrAxjbzjiEo7WTEr4ja07Xq
CGLhc0lQ7xDObZsWMp/k2neFr9UTdpBDaxDpPt8afTSivOVpFVTZzd+BbEKq0PtUEzq9SSrnIdU9
7/e2H+c0lmeXoovqKiJIaALNLyb5beEgKJzfBRSZc+jLhq2vZ0XT+6acYElMeutI5/90+ZPkF6S5
pOpq8O46T/nnIkf/xBxsMgldx9RWKn6Z84FcIY2gViaaRa8kH3SKwpLSWY5KyVvcjhQ8eQCc2jxz
grBYzJrrYYCOfHajdhP9JvnmveA3oW1iWG+Cf/8GrDRcVhjOs/V/xqWHCxqSspnqGY+w9TMSz8JV
m/x3HPy3IrU9RdDyTYyWgGE0rTELmNLg/GSjLAJLTJrfd9u17csDkqjlnJfD/jOT69OAAzY34FGr
XVHyPfCsGCD342xqPZkCe/LSJzcWiy20avrUO/ZKrWsDvE9jDRNpTdiDxdVAzUQgVOH/e7Q6+Gn6
OC2vlqHLZpjJyk0jCg4sRGZzj+IMbghkldL+dhZbJMTzE+N8lr72ByHKLUeWhba4sliiE8YVpOnd
6+RY4GOq+H/KVXBhhJu3xZcTsCgro99QvavdSEPDni3FIRtWwtoR9utGA9e/IQ2LUTx75xBSa9mk
pvY92mQZzUbmFi43G6USCoY3d9DvC2biMGx7OiZTKq/EH0VdkQqBQAGFmGl3CQzTh6wjXisjuz1M
wse8lRBSchUoRcvgH4iSk+a4GB5AFlyTwU5lCP9jNdPHg2f/E1yA8ws1JO+eBE6Y6pifiLVQ+FV1
36/r+6aUeN0qvo+2kt35FwNzc0yRstNk0elcdF3dYCt3CznvyP+Rz2xjg4L5QW134aM7i9NmK3UU
wgtO+edD+3ipl3RY0sZUe5MZYiUYkJiMHI5ilBpAxzbFJy8EAUw/zd1AYk/WcfiJJalx6J02m+Hr
T28HROYXFr2zjj/CluAklfGMlOD4GAUybWoS0x+D/XP0bOIcH2Ol33EpsCBhDjvO868rfIkKAUJM
pQevS8HnMVHa+1uo/pDtceBGS3X4YXvH45a9Axm4VOv4VDYmxj+nnPtp618v/6b11gNDD0KuxN5W
0kBtmmNpEwEnR1GTksFyRbW5UeID83Bk26g76CZKIJueI1zjqgwd8AtJg9/e/B8LetZCxt5pEASV
jCHF4UCZpzaClpuv+Vp70TjdYy6Ole1V5Hf4KvG5XnmjM8YgwXB3Jv5Vn3Kt9aj/W534SPCOR3fl
FqEz15NaZQmT1AUgQi0Repc3XonYJi+8cUxnKrHJ8dBc8O/w9u3+gh4gJYhAzBDr/lr8bqpY4Do9
OmpejtsfVltvF/7mE/JXm0YocGtrEgwAQXvX0rqp76Ml7w6gytBkBF04vDQggH2MrQyd1IsFvR9+
G3Dkq/T2eMxp6gbe5Nng5Gc/M++5Q6WRoGI0SiuYuMcNpQouxoHSihvqzcCr+mxwiwsWzABcwOk4
fmOUGN2kDyEBmdm8YdM+8XoLgsT19gj98w6EBp/roXa/WY4W7+EJQEA+AQiHGCQMLXMRHSyLpVuk
yhGsrpFR70bGgF4MmdsLWKiq5TAc5VlCIQ5OPqX/myHe+MibejW5I3uh7R0p1258l6ewbfi5oJwM
urLwR2/AKfRgziIT39Ub1JS5eKZ79Ff4jbQ3w5T6idu3WELAUCd5aKQ7Q4wdzXZqrsGxww/S2qVU
xHf1xmEw+eCnq4GvFqo6Zt0DNrms5QVPd1MyGokMEaMZzF0sURZ6Unhq5ZdiVh7JlFYek+YwJp00
+2EjCyfOTJWauaL1oAOXpqEuU4CUdfKFOggMhMCxRFwYWrl0PZJECjW7iuIjQcpywh60yTtHe9xp
7qE9SbLMVyiethirjCA2XQqzvqll50BMVdOcIlST3hqJMqaG8jBS8lGreIjH9TmLPldLznUEvYvA
t6KXVqiUkATdZRtuhXD3sIGSMYOmIn1BnWrPEGsJf/g224uQy54VKpfP9Jao9eet5G0syXUXZ4p7
y+6iwA1qhjY7HK+LHWytqOwvoYW+pditYOdP+q3GVh3wuRELZnmRMPS0p8iyfKGxsyglrx3Q0ij/
lh4zE5OZcjMgBkmpo/oj1Vqofwo8iSpCd3arJYoqqSJwDJO1jSVFwo6O/UUlogHWEBUJoakRj/SH
cOJcaEUDpNB72a7iivW1S4wkaRS48Oxr+BiVjIAuukvA2Y2iYs+HIrAD2D32V0lea8tqi9mzFU/F
AVUZShfJkRkXI7FS1gbx1eM09ts55q/MjoO/0GclLlSAEPtUv0SV+C/aNxND7Pc3k0yyWysJRmit
PyyNMtemFTJYGb2GVe1WIlokbWffZWGTyo2dQTLXkZixJultm+xn7USrO74URcZI43kuBmH0gOJ1
vQU4SiQDS/5ty6N/kW6K2nK9564tOcVFo7LMl1cJNH7U+xMwCewJ4XnIkUt9kZ9Xvx7vJE8f3HWD
7EahdhRGBGHkXmgEl/6QF1a926nOmLlKVDD9xAk9VzSpzjl06Fa1Ttg3Q63KJhOeYABI2UDj3+8T
sin4wL5gFW37NN2HyaaECoLszrWX9BsTjtQLfs/iJQ3naxapmTflOXgaCxtYpOomjzfc2jcT65CW
dVao6vAwH0F4Qr3kO64FxayyaBDBP5kohE+NheNwo324yXO/h+PM0rPZRFqkwir9mvkbXnchEiSs
dQ9q5o05DBfAsXpTy/XUoDQ2eeOOSA2ZXQtkTZlWzYrSsIbxNeElrJM3UqBILkdLYOuuDg1J/mDb
U0S3KVBEZghPgKLsEhQhVbx7H4wlPt/Sa34D47PM//lB47aqrPgx2Hy/jvGJs/C9M5uy7IpK/izS
ecbDcUtRTL0KoCnBX1CZRKzhI/s5oFrxQTuR9Nv4vTlvvleknfdfwpNvlgJAwcpQITvrhBRKvMJm
mYLOCCDDvjmMsKLqGHg+N8QCQS+TBR0e0tlTv14PAz4nFZQljs0/+dNWSeNvgZJDFV/lM7pFze9F
VsExu/cGU1jgi/+DuU2Jip5sH0/Fuoq2HR9K3EjDHCJ3iTp8Uh2+DsO5nBOncgrpA42IXHkcegoG
PSS0Zxtu6p0D/a3Na5uANptAftpUXq5d0sekTb/ZCoE0+VxrPEU1R75jG9opu+JamLxb8qH0jVD6
yPOkm1Q7256WNbHJynAZo+/84b7jFnvs6o5CZkRtPuZSFRKqyXdR2AaUV5BuuN/KPdC5PPz1EVCW
zKvmoMtHJ2Q4+eGK9SUvA/coeD2WGM3yLbOeEhYSoT+1Y4apEVs9ePmTbm/md4yLKTiCj3jlD95I
/RBMjSFfUs8vnYneT+v6vRbTC0xMF81Ou+6azpj3z9V1d3IwoNXnJMs4IRTNbwB8huvsftvZgD4O
WEzbt4UeA1NMW7MVig7RA0PcLsuLJImlyHMF3eiMt7F21ag371Xkb4qDAci1Ggm8l0WZFemoFB0X
LwrM6n9y+6QhlOLaf5Rdl7JbJDyi7vcnJYoXOej7bFyqRuWK9+QK1cB0eihz9a1DFKiFDF7rbq1l
KyPgj6V5e1CnJg8rKKPdF9lM0P0svcmRnu/Oc+MdQ76pKc73xQQxDn7Fnw2NA/lmh2pQCToE4ZBL
AqXhAUKC1fgdBWyw8BmHAODg5X4DullIFImmkLJrm+gTdFLf+akbsATRZnRkg4Hcl/UGsC1vJ5Zm
bRLa3XMTzQTEyiSCsSdw4pYbPMl4eG+Fd+nOz9spknZUlwKZeF2UHMGS+np7dKsoabW00HU+ixVB
Ka993vUXBwqO8UHEQp4NA8GU6WHYqKxAeiQr0xHkD1xrKzSLJkiNT0+BNJdOGx24qtpkYyX/qZJK
f0GOke0dT46s03b+kFQG+UAnJ5vQ5+9dL/F40u9jyIdeju781JcwXwIjA5e5PvRQNaB3f7uY7RmB
xg1sc4VhxxWGHq+GHSBZ6qjXyizimdUoO5Xd9rekDz4ToDwd1B7xYTTxdoY90jZxp36k496OXLCt
jE+n7QNTk8VHEU+l8KqY1fGEkx5xwr3cVXcWIQHGCFgyMxMxzRk2TC/sd6mVDyJznlM/qbf8DQvc
20juuPFRrORLaLBChryhsmrc1WOWEzg2xGlOvce8C1Br1Ts70syYQHxj/Q4dhyAXie3TShTt4/Xj
abxZTwYsCynLUQqFBQQhPMbRTIGtMrpgLXw5ye0BUiGK5LGW6cZ4BVaFgdNB2ACA/Uu4SGhXKev+
dmExcqncz6FVVF8XwknbBkUbSB/GDHVQPg0Bpu2lt+xkr1eTumUbxR1rkRqczvqDMkQVyllFEaUH
P9tT7klbgMBOkS6KNKnV8S2GoFUzwPC0F+YsKZcobEukEwvxKbH3FBDpa1qEi+5dBY+loPTJSq+o
fH9w/mLvxbxAYIlCOBCTcTKPwp1dSjmYEd8pr1xtjBYsMgeg2aJwzVBoj1TrF5YMZiPLQpRpRUzP
5lzXzVOOUhQOAdU19edGMj5F5qlDGLbIQdfeKzN5O4rqXo9Db0Mn3GEnrBqo4McUShVJmaj1nf3d
qOEJjOVZ4UIGUDNkyedJdO7e2HW22Stw5bmU1rCUv7ecfg61DvKggl1zJlZsxQ9fmA5Aaw2TBvGp
cqieXVOQYbncBg0z6Gx/qSF6Q/B5WJ3crTM88E03GjHjGpxNNvZ+WpqJi9ZbjSx5rVp7h8oYuFev
vKERxCUOl1XZuHdx6v+r5Qn2/MbBXwk44vjKlw/8Pi13BiBEiGi5iPX90wt0ss9NQhsla1pL3Owv
fOP93zZGaLxx+DBwFdTXBgWQZVFJztPrJtgiNyog5GcGSORoe9wcHSZmXhr9wjWNfyoxSbraCPrU
AyDP6eXpTJ/yqIdzsHL9sq/7x/CcEOC23lg6+R+zF8BIsoTgeXcC6Pqcp7+mrA3wXzrlBctnthww
HkA/KPHlqt1s2Z/L36vw3Z5Yqr5C0gFETnIrtEdh3Ee1he7UO3cfopLUFeM77MPk+DCX0yKdwjO5
Dr+GH1E8ZbnX8tqvfZpGFXKsTO+QVEDc8LcNH5N3Hzgd+IJ7Ejv86B7FmO3YHpHGv5h2FMpZBAOi
BA40njCygHPsBA52t8IUKEZB81oRjV3tuUheaMOOwUwChd3DGq33F52BxmFiQG91OHYEDr4YCCV0
FtxnUVNnjn/uaxprmtbG6z2amCYDnCvFEuxH9BhMGSnOUzrTuM/zhnFFHDloxjaH4nuydgaJc9Fh
YiyZ+lsPYCZxdIvIE3x7vAlsNFu3XCwZ2jzwF/l14BEdaDXPoEvMue00jyKhIaNzNiLRFNICy+Wv
MgGDelTOmV+7ordPdddtLphT7ocV+5jB8lIViBqE4kJibP8k/f3xJGvMWysdwvSemDMRrStkm5MD
yb1bGrujJHxXtwqDjquEgioRPeYMbQEY5P6j04z9k4H3F38fqCrBCNKhOH2lSeMNbIMSImzPgvj7
aFKlWPfZhKYca4vUcs3+oXVx7jHnSTbEsJjQB5s83y7qIfLB5+VOsdXtuEpVXdsh5lssLVKJ0K1S
gqahb7o1eiFGJPXyooEQLHTYKtOz+s3xo33Sff0Zf89ujGWCqhTwaZ1I3ah8VzzYZZCxXEfDQ5d+
rx8A6nVTyOPlmnowpraiF5qQ4aqkfFwmilzrEepx4TtnSlkCrQksfRucPOyzKExquzAXSRjUnMnK
FGadxbM3e66yY5ZZycdrEtq5UTYtgzfU++zyY7zIfHeHQ+BeNXWW3lfzXQjynsr6fJEFpHz9PEbJ
n3Fu/QE8cYvDcu+cGLVbJYTa20u4y/t6JaKO4q2oacYhXGJnOSwe+EDwo47LNSYk4cQOFS+l45DL
z53YJPyuUMMf0599kIH7dhGSQOBDOEIDItPFkl4SyQ/qo857fcWpyipvYDzedDUsjpEoEoOjEkKB
9YEpYaRYQnFYP7PdUt9BLbYBSoZHOXwMY11RY5egU8xoCz2Rg0vbr5fuC8aff81HYL9XyAC6SaQD
B+hne8KQ+PmkLCXwycXIBXNoauJ55cFJyTcKUC1HwygQtis7iIT+YIV+57AkPAjJW+Vno/gCgWeL
SlT38L4+QQPcjfpUbfYciLHQva0UYk1MZ8lJeOffa7pSET0nAjgAsMq4cVmOBqz3gciXYTSXwKu0
fOzEpUxZdFHEQ2dm+l1hg0btvGZVBFOairjHau2a1LKnTCmOCpe84KAUfqec8SV72CPo5AQKPwB4
hh1fATGCb4vVAoArnuIoAALM+yKkUuo9caDca/HsUdqbp0I3mMMIY1qMmOJHCt93DWQIbFpw9+Pv
eo6hEUGKzJ9/MQpJtPkHiki3QxzLcBzvCsUhzS2XOEZn7dMVQS3GPlkrj94grgzXDTI7obIK33Vu
eB7I8dV7K+qhy2/E2KylnK8dl4czu+s3E1AlM3muF25kO4Ljc/wl8wOM4vwFFW0Z/OFh16UGytEo
9Qa3aJ6YuKOZbDAbWjt1uOJ4nMGPJzjEH+HJ7Pb1/wpWszAYVnWmDWWkgyOcL99iIrFB2JNlvNcD
NCJG8zDjsFA5Yc83cYDICCdQPjDg4eUjAmqk8LlmE3QOL2EhK83pumDJDQRkDpCFx8UKTw3n1efS
/4X+oJ3oyKqmZ41sydQHSMc3UifsCadJEyI2IIPilp/felMDyxYtNzSAdWXD03E/XefCaVyMbgpE
86ehzbYlpvOuu3I3uOTRmESjSAwTEeE/mAZ9ah0PlrMK+TZz3Ch5M5TwRt3NbZltCvvwobOxD3sW
FxkxGppJt0rQAEl4fp4YzEVP2CVRJWe71XuXwQSXgFHifcIxXGGV0J6+tR5xMiar9oTFGnCt8kWj
gWo4ipsf32qN5W/0Ot5g6YoYHjiCatcAOphtFAbGrjp2c8N+fDYrnhV08mdb1Akar5LeBIdtKf14
iNTVUwlZXIBpxa/0CCUSgwKYvLwy4IfeWVGTBLZM/zHPLmtHulHx6iTI0eg+JlsyaLLxpmpvk75w
K3Nwz3JoG5KmafUGYYS5o8mPeW6uzhoQ4exlAZRhiEiNI/sx34l7oWznASRimirnai40aicSG/gN
zKNiKPv3wp7cov30kHoNQOlxeYrZ6thAb90rz0+8tHuWd3be1UrNMs1RbFHT5yjkOaN5zvbkTzPz
BZtpkTJRiUIrmX7iSxY64crDwxw1y5WKz9dhCo+ZHGpS09ywAfEPBQMmuORbvA+OqVgfwIi8/iDN
PMeZR+vI3nMyekWNjxZlpjp8sjKCuy7qrOyAz3LiSwr5n2TvAmBlNOQVgijI6fVfYpR4w0cTARRY
YP5leT/KXCx/FPG4KPd7YglF03WBC4uERGWiHqbonTmc2LCrDEuBFde612+ZCbu/o9kWBy7AZgdX
kyRZmD7x6eqj/qJgqlYBZ9ZHc+absDNZFL+eNYVz6ggNHQGaKx6lMY35iaapKIYgtroLQWPCsqEl
rbSXrCYYqmGf0xBFFliInjWD7QbLacY/2UoOQmPc2CMyQAzqIuDGIj38maqG2OKRKxZMtb16iFJ9
Q1aasF35YXETQnVn6PEpgxhksekf8GWUwGBLepLlidL1WZMIcx2uvbMWCA315p+QxtWA0gjOArmu
RASWRU44kA7Rv3/BjvycJ7PQBYVYGPyHUwGubTLuFaCV6ZHskEoTTIGkGJJQAOzqfWjRiIec6+3u
WuqfqT1U4L0yGOmKm4XXas+fSeHiQ+DjMcQUjQnuhKffm8BSYrico3/bhEmhc/Pxh8FlqbaAPWvI
IbV5limvbxUTBiO77unbfsZ5ue8G6OX/MKARDkVpN9JrZxuK7jXtzj/uG9O3On0VYRhTFsLIOs9Q
CLymj97/aNOWYFgHip7xtLASLquvbJG54br+zfBVvxdqrJJucTjgkve49ozjystn/oR/ZPyWDxgq
2pNAntmRsKJZrBMk05eaWCIed0U+z1xrmxsQyfq5MFggABzSMqvrwcFG54Z5gnOA99lgaPUxh77X
Um4jJAAG83spV5MlliXN7q5RF08XYFyZuvLhlILZuu8qrzJ40EIZsU47tV2Gu3/0KjK3mSoN6r4/
nATCXZmOMKq5qW9BI/SN410QTK+MCo4hwNAtLYGSvW1lABqo7B4MlotByHw4dXWofBFezLPxJL4M
s6DjFVJ+e/RKEPWSWrVAcucn0SSI+69oTwFsXKEic5k0i7/uVF2N9Tvx7todYxy1QIwuzJjrzvXn
AtSjtcW8uscTaleAxC92el2XOCFPKw7BycWeB8MHbiCU4FFmSbbe3+vuQahBRWcAnUT7IKPgcN90
FyQ2cfSwLrfrjiN1DqqRPZNgr6bOuLMq1qTPzlExHcGgMpUdVczLweCWq5z+uG4EaJ6Fgi/LX0lr
g5e0Ll2xJHfgIxGhJXO4OJivfNSqiuEfsZUTbzGY3mgG+dvbc/ToEYlbVSAM897z+ALzAwnl/tD/
9EOiPqoIxLQ7dFya3W4x70jsQqcKosSd7SRrVm8PGoM7ILLwEDXie8kDqWVBry62SoxnAOgf266i
Rb7pLN9TLD+Z6igJIPUUbHGj8z/lXEvqRhe5BTZBGpR8C54Drzb9SJX6ruI04xwEDmXNoUdhhIJt
UiOeUpcFC3j16ltviMY8JXQMwkvWWHjaekiwIzFAWBznHw59/ukT1lUyUF0VRgd936I6VWegkvRJ
hVLhMdXRebfZOAK5pUY44Zdl76qzyn+oHleXjLWI5fE34LUN4UB9ehho3Z8W7N2gnHkNntl17PWj
M5FyrMzFwwLonWUyl1ihZ5pz/lO4yzI2hHpnslbMaiW1Uod6cjHS1mMgsKlTfzujqGySeWDnUjCV
8tK8UzcU/1koD+G+xvxfTXbryZncl6rG1a4pmz6CtFUxpsa7wPL/3/5MaSyMStMbXDW1Ro5/PNbc
cyJezRA7Y/k4KWRWapj9+t5FbyUhQRhrM+1MVtotr0CookNZH6mLJzpZluhReUXbTO36Bzxqo6s5
HRu6fZKa/bnvupP1DjH2rXa0Sv0OJDRWNX47AmAK8EkTLbITAHVHctfT/l268JlllwrYKThiAvRY
0uYFrbpSxlkNKQN71EMv0jMQLi9l/uZok8Q3K9qud1KGsRPZ477zmbrlARZJxzcos7p8Kc6/sJYH
LnFoj/JUMPEt+eSetjSDLUk3a7mozLK65s49izq+KeaL1cr7lg3cbfI8AuZIuTy0JCkuSnb30Y63
llqNW50id4aWjGD4r1r7ShZGbLvj5J0Y/ahJssJDR0upHh0TmLNFifMlj8ngvkulXKAvtAVuhCF/
Dmy1xJQoogxaVcxZ9qPNNcTK1a27jYmFco1qyJVu+bmDQQwK8ScfF90nf6d5GIWuhiS132RrE3el
OvRkn48dQRCzPAwWPRJQSvkhuNyPlMW+oTV/+vcuOm83QYG9LFp5g0uENQbUdsKoPwpM2FXXSvxi
YYkbqDjzRbLM2UVrDYQQGohb8WzIsv7QUmd2kOHHlFHVgZwq/Vl15wrvwJZoYwETr0kA+CPqmS7J
gX9MsVxkApRREHb6BMIz9ilmOv4nTJZMJtTkYKQQZB1eA4gPcUej8NZl94XmWWVxHDpmYmAwajL8
ec5cekQQiYZ4QpXVJor9n2/dWQOOxa1m3D3eZwGN1FiU/wmN/Zq4ixOfbegMImPCLSbWdY8pitGA
wtA8juucUQ+WSlIdKtq6XTBe8Ehro+IFV2arl324ZGewu28QxVqecKgK9rC6Qmm9OOUgqGU+iWcb
G90iLeCfCcL/StVh8IwDSpopbU56eEzDbKwF6Gc+slR6M08UnIjrxnPcUJvzJS8ppfTUGvIZ73c3
w/nz1EVWgfKB+OP1PGOYSOohkoi96+/qFsu3HHiu3MerRlG2jHuln3lBSVe/vozce9hpzHuJXBa2
AbrKOtDY/VAsexQWGdYCRBntYG8T8X+mbUolbGMNBsIg8w7WybSthbRQ4cYdMFzi59hIadEP01Ad
hiKQVdHHQp7KesFDKS5aU9CwXof/j9yCunyM4ALFj8nZAYO96vGi9T0B/4B/IqGyreiJ6/pmtQWP
r9Dn+dzIB6wnspcPzz5plFfq6nMLbWC/N4mva2QSAGoKui0kNzPKR/9IQJHGPf5XwEdELo+Jw0fr
db5fWvJnpLGIWvOyFNs2tSAYdhHtYbmy8SopubwdAq7sUCHw+qKfLfMYM/+1x7UPxrSn/u30XpIf
mTh2tlFrDleTOOuqY9d/TyfqGHnkfLYtp6HdjgZoEM/cAIBLye4yJNqWJWbZXk02fQ8ZN1KZjWM2
D1xqghvBY/78w38KfTNMdP5tauCNf+L0ahr04LAy9klHpLtETvqEWyxA6rNdIl+1Xib9AxLLjMqH
WY3xN3PEMQaKRMS/eeTlxYS1tmCqipAPnta2q/Y8xmKTzhsPL/l3bJA9FcWX4LKhIXyDOSnrdUyj
Oj0L7K25zu89w9vrbrCQQrtIyEV0iwXNtNhr4HvL5moDT+xPOIr63WhBS6WDSsWAbex1ulwhVZds
3ubCRYAR8c6fcttDdiVh/lgiLDVYj5IT763/QDUar18yv1gWBY2+WucM2ZtFRfqxeb46Ccg1TWgV
jaYjuhL61L/K+tQFRz19LT+j/tOM+Zi2MHf/9CcMdgUpZGTW4ZSht6PtvLhuYG5CKc3LuWooDUND
9vexBqr0yQcrKJqKootr4+kwyM9+xJY1A6TptoN09HrkQgDQkuZRfrIt9joFQBwSkQhgFLgVwEse
5SapceYSVi+lln/+abmyVaw+sl47iCGKNHAP4+C4AYP2x/Xi4+g0z8Hu8XxyvPsx20SAtYKvRNvU
vuioaV/M5I92LHgbYAMQEVX7BeL7+tQzDT1mo3cCvqkGJuM3glTBnDyuQxLZcSM4VGs/2vjyqnUt
65rgA/E0HXRRjFd7jSIyQcVAn2s3HlMG5UAmPh7f+D7hRIPWKET9/gVrxmzjZBI6AuD87RieDlwJ
3s3fYg2yQsUckyGaWVLTzxrjsQ2ioo5Vm8zw0dWnxU76cMTak3kQUm+Z5i/doX7XvtqQbV5AhoRK
y17eytoRmz2Pn0v0PjI+Q2YiihMvzPgaDEwXGHisTdzyGTX51y4h1wLZarQivxpghRWeRoal43uA
c17MFGSjsuGMuVT8Jte5EsXGU1aHNlGbMC6W+eTA04Tmcdc4ykyIbe3sTYo3wnnERp3yPmlghJPt
gJenHfH0wCzhpGpycNKGz5RocefrUdtd14ZXMlIIRoLx/oOl5iO/Kgr2cg1k+b+YVaI1yUiVySVl
FlfZJjdZBhyljbduupmpwZ1NCSqEMuQfH0AlKKGXnOhPLK1go5R2gNcx+1YZgEvs3sAqzWlbH3UQ
dy5gqjv/v3dEEHLiGlJ0oDXDk7CkaTsnub2PDDRGU/fuaCTiGlfNuYSLG8cVQ/37GozFbJTrKTl9
ljbPZPQIU8m8Su6zS4pqoKvZ+RFo/hrom9ipOeo2JbrvmJ/WsO66NXmZNr8E9GQ3moofDzHZjg8q
vKgDkCWl8fL6nWeTbgBMiMQr37l/V8gWee6IqVYqNIZjY/ngB9nbdKexAGTxUQlh9Zp2uJ4cB5Cy
nE19S85HSh3DEkI5JtwvgEmVasCuc4ci0ecsSEWpgwnUH7gw0z4w5c42w9C/G9+xP6WCqRRoIsTg
T074x4WkeltwO6kZKGfAK6WQt7sxsMWoJF8Xu98iBCgjDFYTkYZ7vgEZGT45VLsA/r6Lsfl0djRa
U9WYewjqHVzmWBwe+EUdc5hoq+InVnWt3FQ9VWtMi46Cb+nI6a9xl7lDzgfl3cH7SZeda6kV/qgV
75DT66v/a3mCNgmqtGbXrwqy9Q7sSSna/TQpfKtLHPbaetTY2r9AMTWsgsVcyeLpYATnSDBLadwI
KxfKBS3A8TKXzLNwah0GIvrIuvdICKr6QAMydzEo01l52MnDGJV7mHKSXhwZCtDae4nXqhg+bxvj
wVdelfvv590A+iL4OWuHgKqrDQVGPWrkoSswtlm0/nuPd3ktpLH6uTirQuMamWtCfAKbYkaADteW
wj+A0sQFO1n6e3Mu2cm3AHJMRJvfuVYypvxccD2AKaRRikb0cSmWdKTn6XSJwvvPc0UQ59l9XUpu
KT/IV9oqEVwJYNNiqrMqPfUW1YbOstUAs/pGjyqdJAMF2ufz1Vc/UwJTG/C8cdid0wfjn3RVWzro
BAcZEmBXegwYR0iwBm4LOn+mnZqR4fcoDCpgMP7YckBa8/hiOJy6Vl4zTY/lnfZ6KBU0wvfWh+XG
s0/ccR6CIqmeLctuXpwrnu3K1LqrClxelZDVKa+wslmwpoR8g6BHWTK0LaTpxTK1F6fAgwNH88NZ
bcZOWphN7hxp9+CacmIKMV38sysdZiDM/LJFI3NxugkxjfxORbU9XCYIYeDrjdhmpNuTiLZ8g7Qk
jQe2vvtYdlScg8HJBynG+qhpixGV8u0Y4xPHAq7hTCFJHofEDnf+5r5iAPe96IOBc5C+bPn4A0Fm
JShY406BypobNlBncp/kreMOL5f47R+oI5wNgirJHCCFHnF0SWgjcB9JEfD2V8vIyNY9l0qN7m3A
VfP0t+wkMSUs4JiyzGWBJ3KyZTG5Uq3sDLk4Xq+WiG5pLDY9LH/wDqvgdAiyyytMnXdBmQeGsFj9
xb75f8L9woEbFLHWXWxQykllRLmLOzHoK1J1ImZIRouP3Cwd5y2Gwq4fYIvOek7WNwVC13J8QtLI
YpIVVy4a3Se20cqDIr0uN9w0XEmop0tXeK3pgLMFD8iwA9wCAUb9hy1rlZTCf3vWE6qTbWMyMTIV
K6/PXZa/zcN+51+73kKDwUt8W21gyVphBDEEJlxlJjs8p28ySj8uv/Z8hYzkWlqYswjqyKfN+q/W
u/7fTpSE4Nk+LK25ZMrD07953fv7uzlp3o5Fo8UCdHFsioQ8KNbPhDh2PmdT0UHpzO8Urt5tjQI/
paaIjnY/0CzJNtBsdEkmQylo7EeVIGIveM12dJCehV9nPrA9BkVzZqIzdYzyKlDqKMwCzCXpWdur
Fac7s+4G7LlRS8ayQM/PWpqiscTQoEqClb4KCwnH7JovXoTfVx3LLXMuIixF9fV7puRE/Ug639dm
GxUHuXy95fx6BR+rVVoxvKmaFJl7cMGbUOtLWhaoL7owGtMcdlSLxS/nWHJ2mbfCV2dVP5BAOJXC
P3Pna1IBQXZr/RZZ6Bgoh5qCKg4aWDKa0Re9YR7SzI1bElPZWu81lWiHRIN/+a7FUM/pYcAJ67e/
Yu2KdoOzij0b3GlosOt9QHdWGdrlLq0wqMPYDyqKDv76riwcibj3pHzMnRJfuXRmOMo0ZufKTs+Y
Y8md44TsyeR9DX4zj9X8XKMidrLQInLDpnqHszDJG30sbU+pxZZZy5T0p4Iwdgc6GslfyWDYcF3Y
KJdX7g932a2ksgrNclb7415mIy+RVNCPlqrKu8i50MULuHaoXfJ+LnEqvHhvo1zkkHXCYLPVioFq
1lYFNOqBuunvzphqMKkFJPHG+Hpcmtfju/XcROUDsMALR8kEyecQYzroWWBdmzxGL5Zab8Uxy+db
4SKFc8UI007jpo+8UIBFupcJQ65D89m/D1AlfMXXFtuyN/7ZJ1LA7RtnGU5zMKbze3HpcK0Ew1QD
/lzn/14lCKH76R91dB5DEEnL6tLssp3URwBDMuC8NGNhKDQfPhRIwPNIZU3R7gtiwIMgbXXnIvqn
hA0MIxBWcoGFz9GH8RYpm65TIjKQAi9N3WMLZO86Ma0ehCPgCKpdyYZrbcHWKTMwAHW1aCB5G17c
QN/YQIp++Xors7YI3ynagG0ytQB7PafnTfHdp2wdF1z2R0Nt1CwOFVu3ZylMy/hF/r8iax5K2bKw
Dy18WzosLze4HBTk8oUpyuHCPo17R9Ebdl3uUMaDfMGC6jvcn7BKyzUWstm+UCJ5joZkULqsXe5F
0aD7CDmpJtcUu6DIhfCBQ8aMeGB0ShI4WZSbWUMkoc/b15sE/ZCRnQKiGyt6ETJKqAGLIpV7J3MI
HGkGAOMt75yZGitjjeivSUqPZLXiOvbAm6XsWraET+QNGPwnsY563u6ZM33/vZzMtfCcBN7n3ppJ
Bu+4PfKa/fv4eC+iXwc8aMxO9lFNosS84LKOvfboNRlvVEpu2OTBQt4Lc7hGyAaeAF/WwrFLItyR
joVF0+pJPuYoj1fE5DblTj+z3LnHRRtnBpgcAN19EyxcMu6UxsU2u/sW4tkloxkKvFxRCd8Z6ZaA
ncFetdUjonq/gioJp8JHYYbHJ02MGLh8iwod+XiF/ncSAS3QVBxBJmz+XcMG+IEAKaLmj5zNkM/k
re+16p6x6DkVNoyvmz8RwYigIEx8qG8mDdtykCny3DBXtg55hnHpuw2bU3V5D+p+r12SbLcfCqJl
5Owg4QAk/PVierfDuD/2UVVgqP2wdNnKuh//XsQ1uUy459Vo1H6KjCXh3G/Yci35TEan9IjCdPMF
REdu+r4alWfzEAtzhXV46L63tnUR/PevfHINZ5VZ3+9o/WHz07ct0sCKzo3yW+xqg3LGAutDws0d
cob63FLJsy5vfXPtgeA6by6aZQ4mAD6erQ/FEbVE5RZ4Api5Qjcl+d97zrJ6CCzKXF7p/luX0+LU
CuOzNPO8y+b1KL/2bCJm/XF7FAUTLs/BmbZU8srMmYwP6iXpHE7526kbyHG2NP3aAqBFwTVJBYsQ
GSYoXkpUQJVoXKU+3NdOY/NuEFYJxeDJCA7AiinJ3QBVRyqeb1hKOCtQG09vedHJfFzopbvkRv8o
iukmBVwe+C6oeZBO53uDAIUzrmLjGiOqhqWca2pPVN6l2P3qNusP9Ma/RjNzPNkl6xEfar8oVC6h
LNggj8+NmoH58JE4R9GZfPDWuNjsDUku7Z39yDZMqfOMDzrQDLbFRJkFk9Xgf1aBS3s3DQHnR/AX
+R2NMi9wLIfSYiBb1QI5jREhqiECSqKjuACli7TzRFv6QsdJIQEKjfFEG1CPyB1mQUeLvHH8+aEp
zTfN5SLh/zVNiWTlRmJc/iAOysRzYvIrM6O3ZF4ZpqajgxEiLpHp6pCW9mIFwX+HHkw/RfrU6z9e
JNBhicQtDuQc96jmk3Lxo5IRoxUBGVz+q41F8OugNep7ywfQyK4jMLnNTkdUmRu78zIGKZclrE9J
qqrQ47aGbQgk2ECmuL/O4FiRM0oeYNd21fBayDYLG982MirxYz9+FJzUD3v+0IJiriOSJ0ejPk6/
dyDCtADwfbFwChG2h2J3y1BX9BpykzxGbqF3BVyTrTRDfBaHwtsM3Z5XBBmcVnkhSjeb30jBaF03
6PrhLYGleGZlsaN7qqZf68eAot9OaI/BFeDJCIUKgKBCNPf05wlOh1U0SfIeuPLiVdgQXX/pbFHS
UtGA5fWPTMcWKCwhUgr1Hsyuqnc8pO2kbTRkTmDtcX+7IJaX4lsvkEIv+DJT6FUPs0wVgh1GkGKw
ONRuki93syS8OyzrQOB33weWUkp7RbxmxsYI65m16crhZFLmok1YPc6ppNb/sC27gAfe7J17KrYr
t2O1/D2LHUsgtB516lAU7oURzqJggchxUUgU1LQUK82Apo48+bcQwopiaODyDdgoC68u74SSqLQj
I2Awmu8A4b3q9OfaTXitlPm8haK+Y11IWiNkTz4+RZ8rKtVrf0+qx+WgVHiznBYvvzPTaiW0EXQ4
NNJyK2odF894SnKP/4ND9acKPesYSyxq1b8Sf+I/W36JgLWHMCJnObCFBH4j8xMC9Cl0sg4GAM1T
g1KA11wyQrvd58WlQ0w6XVG0QGQHLQgd4Ah3WykFGsc8c6yXrfKhs2WsyhZY8a8/yBA6FiyS+mg3
MvAxGWVkvUzQzoPAJdhvEQeySA6LVad3LxfqIPkxqukQQmri6tr6M7T4T/nRoPSGZ/B4P4dLRvdL
xB0hyzpf0eW38Q5IWHk4ymFHIYW+TLSh5D0QqpMf/b31/upE04Y0cmAb8tJBrsXVrLKqAJ92mALb
jzVAlsNi8/0py779aYKdIcz6i/Ni99b0Qt9w61uRPc8utaFMOSI9o2d8SxmqkKdUcisvMQOXlW+B
4S3Re3LhB3QGEP7RCksdSJhMS6Bn4RETbb12D0NV9c9h69d551alouti/gvRZOc24kq1mRsH1AUK
oL0duvfUZOWW6Bt5iLmwPfOXy+yLT1HlTMx3GesLMQx+o0+kppMRngIg67F8Hy6wRkw6RiMP9hzR
QJUsBUAhXh9jcrELdBJInAu9zX0tiem7hZLVn1odY8kCSCbWQ0ZQKqmQwrY1TiLPXTBT4z7xUxCC
H2cIzuz5ESHkSbZQrr5NxaZSbir6IL2xyF1H6Uwqqo7U+6ZoOjQ8RWHleI8dJnu4RlrHqOlQDNaD
Qh87UaSU52/ssnkoBRbpPBQyUYjp9CXTZR/3zBdVVp6ebUcYV4uesoFTIa2OqDO5CAYeDTYxYmaf
cc50ZVZHFNJmTnQ7lt/Uf6w2m5HeZ4/FWzmSe8IFUGYpY0psVY2SMyIXfoSNy+G46tEdeYV/jFif
dRzItdSfPfnM6joffUG1go6GsQJpMnLOSJ13QSilLasLGZFcQpwqTqOZ6gbdGQeXnep76Xscrjtg
Hr8dB1HnsMQsbOoMnPDMRdB4ayXg/5fPHzyC5EWOt9sK+fgyDnI+ugYPpU503hsFR3qqMKrtJywS
iZfYKunv2Vt7obr4Lw+4H5uxraYMCc6qaaw/YFeRlsu82hmg2RvF2cqNtQbdXcsiB0wtP69Afvec
9LFowIWU58lJ2lqHkQLBf6Bd5fVHdNzuQ/ZDK1+0AfFUJpxF93FGii5ua/fLc5s7cC5yHGmHwLCW
QDLmVlUPOEtSSOoYqfPHCz/DHzTpVV9AAtz0ACxA6tEoLgQJUhuKUvDCoEdT2XI1XvbpGpKgaFgK
FfYgW7atcNYm/dJdWTc9ZaywpgSx9sX1VE/1UmFWvU5iMEJ2cvSZ0xF9PkAs8YDV1PugBTa4iInL
GyOtUejmtwt4YwzfYIAIgF4V+kuBMgxqWMNM33gBqN2JmxzJm40duuhCN7tbdf/vGgE+HpPTznX+
6i75tF9ajdFLuN8nLgZJaiabCp+4RAH4LJmunO00V92Qa4R4LaUQ/Uw1pdEe6YdUNjKDlQoEZrVY
/wnjidFeJX6Hb5Rd7fhFRsx0l3Ga3UxoEXe8kjx4xrCYBU8c9TbgwppGYF8MspavODCWpkLz2KsF
jW+Rc5wPEs2NptH4i0AIIdBuc5c1YjMiyi39abpPT+3HzpGt3J0BnTANN5vnZ1UTTs7o2QLr3o9g
wQ0iFUWn+hd4jMQEJZDS/uZs+x1FwKRhn4wPL5rp4b3qD1wVodJGCImx1At4JYxLkYvCnXUPANSC
jXXCs19/VgIr0YLGp4PXgY76kSdTsW5TDP8eCH3y9z22690IRoU8FJAbXcrvL+8yHFJHoG9SrxQC
QDMrNHKux3Ll3boy5Dp7gm70bS7xvo4jPjk24IcWEe6pN36/zhrIhOqvM5HusT/wbbt/uFJVa/Iq
Ri/yN0JIC2QHS9UzO3qTIvFJo7NgPhOWbPdn/L3ytrhB6dNT0U/uN3dzUqL6ycCIdmWeGsxkUQLA
6T1F37/JKwh0NAokPWGN2cVsevCbLgqOQtY6mRPfJK80wEWSBhKE0GCjVqKaimXQ2X/taqwx4gk+
vuhSMIy97KxWsnVexfQ8GpwDFKUfdNPGrEE1GjbT8UtfMaG6WdlaOz6fMbLLvoyLI9FujGSlGNey
8VO7y+C0UvugciMlHBl0ORC1IX/cVD5rWx8uknUdc0y9d3vmbpz1UOcGv8Dby/i0zmFubqQAnJmO
oJMCVKpn2/qNpuxADcTdSnw3EC/dPgNX8HXeWp2dL+99QBod/ML76ImtoNkIYub1A3rlwHk7DQF0
8nFbsZ935J91l37LVryhTAI3SERrXjwnbvMi8bR2HgGl4hZWbfAHAmSyf959G3yFVMCe6nsVfcLD
LgYXvFb+TVinfUXf27MkLbojD4A3Nte5lxWYknmyy3ntO+sBrRVDTO9kx1atOQDy7PCsXxEraQ+z
DcUG3hlXaPUc0eA/gL5jGh6EZEyQWapQXCOGedm0jT8xrBrE1fv0njAeisdejAT7/kul+At3b7Rc
zMz880grC7RsM6t3aYstrsrb3buZw8GEmcO/uJmw25H2XdGuyp6Cpq82n4iXCVk1ahTxTxWnWLJM
FMwuQ04GVH5oTPDOJjA1U1V/Th3W3C3RFuYCXfT56uKKlo+HhMFHYOPa3hwTYFrRP9o9s1bXMRjG
OYLVLorHgzLuJ0vo9cTTYp94wmk2mI0HU3DW/kq9/u/xsvmea3kI3irqFcQjicanmfKbYjs7K8t/
CUsaENnfZPQ1KEkyUQax7CfWxlXCgXyrb4Oe86JDhpRRWzY+2MkWD8pfVL2bXfZe1qXTQjOi8+/c
xV7ACVajnGIVm1qh7TBU/9Kj6EXKWRYUHhLxreJJwt3pBiTCQj2fEY+pfkR+1NyB4I7sXoWDsLwx
X++jtv0vucfX6mdtW8rmfcps9qH6O86dkTxNDak61b7UMJ2TZh5rdIksohKmG+coV1khewi3MgdL
8d1NWlOqqmqBCxHwNW/d1p7KgLKPi0jBacqd6WodXy87fmuqpZ1ZUT8ai11cEXH6UQ4TiNK8u8UV
F6G4QIwLIlyC47xPBFHnhuMwLhubcAu32zpjUdR8Ljf8u1M9JulBbpnUpA1WOzbzokUg4ReabZQh
Xk7M/1RIyPDTgeHfQwjx0AB3zNpKlw7YToL0gHz3+qS96/Y2Xtzj7AkqZHVeuZQafaSEoqFxrnCv
+DpUmMGJgh2I802MYRJU/dCZNVN+Em0KSX1jTQikiOYScPiSCYQnuQCi/i8jpaDIcZr+hIlMfM98
BvOQaA9K/Th9MHHTZ8Bhp26KXSwwwRZ0B1NERoQqSHVTLOdZn9kQmizAUo4QbN2L/mrXVV36Hfj7
GOEEIYPqlD3xweairwl3LL8gWU+9NGCDKVesHzpvl4bttt0IJezrpHbk/mO6c2hxVyEYjpzDwE1A
eqwMOvbr1hepe/Ym8vX2kfnmjKXOyEChuv5cJDMufGFI3i/PwW9koTO2moiDSBeQZdsBhvoYWRNi
pfcNNDFOp40YanoJfLjWVKvF7FsjF6OThx/Ycx/em4RODPIc5c0uR8rYjaO5l/B4TfpEBoBzD4/I
Eb5nbve/jNxzunWmliUnfEYN6/b8yo8tNtv7GucQu345LsDZgiAA0IIHDFD5jWWfYUNFtsqoNi6Q
RrrQZOf1k9fCTK3SaSvqAQBHmIB7jeIJ1EnvoUNZskOJDWACSgsF09Hf37X6TUml59A3xn6jVhkY
z31hHdvGKD9B6ubdSRFwIaEOUVwEtpf1bcRMNfFNCQHzJoSnoPsDmaXCpB2oFRAfiuLIqIjZqx/+
k5LJ/WqOajwr/A2irEGh87fUBNXkGZCn9vzeWNKWWITSnemdbUD34bqltLF3WzyHNY/gIuvVpMOH
xZn1XHpzLwBeE4tlhSsDHwLZq+s78+0j8CwpPXBOynbckdFai+gFUzZk8jLpb3PVPVvd6A//su0W
nwyyYAfs0sIVl7dGLPfKj75Y5VWoKpnAmaRRY4cWVu5r1WtcLfmB4j+C1EwkoQlloenYTE+Ni2lX
z+TLeJr07h6OeALpavh42pmp1l4pwwWVGvjRfgyHE2q/2jpjzrBRonlb74IG5JK0jYvBjz8/GEs9
kfJODt1PbbqTGsZW1CappgooMOE02F9p/KP5EhB50zUimHXGlJVVjQyRRh1CWbnKMso+9EOcskRw
IudVSWaDv7FLjCyC77+S87jfVuB7+Ayy9vRYrz9dxxLHsk1fKlvi3/pYJWRUj4FXXHKKC5y83XxE
tM8hpFsfNmYt8tjDUploRHncOgeTb7FFYzmssS2wH/+s73TBnZv0D2yG1y/Kn1BMRbhOjQw+HHR7
Xpzgsm5HyGf+SWyLPySEjxsU158MwPlVg1T4PBRAq265rinrUGiV4kCPU6un+lxG1p7tVlaykufB
2NACBKMLr/tefTW2IC6Xl3WcaNHeAe/db//oUm7UKtxRHhiQYDtO6tfU5ZKlFJUAZG6esMmjuJem
zcx+OhcIvmyT2ogqF1zcnGBNJEkjlS9UwRvH/yjOzrLfgZRYej9IkwJv0MSQKp5qBdLMF+b8DA4p
oqtXPoFmN/PHtvANYv6Am4luaTyIwIMSUnouvjAiWjfo6R/KHbQHWsjXUM7xghmdh3o1FndOkKej
oQqsmgbRf1qFSuxG6TBqnQPl0gDr0oUC76Loxyph5FHhVoQaDo5giLIJLRMyZVYZPCLlU/VF8Sfw
f/MR048PRUn0p2TG697VNtiFGGXX1xRkMyD1+BSC7qrXl+FgWYDmUfB71ywYGqrfk1bNendBDGVS
Ohnb6mZijW4nFvzfTaj36NtR8eKIw3ZMjGBrUKMTxkiJOzFZC4cdkfXzGAFJC/mzXxXlYYFS4/3h
sq6G5/GmGmZXsghVzav3uKkNvUKHoFVBal3QXaHMWqIN9ur8UxtyHAbduuUGMVUcC2Dv50MyGhf1
Tt8NTkl6ib9yJD/Njo82BZtTtGhYKdOsuDSrBgQ5+qdLAyh/S7CNbX04oYyaKLfgIEbN64famn2A
OtRiffzCDdZDa/mE9lZbu+tWrYYyUDTBUZC5/Cu7hy8equcs7nN+ZYSnU40PAOnlmb0BX2JM1aK6
tDN7ans7CuM8sWWiE/IvO0t1byaN2ZXv+l+dkSCtg5JsV6ZQAgS15kvCcB3UcBLIfHsJbINtvlXD
lTexKt2yTx6U4qzLN0SKKDeIWnkBfkt9wAQhlWqU2kau+zApNVYcxEEGT464G+DxwJpBNd5JJ2iV
bYe0BYdEbdUBAC54jJh0Sd3I5IqKuOLL0IJDgHrJLRrYqRwzJgUlsKhIOSDxAwRcrKGa0/5gB0Ar
7N27dGJFIERbFoTS4nwNj3aWttk7c2bV7iYEkCygfuWkr14O0qbx1g1D7/4c005pxLlwmWh+oKri
Au5q3TZrQdxrOVhfeRu6QT1lti/A9TVMbib5umtQgdYvYm9LfuimSNtUcxvzWWDuG1WY9VglEt/a
8Qb+gApYgDkx89OCKGySRrOOyHu+sObUkZVgnCYhJRy3gExJJ3ugoEbUWp0ohhVhBTmvAkeCShtP
I60tdZ3PrEoXB062nEgfXpDCVdUVJi1Nvtb48gu6Fa5bHsbkfNFcoXIJmF3xDCkfuMVIjUW9pdD4
2EPliJIl5YZyvRHLrEZqpsb1TgeDmQSKA9QQOEW4+XdtsLjXo6ESJI3Qc2svVUbw1T1sjDTiVHWk
QPBfW7fN3goAUGfEjZ1F/hIDCjcYUsY1ojKHPHhKSzPqmQUH5f1pZQ8zJeiygngfmX5U/Qjhrujc
hKwzSSA2DbcljNWfesXJM1FPMenAPIVlik3GW8NzomGZz7xqJK5UJ7OCWLmrRtlRnP6/vzEVBgpe
nyBt3ihMC8krELXi4FNp6UYOWvSoSAtDsZ3/tEINct13XmNlvjdruyP95IqSJBLSAkiMOwnpww+z
EN7uPruXxp2Az8VaRLP4VTitk1Kv7ZOAAyTVupDWQsDL70mLYtfp8FZFpgVRN0/ga7gfUfqMWUoa
o8n6U682KXTskPT5ZO6do+XY8z3bMnXuSl7NdtckArNzLABT4RcrIObYGBIScGkGZY3N+06wqsmA
VYY7YljQ+09M50iOrcsHd4qOyyKlDvBIP8xCaZssZZPXFt3f/oZi6mdBzqq1hePYEdQlER5ThtaA
zOQYZOzf1Vkf/KiyX2bmcC4WILT+7RLfQuyiokXXLh+p/WLa1KhcEETUCYPdcwaLYSwrAbTgYO4X
71Xg8qzD+EK3DlRG5//pnoKTPAiOsN1eUKM5JHLqFwpf+DTB2Fk3+jV6kzIYmmdIKC3IeMi1g8jg
YV3IhwKgxwRsdS8X7VbmXmFzffrW8z7VCRcSBdP9s3FZUFvqjCNvuQQ3PRqk9HG7CB4nf9tCpWF6
3GnqIhblrdcc0sXmOch2pXM3yOwKOVx9Kcvpo8eN30W7zExfDJD3lSlvGY1BFQeZ2HdBKzpcTsmq
43GUDxbo4HXHzv/LQaIG8h22w4MpNSfnF8NuTMhxPivwI5VK7xgmx7mHAIV6gKoexB4Wn6KHcK5E
mVze0z5VNymhxuG4peY7N+ZpYBApfQspF87DOnRL6ZWakXD/CxWPnciZVjKG3Gi2+Muspe3ZhKT0
mVl97W/6h+EjMcxcarCmyqkEYoe3L6IBX8mpJIEczQZwG9cdXXJbrtuAbt0KPnizGIFBPHQ5jCup
KKZVJyx0RovT0vJLFvo1fZ+2Qx67K+3YD3HKeknnrKz0yEA4mtAFDYJxm4Dea15g6QFqXuXDz3tY
ezcBvqAzfOGiky0yE65yNoW8zojoup9FnCQ1u7Vmni8bLZ3LdeNJR8PimmSVywCv1TQ55rp6smHL
208XbgKYLqQXuXpY+EjugLNeh2OnFUoVamUrUQukNXL46nsfcKdA7NIXEbQRj1k1Q97mlO5hRS/h
8KKSz/0QuMA0HBIdx2zD+n7QYRfHJeL9DTQR0zYaj7h5tUxTZBmEx3v8rAZFoQnMStgcoxsVZIkr
ZUbZlC3z6Gla2fMyy3achWorz7fmX2YqXvgBeatespBw5yxU11hkQshRfKbXWvpXdSps2Z+8y7MC
P5eS4JkXdM6LXBmwcw4o65Pcbar/waJxt0zSJlouEEGHvBRRav/ZtR3Tk29bHKJPJQm7pdSMr0Y3
d/ToNyMHdWgXFIRZO+mr3B9UZYGvSpLC75p+n2dCHzKFD8PlQv0kfp60LWWGxfgUbW/yqCUubv1Y
LzTNlZTnG8q4RhKZZLMIAg5IG4yUPLC4mLO10v5p9zr3+99ygF5NEIqI0fnPjI0vBEhEthGZ4iu4
ljvAOXT3baWAzGhmSqUAyUKaj7nBDJXpI++15tSG3V+Zt48/+HOi24W9zf4gp3lJqzcwesqFqjzK
o6+SgezbqNHG7ltZrcghD/S4UNyM4UX1C1x0QosV7pBlT4B6glI1Ujc551shPg65mhZNowOLIQqM
uG0QSP/M2FA4hTia9yYmRtEgUKskmcsbEvZOzQ0m/+vEExT6y7jgkK/6QR1uAGrVsSaqPU25VyFW
lwM6vkdnUaK7PKBAwo/exFjEc/H3wYACNt6ahh/tV4Mi4eEybq7HijLiQXG8ws6NhbawlqtEEbGv
UW8uJjSfmCfHhR3A4HS4y+iTyEb/YpPWCa6hTBsTTmWyveeEV18YW2CusbE3lKfgeoLMoT4mscah
zMAXgb8v+msXie9YNwDxxv0jgLQnwW7A60/Awo7xWCF/HqtiiJQ/cZogHJ2LKP4oF5N3nFGLZebJ
lM3QRukql6PQlgC++/6Stf+Ye6j/JmGEB1JPrnxt4gUAl63BhfUisYZbxKYkSTql4o+/JmTAFcPS
9UWEVtlWdS8JlyAfrXYZrIrz22a4gyFDd1xRxZt3M94J917GnW1tita2WLwkeFQhFvczw2Oq7WXG
zz5xvxEBI9b8pfEEbM9isUfkX53P0t5JdtGzUpJ6ix7rMfatiAqNQLyOSuL/S1M34t7W+RqH318p
nwaaoAN6GYRIB+Ks5daiDbGXLrYXabWiAEfsZxVMJ2Z8bndi4elr8ecydQGtriXp6kf9FVOuXQe9
aV2a2k2Mk70utR47iZyFMzYVTUi2md2EPH1lxyzqs0yYTH5KdcUjXIIPQOk8JHRIIHHPnYIwSxTF
LeBRS3g8i2Y+wDU2iyoJswXid5z30y5qYWA0ezfMG/qgvVTRZjoZNM0QutFfbUk3gcXfk+esitqE
9tErbtkGfNbULnn+wGm3w7f6rbbaVbukEZXzkw3a6TVBj/Mz9JO1xowqpOiJQhJUvwd3ZqQYqhVN
rEw1GGoZQC0Bs3tpKC3yriCbah54UeM62vDVsAkWKh2/Dw/txH58nqPpbL7vOsPGRjaaPcx8uHnA
ZBTDA5+sH7bRw9hvq5ivE+DkZx9mac4pwIX5jTItdPRE/U58Cmdywi+bSt9hPRaSOvzoBoHrNXQs
cFj4UlkKXOZMpWKqiWr7TC1ThrbBVv7EetlvQZ0KfIlFuSuhw7OdCM1KJ+N9sZFyzIG8/ZlqtBiK
deEP3DQ1gg/0NP//0ka0MDVQCTa8Ae0g5LCApy7kGF5UFenZkWmnRiayLo7xEyouXL30sCsnzYAO
ggos7z2Wky6cqC/Q9dtUDhYRLx10rKzKiWDKpx2cYxZbbjKGaTw+GJmtfFrspBGOV83mTzSclGl8
EQUugl1fOhN5q1JVhop6Sao0eg4unP0xUeLPFeSKG2HO4NcEkr6QbpncFQYejY5zORc014kGWcIf
Zhvl7LH/G3ERbII9/EgCQozQwKWXf7vHslveC18JhTsr9iQ1wWEcu6Tl7+EUrTIY76SQXDR274Wt
y90roZ9eQNLAVUY7IaxdcvjRAJXIgD4AbXGGSlFSc44+wZBpPomvjjf8WEmMGlBrKoK4CtfYvNgu
ADSPDyjguzk9VZxyYtPRZLz57g5AHEfrOPewUXDxIaoNdMja7bPXUNcxf6JqWxaSLWNdXqpjM/6Q
BGS68wSzurbk4f9XV5E3IB8amBAGMD9+CeMaEguiN7YFG0Wy/yePBKDU9cgJkYL56D6qh5huM/ug
fXszw2u/21IUIJsheMPZPLPJVhAIGmyptbNLbPC0RzvSIcZ5JR5IC0Fp3tLU17HF97jb9IJEpEdP
ZY+aFw3iiLyRq9Apf6DNHPEoZTBpyuUQk9OmRjSOcw/lVj9huXCdFGNBd17dBUR1WtvfkpHYw06P
z0SnttrHtB7o2Gt/Wm/B3UDohCDwkh/LAxsK08h+FjSS4RKIJ4XIisvSPwEc8LQHJQZNuYuHay2M
xX/+aZbAI/Gp21QxAxampNyFBtuTsVv4zA7Se5dCxOew1CoGgMl61FAcjQkbMin4Nz5xfOuJKS/M
NGgQ9oTXc/9YMkWCKQqHKFUVIUUAT+pKhHgTo9t/vynpAwHTnez2kmlLWns3zyAxaUVNtTl70tuv
TA3sIsHgTdmUmNl+2fA3AOPN/9eubJTbYBOrZDrh1Jj/T7NlYjmS+mJbJ0ePtiUdGEk73Wofb2hO
pCOXGEe+oEcICu9S41pqChV3MPPT1ZE1YdgNaN85SQgcOPj3gL4n3tmbd/GoYEDbft55gsZVEzsx
jU6SC8bt9hRR8Hu+9FadCDN8wO75VR8++IMON4RseefpiI1UhmA/2W3lk8gpd6/QsAYNbxZ+Uo8H
yp8iFaImBjpF0uFSRPMP1fWuyos8/NSfBDcDDTH0F4xuz2Nsa3hYrF11rWyxdnBqN3RndE4IEQv6
NpwQ2iRK8TshHrLO5+bdlhVTj0ThRay/haC2Y6mSET+FJkxpGmNqrMbHtoci2q+ddnUNA9ApsayR
f0+LjOMrM2ManXVw/cdCXuz3FaNJ2WG3hu+MwpuNjqwNHoWnBmpGT+TUXu8bW+ALLOeSJNUR9SVs
PMUqk3iKOlcmcrVtbazQogRN8lr8S7qLWxXZ/M1WKOP1J4OKGCfM30O/yrNPJdhLneNPu4Qv4jUC
Cdh1pzyH6xalcVrOKIbHMiU0jerTdkgh6MzzKibyG2NybVEaODKnXbQyIfUA/KeVS96FK53ctyZV
mpTsBrbRPwgjd94g276BddTCxPEwKqhIKilD72LUqnNwlmAf14HQO8sknyGqSA2gVmuZFXkRmOr5
zlgMHH9K/0n1jHXPTnUtZs09dap7lu2RKOA3tcPufbO2YFtsEXd72jgWqmeHpopjbbUmuY5VEP5W
Dgz+oqZYbK38Zn2PSkOzNKzBLzUppD1DsuHLj0r4AXGKlDP9TwUby017RZlwcr864emUKtF0r8cE
7sL3wHZCrKVh95aZXHGjaelyeMM7hskTIHri995Yg3zDSI7qUgnxwbhoYdt1EqZphGhGSnaMlq3R
2TYuta6NglgOstaHwYjNngyac3b4w1wawARbQsH1XNbFBgtgz19Vb2OHEgiM3aLfUfB6dsfm6FBS
vJ449d1t6QxRhsvbxHxJB7i7Bp0p1tlhPNXjyPLqhQFzXjUHLcyN0SsXbKEE7fylzjL6vH4zmnlL
6tngHlINPvcJP1WeEJZSHw1wfVuZYxWyr+7zKTN1cX4vmKYIrslM9LkANHFod1LWUX9y5bAAPmko
PFkD8ery/6YKsV8qlwZ9A8yMqFxX0EF6yFwdc0CNCZ9mmgHgs+HNx+GmWLVUJrp207/DbDmYs4Xg
j5RSS2Us5x9Rx5aIdJz9EBVByfxLw8phHqn2E2Egq8MyaDPuTiEXTkV1kcjZ2IjobN9g/qIoJTT/
UR7IW6kiRhyLz08pOPCy2q0vvcel5fVt/wrX1BKosCrJqtfJR13iIhdP0Agnd6TmdvgsFbvEARy0
Z9Uwxee82klmxbSiResasXp3Ei+4s68qp/yGywZu0l27HTlUjt05F+H3l0B/s4EAuFx07jWgKHN3
RPRKCsHYEY1yIj0d7o2EP8OsTmnCN05+RIKhBfXP+bc6nR0ypJ3wGDUg/Uae2fXEvik1AJ+/M8Ig
CYbo/gTnNkv52miftsk74yblPmBVSpTD1pdwS7l0QywgJZ0gLMmtxo0aa0Yhfb0JLNbigphB5HxT
R2cer/rRYYeHGvWIztqx/Hv61NXWx4JuRGYh7Y8bS3xbgah4LczMyDtWVrsRKrwUNmmTvvZNAeQE
rJnPY9ONzIeHBfl8wWa12U2KZd8RCv5Jaf1ejlSHomZY4P4GipSERf2u5ukp+9wQlXQzvpemSOQD
CQYD6CwI8kzhfa+OF6ZmejXNdVSVR/NbnmY8w3+AZAZvs/1L7q9Iwy0mkR03i03/2pdjFT74BrsP
OuONEWhMWnM7+iAxc3gsQNPSCjNoEreT97l7LrrLGDBjj55RALgmp0VJjxw1W4bh6NwGXQa5S+iA
CgPYYD6Ih0Tbp1rtvDy0PqKkJCu/h1fFDNuZAV1GpjsCezJJRhQSqHD0Rwkt3Gaq1YaKU4gzvzla
xREANjhW4Sm7sSiNlHIiDwYQ0nl+/r99b7JZraFEmpNczYfOgRYDNhpTVDZ4kRmJ0dIPkiz5J8Jf
0CqQWWIpCxnC6dfsYhRIB+0XevsQEQHuLleKZ3B0S4Sx82YVanRbA7c+99Woxb6rcc5JcEFTaqSU
NYMl8ndypGcrKe/Roxsu61O9bcametUxl3Mpk9WkpoOzRA7DkyGSJcRIPdSXDGTi7YPNwuPq4v2z
ulwtBXC+cz74j4DYOE3HTArW+k/Mk8+Yepoz2FnLlfsRvIWzdtZ8b51JffRDka1sF5674UhKwfg1
5ohBp04FYJOH5AnKS3O+NINeufCMNFnm/Aqd/dCbS1Fk67gfGSkHlwe1fUhP40BfkKSO8pEkEJVN
SC2n7pNuM1a0G6/JNJo3jP9bdE/fQ6xc7ONqbsJesmHPbBZpvdCy+wL4M1D+ZTV1N9Wze4HaryxR
m3ZZB3+Zklb1nqCYlQVtlVlx2a5Q4wvHZRCQAf7TAo8av+30g1HdJ8BvnCgIBphBzePUYx0MlRxs
n731+4tncOoexAk6NuDqL6YyTXlGPV7Np7dDl9st694DVj/uh3Fkd++i0ISBTsUOe9akrtl97V88
26RD145EZVgoZN9Y6SmFtNyhJem/BJH49h2i8PSfxidl5xYV57zdH4cpUP7IGE3Qn4PrR8BtaINA
AHc9FfWjRuB0TlKGAli0ERq3QHwx7i0zOpai656kUY13xW9+4e5oX+/yCz/S0ltV0hpGodmju9J8
V2fhsDtuEUSpKBstuEdaqASg/YrmIh9t61fMiBmLWXJNYkDb0TNJZVCfcXawA9gmHDHFL6zRLLEs
lFkZJNbRmxJbm4oF/GY9MKrrbmSJ8tt3tQrsKwX3aaltNsGI6QbH86sj8Mj4Aa4wY5P4r9ke5iNH
plmSgbnBCRowTsxBpASOLrbYqTSOCeGJesikmHnEchNDRkw8jmiUIzNEw8JCmWa42o93nDS2Mk+k
XWoumxjwxRXq8w9mrujP8RdbYp5IxLyQK9W76u4qbUkjaeS2IiXvjT4vr9whcXkHqTCexMg5pVJp
BiCXR7uF0xEFlY4MW6OcRQA/7S5EZZyT7maUcnIrDbL/CfopoRsqfRq3T3m9dm0e7dCTyddaPWQj
Vu5CYLJ+fc0u3yOhttdbuJWiPFdX9xbmlk6OhuALYM6h4wrQLJasp+E7H8+u2G2N8nJCvrlBgLza
L4voLN9fiHutYaxOpioab/5ArzMpUp7QhXpoaXqstUXzo4xhpnk5n52GT8iCyjqbf0e5b8ka2C4K
yfPlmUTOWKqe8YEyep6/6Ia/7q9JIZh9fFfcgAPkMmY+a8QDEK/HD144e9pbcBu8QkOKgYUdsOJ3
SMOmt/Lv7jM9D325CBuctUJuUVyn9DR+F8YlvUXvCT4MyHiTCdUWjCAucbZg/NhHgDnlxgmyot7v
W/ay1hdxgZkV9o2FiZBGUgNTfaDPk0oPHxTJcG4j345xFrj2J4RCN/zCc1vowgDt5vB1U9vhDm8e
DFbyoufGo+mCCi209xxQ9ibe6fMHuULfUIBZ56UEHmk0qzcmQSiLafDIrPncGaKmjBxBUYOqLZ+u
7EJ6ixlvrK/u5TBJO/q7LxdmWSIMz241kv3TJDajO991ZZ1yju/GCminSWOM47DHRvXOBJTxpFEO
ekSc1+U+S6apco33DohvNca4w5KBcRNmM/gIohyD4n3u8zFZWsoc6PrGHufPpovgx6cJMRs4kjmh
2TFOtLiaI0grHIiJxj2l/kB6JH6MSHHt9PBUD+UIF5O9NJZNJP9u3/WOFFOiY332ZPfTmUQZMf/A
N8G+SInvjFdxktKBa8kM6J0ykWHLUN3F2Wz0zC5tTYt2XUhRm7K6x3dO9T4C600ldZszy1RB1fIJ
muHR7wniQFDypBNSyhNvAP73VkKHC6mMZm6xXDfxEc8S5v5kNMzI07u9ms4h+IkEyWAoCDrKZo1S
kwDS9NIzZ+pLFpQm4I0CZl71/8GOY1LshidKC3t34uZr3cL813Wvm0eL9yg9Js/XvNsCpL0RVip0
gH2wOJ4wtypMk4z2eTNGK4knuz1XV3n4vnXKS5lOSb6R8kGYE8192AasJMzS3godxmkB1cd0NKUX
jkCoi+5LfpPNgsU1HSl/yWOPFs0sUR7sm1TlgMEUGlsLKbiVOV1s0UAa/F2bjiDPcz9D6mnnkIkq
rlkxQXhdsxnPM+2OLX1FIvIsq4P7qcXZNqeFM3TASWEuJu1pAQad0MXJXuYxKMGQtZbZHVLxBpLo
bpdWk4xW+CjgZMl7FuupgTMjHAAsKsb2DpmFJukNvOYo6qWexSP5pMaN8RCx3fdqI9kNV98TKYjA
X2oydqVydbGtqz6OHfa9++tqgss8Uj2KB4jndR6d9H74kC0b52sWfCzJa7yb3l7D73KZJMDicvmH
AiGC27jtEKwyAZHh+5s+sOeNME3LCzbOgZ42DYmSDXPhKLVm1ztJNzk6CE6VAf/9Zj/FDM/rZohW
tlEkjStbyV3xfhvmORigTELlTixDDAs7yLHMyPdKqfzIKtW/HX5mxhBTm413t64iMMpqEcfkDae3
81MkI0Sp9oSDa8MfVBbr8Tf4WAF709+iNyD8mZsWB7F/icfdE/CD0pzP5EUhB02B1AnCzKy3ITPp
sDZ12L54jNy44MOqzcXG9XRnS6XiOnxszXhrA8jnl2iwcM6Fuk3l4btJRH0fFgwIyvkukidvVZLd
/AUF1EOfiwiTPtHP1S9NnwjTclYubMBc+0nDpMEg2uHNpKKtSEHWrK5ohVBQlzbTGfmNAMSGVw9m
6gat+EfdKjnhuRx8MRO/1bH2y55tNlCOtYrXQIZ6Jev3p2W8s4Yc3m7ATBnQJUilGzWp+XZhqLQs
mBoXjJ9WoNoOTqj4v68B/BZ7Ja9Me+WBQunJWR5nn1nZ6anguRqfBIfmGrkKLQsCBLBCHHLSzSo3
B6Cr/o+8H0aqAXEAF2VvBGvlWjrVbZVfaHnAGFw2TeuFPDa273fps7xKFNdIht3/fa7HvWq6z1ce
0dYKeodSV/85k0CqQ56JKnrk2kCAjLaCldzcf1RYp4HHJ105GUZ15DeZ4qEevQ1m5xnu9nLFHQWV
LY6Pjt+Ng/lMl1UaNvO5thUgR2TKhSQ/981Uk7ZEuqZeC2z+wFAXTXi/Zw7IBfu5D0uixpdcFY7d
P9Q5GAIyTe1qWhLJnlu8rU3yxdJ7WqTQ6pLfHaF5eajGa3dzvl6KCiiQsE+2RBtHuMNoyamxIhyL
O5ErMlRaTLsiCDtTgEA7VshO2v5vC9GIyNFFeg8tqbnQVw3uEAG+dV/aD5fkvKz3tfuScu2onl4S
Y1MvHXHbH2syR7JOYuT26ap4lPz9J3hDk7dlfshJu0nh+PLJVm8rMcu/pRuSKpE1sePijOEBaB8u
yHNQj2j6RNf4JDvOQ9lW8utVEHN6ttK8bdwAbOy696317rLJYM+SM3G1OdUykvQ5iyQ0/LqkzQJc
ibSVPZsWGYtH4yk0SqtbtZbVVsvI3FcX7KfarkIl03jROV2+8/4oo7WjE65G4vgsJ7sYnJ1Iw+xS
YWAOELS/mZFo/9l0RyM9imfST8Poj3YaeWuaD+5tEmhQet8wTpRFJtvyRS/Ys+TH/aKp/WZysmp9
2TyFSjW9nv1UJ9nL/E4+wkN7DYFhETlX7Oondvv/4XSYQAR1chuDDo99lA4ydhTgp5/hgnrLM2UP
KwDCVSO1zqmELhHOcsVah4YxFZs5SLcZ+e78aHRy4PAWQzQjTRr/A/yaY/dYacWkNbsI9ru/x2bF
VczQu3+vxPfesL2zdQ3JqAX4xxEHcydZj9sQIRkcvdw6wk4SwsoHxY0RfrKrOwZFutUS+p3MZIjM
AkoYigJcbLAFAm9KYy4wNU9Qi5S/z9xgi7rLxPtcP82i3HH/cf0A+87PIj8OcZV06aO87BM2+4bd
wciiyQCp35SZeM2U/FnrWiEd/b9PIN8FYLOt5dM+rWLA1TGYLcgTu6URN1Bz5BHH7lF7bUAtwKTY
Ot3AcPmoafwuFfeQn90RTWQ5MSrRgWyVGwBxFnhnB6s7+ubn3GeW4SrfJnO2ZOT12dGxZbhmWdgr
5dKCoeyTWxq5ACvW0fHYrUbGX/x73rw/iI0SntnqQwOpNPxyuPKl31S4ZndYY/V52IbRxmBImzwq
BeRT8fUtq7QBKp0BeGFc73DjJ2tMMeJySNwo9T+RuMKjizUK0bmwxUacrEYbCLFFOC4MNj+RrChQ
AdgnilWS2HJWWmHSGU+xRSy6aUC00Eaf+ag/etOmFKD18Z47xOB3chriQdpP86mRJdXhdnuQRUCL
Me/5DcjGqLyz5I6cMNl4Q5D02SZtPAUdj0K82ySnh1U/uObs3USoHIm5HZDgHIk/1LMYap/ektv0
obs0RybH/PiOJbWW3IBbPdtvgJfuyZKt2gm6AIywSijROHhqMigYFji9Ol3nk0FjYNYYllF2iXiT
1+Gs2XE/5rISm+Axfp7cRv4gHBR/pAa7d8aZtLRqzCXXpLGul8ym4UtspwH5w2091jAR3/IVJO0g
kQ30RUuHvXVX6X8AJhSBksTQc6hqsEJy+dXtheZfvn0EKfQriWfin7roISiymKiao+wCAGCNdmW3
Xv0oFWjIpKnWapH+s/L7nQg82C9/bxyat1rtgvLuRiJINV2DnxJCeYlXrvVJV3082JfOjpTkAVaU
So3b+npsrPvA3XQzIqBdCVg/BqzVRIq1vT0lwsLB2EvUG9rNegOSHiQ/xItcpBIcJLE+0R0xekdV
UTbpHVBuzDSiB3vtg7VmaqhWmSriLyQnZUG0dmhNGLAgND0+tzB8mjCNVXCs9v84pR84TsXVnxkl
S5sSb0eo0rkpesZvnVP1PmN69CMmWbEqN2f6M8vtILbAmUslSfRkj7VVa6njupYwgPC5SnrNanVP
Jr1FFLK8Ckcc2B5BCwEOzbSj/t6znuBXdm1CT9+AxfKECfsG7fcyryOZLRtl6ShCN1dGelTEiSI9
QLfUeuY3WgYkXElTzEsdoMRyGbtG2I4FpcKte7nBZGd8garyNOprRJ/OSebuI+eIM5p+YHbWVK2T
YtcdYc1XDtpfs+X4X6NfLQKeyIrO0Lrd26Doj+vUkxadpgxT7QU/reTi4/sNc9i4iuIroeYgt0QN
m6OS0SghfsUTshekA/pmVUqEqHs3RZpA9+NNpbOYVznHPJR4pyb0JGj6jQ8Fsnj55sGWgTIu1voM
O/vJWu9NlWRBmBYlts74yX31HlBtELog4Ju2JrDv5V2LNTva6BKRkGuY9GXsO/nzrdiHzgA+xlMn
30rFxybFJZc7dqJrLEBrm69lKuncxmM9wTHfHIPd6bnVWf0YOLw0/+/8S5SZJoamiMuNwIhuwCka
Uh2peh6HnEO4cXJu+GsdKigJrkXG+6jwgK4TmmNr5i9GQPkrbz4+nCxH4jFqrxTMi5+D+Ny8H+Qh
Z3az8hlWXL/PhmLVW2GXq6hJz1HvCStMpJI2kX8ninkL6lVh1eD+zkVwZ/6gWMnvlx3gjYndXpyB
Xw6opUQl0YGMcy5DpfpkZas35bgsPojbsqC2Y5XLOX6VRZrlzp+d3/C25BKFG8DVWs9/b/4VTswX
g+pgYSTXUUXiNqj7CE8Jhqb2I9sPwVmmyIGh9j7j2dfNRcuBJ1+2g9eo6inDn2LL5B+0WiwaNsqT
G5KT3jGkUN5jcW85stFPmivLeNCZnf8o4OuwhGR5503BNBd/YuXeyuMxZnGwTDAsb4313tlyHQQH
ML0uZObjEAhRPzRr1NseHR3ugI/e40jRKX8W3Pg0TJCDdrkbRzLCpDI2kc8+GJcJCoi8dkfjBmNw
VDwpg0SaYwDwoX/v23/Rzyv25wVQPmVabeMgxMRlwikqodDsatOItkD2M7KRb6KBjSdPQgI5TQ94
pK+x7aLIaelNHNNa8eMuxWeazlKL1Hy0OWMU3HK3tw85EiCJrvzMfWt04WuGXlSykY5p4fmanWwU
kIyenxb+XefcoPjenmvgGwP3Y4jrMtfJcAGlaoXAip+5iOg/LsL5afhrnrh2GeV3gko4/DmpA/5o
rkmQpkt4iF7/umWy3/89MtwTAbdcYh1iHE9fUCinSvELckqa28+e3KkOIZHDP7HABlVfyUPAiNjn
UtOq+6DdqFIrg7n/WLQ2EMrTQclO0i1IoqWtXcw9k0HjqYx7qkYuIM+4yNDIWLuJdlgdC/qLkp1w
OqBbeqOUoD8D6sMjkZqSRJ8arfLzFWf8FC/4lhyFip33iFA6v2UrNXDZiFmoGBxEX+qMqwzKtCff
iQdNg/+eSDLjEtWuwl//xrlgfDOJDrw2VMV0YTHxGDRGeUunWlMoKe2uOBpkZHo9crtmQyY+niOk
wJvBB31B2u+7QQqgAYUO14WJVVP3eE9kJ4cnKLX4med/A8NFOwqVzKSRl0x9yiAYLjxCmjO1lLcG
Jr7myLHbIwWJpBICTLNavwd0gbjZ17/b3byapmv2rs4WuziY0XFX9UkSRbRiVQM6lLXmASeKqcSb
DdJYN8HzP49HeIwaDMn5uGKKj0RWkhx3fOjNI7xXGVL0lHUHZlGQRUDzfmG9Kx8rArZ68nt7hiZE
M4+VsEhAsMI3nTtvHIdopwA2kIj/ZgFpGpMBJe1cDULKe/eNrA2p9MBgMAEK8Vp0cg0YYIwWrCxJ
3Zv2N1crbmqiPjgXfr8Nmci7pz1jBfDVjt2kft31Fj8jPYmQIMnF9oRlbhybcrT94Li2MkQet0bf
6jNYYnGxZtE4Ye2J5CmBhRoATPWFLanOSrvmXMdr0A1qLWT94VRj+Ev/Oib6S/6rhgbo1hs8RJiC
rD0PS1kKYfT/oZ0DY2hfa8EKPr2ZNEwIRNH7MWbd/xJcW3adqPG/Ltcmw9PsjCXTLDOoPLwf6Wvf
goREWilEEmrG50MsaHd1vEmbJmttLQtsWinkh+lir1zuxfPDuXuvDXNai1FVfF7pZBgwuO/3Q/L/
kXV2qKhoYy7/PZtZsion0Y1H8s3dxbL6PAPSrim8L+K9ufl01CGz9Vj70xKbdQhQqhoQYCLLI5BZ
IWxszpgeKbhxL/qqByTiN05neuOSvumQl8RCzEK45AedxwAlmHs3lUZZpXanJhRQEqR6UJNTzt2J
PKdQ4MMaRdIGlsoidFyMydLg3UoXepIHRsNXjvbZuUcYzyDnhDHjhOZ5K4SBAYABk7jvHZQwzYqM
Y3EDo/lA8cfnt48N7Gec7BaAIJEoqOVAbci6+1eu89KN+oOdoIbjlYOaP7l/l3J3qZJFBqQWB7Jf
mCElh76xdgkNKLj5apF8W8ccXiBcePzgTc/uLytG/aPB+UlHlSSQWlj1WPutWIAYe32NJBda42A8
FaRNQwEZo1RBzKAQ/XmitXuOUhrD2tpBDVDe2GCVrBJDjYCvJ++NQdDfNyfmRk52EfY2kBhOHgKx
/GNtwkDKXmrcqjHClf3w/t0q3HkuLLZP9Zw0fM5To5Ty3mM06PbQdZpY9HdMhwAdc6chDwpJ4ItG
4uxCwdNoEvgUXYFZk2/daTZ2KyC3hLssk66pyiIPeC//3QSjwcNV77oNOAE/6YVOmbNxnaPsBSd/
S/427nQq7QRerurRV8EOdCpm+awur9UyOExr9Wb8RiPkcMex00nj9MrvInYHD1UGRaZs8exq/Yvt
Pp2U9x2v42GFOicU99zA3l01JG5KurXHN2ct0nicbyO1w8n3TSFbRqmmBG3rzqGfmVkkfXSYHvTW
xNP53Mse9pCEAn/lDb5NAVZLAa3EK4s3FgyRwVwFpXtGiSnw55ndHpkHMu1/TDrMS6oSwDo8FNq/
Wujuj+1Dxv3qjXEcwVdJwLE6ajynrIfe3tDQt/wM+zjLA3Fn5H24Ee3IltSkzdoCN9G0+186W4V+
hgOLwP4OMXShoGfYgZYVcnHL5KW5/ABaaPsFGS4jVzhdIwBPICoicjtn+YlpHCZqe1nIZUwqJcDZ
9EmirR5kHF/PEUDEEaEO49VKtF5Okg7zmF5VpkVm4qLFsF+EGvoUDvTjLpSZAdZf6foRrKEuQPvH
g5YVVXVvOQHOLY5SmaQS793RABd5FYP6QpiUSKdVeYuWwQ4j5vcbXfbj539yx2hc5MFTgn2IMK88
i9JR/k0ulCEU29WdfeV4rtdINVNoynxWgN6uQu9AQlyJiXpxLrTrfxWeVdMaWaNVrCPf3UVwp0C7
CkNPIeE3TLc1nBmekU9Wed+vE4oNf9gpVagPfBdGMVE0ZZ40RB7rgwKX+8uCvpxmq511frA0hIh8
rfnGBvcLHTqTMKrPb5YqSWmaP5bqas6/GU78Z0uJ7sTGGSX8xL0vbNXQ+ly969zo+FatwB8UxYYo
3UTxHbWx/vK29JwysN3svWvaIy7R4OqqcZ+8LcMBrxTSBJDI3bvIKiMZAvnz8fxx4VaeW3EZ9TIS
t2XeGWkcZZJ+2/L9gD/35lCnmdKbL+hdGGVhFfXCCZ6OII/055KYny+9XRDqQeuepNd8+I9P84gZ
sevdVnhUGPGCGco0Au/nN3s1RLYPvoYGRLj5+omnKWT4Gdvm7EofULkcuRcv0iurQaFr5bVM3S3f
Pb2vKLBPZ48rDR853bvUE1m0nw9ArGB938pmnVJ1LjrckLnNVRx+y5zGngQjoXdxhJjNXV6RDfsv
GQ0LnZIq2lFC1RnM3UPKDzP/Qt0q+rn+6cfjaHmw2wp2RaRi3aaRZr3XesgoQEgnwDYwPSZ5pPFu
CEV+k0UB5SgqP+gL4riOGh8Ux5alCUs7Gx0mPrsW7XTOvkf5mWlafyD3q7VPzUox7w62hgyYVHT9
ky6LuqmZLgGYgY14cE72ds4WmPhB31cWLfMNNObEImQjJDahy5cJqFCVmI0eP47NALh9keoJgT4F
5dIui3OUBIsBqO76qc5DbA1+xX4hyEY/8P49BNZYMDX6aUVgKQsMxa7XkYurUjn6itn1sPXcm+H0
nHKPQhakZ7bd7D1qPRc+cWdSw2WXI0Uew030FCsMFrZstTxIAEINbCXJehgz8AqpBAVebogCLyOt
vGC85Ya0SCD0ZkWQbv83QHZOHeDE+vuCU3JGEDEXuqndYSrsSdTX6zMtIJy4VUMzNpiD+6rSb052
ka3xKnffB1ChwlYLYMs2UVOuIeQaESFcZIIkjRd7ubhv13dnbwpN3oxdDVKVCA113kxaQNPrejdo
QFKJzFTi5re4XostWsQrpSPHP3+8D/OHJTvunEh323yS2ZsZZxIXBKnxUXUc2C/FLmQ5tEA21rAx
DgbgOhSPo5cznYNgDp1VgVOfADRnMW7rAXHHoztvo6SqjW/qkhxggjPDi98zLj0TCUO3zs4qAz8n
AIHsdgHtJMPf21h5r0J35cH/LiiPak33XJHemYlVd2uQ6FxQOVu4P4rj+9noPcxJv2kxRBejnGdW
ZDzzu3y6yr4IyyN41W6b8ePQSmK2CjloH/YMLIP0gc8qvz1zw3BXy09lfxAISX2thWnfNKtMeqYV
S1T936k19JaN4Wxe9ydFpy+OWt1z4DVCUQ50xmlgNQd5Lhemn677iSk95+nyO04TtEQdKS8Jpj39
tJjTOL3LLf8KhqZ5JGFenHqpqPgIuEmSR1Wc8/ABziaM9jyxEP9Ynl0BPkbXSHLVLu80c3CwOv6E
CX1P/OsisMKzgbJ+RUr0a/Bixfr/f7rld63XYWJrkcc/g9zjMWpB9ohcGsfBI2bR28yxdlhtqkXT
dDvCQINDHAbKkKwK6zCiWZZXz705uLZK6KfsCwZx0jIQz44Me3SQW8/pwWlDOV/dsQlA6+D6dlRJ
ZCg1Ja5upDJzjSYH+9GYCnRr5q1iEA54wxoe+94U1Y5TafzJdMJnmWibXD7nx164X2ZD/ycbfdli
3Uqnv2iRpgtP9c+FimU73RZKqdV3H5XmOt2Xjsf/0wFNxCQcZuWGUp/sZ9VbQJ8LpzmFvQNi2cY8
Llg/h5WNy+MrVOwjxBjL04nrMthG7WZ4w6G6I+yASNgE4hFx+6voB6EpkT1FU7QNv+wyftLX6w3C
E6v31BRxv6QAhWqCy5itcgBgNVLtGHsiShbf4BH01J4+dEGfXUfIgoF7deMeWjCH6/GtuqmunmxM
sN1onlLWYCH2MxvtCnZWZt/0mMbye+Dnaig8gZmjpcAiJf9h8OXrP45ho0M8t9pvW7rDsS+ItNA4
r9H+vRhXFCMJZGkvCz5oH1lonnwR6FebNGWvhtZm0KVnsVN/vs8mYbwJJeTlekqpnQrnxrSpOoc+
e7fqqxiMCOtfk8hSFRXPUK/ik+xrKQeriPQ3+9aIGk0/cg/KuUooyIscncQZ/+VMdgsEStWS7as0
hTyJcG7XMYmOEMmNypcwzxKzKyLYxzyucNKq0NEePdO5iKM25uFygqDt5wA8XaeYYsD1KVIs3akN
FpeRJmXny+1SYuWzBTm5j6YDYi/IQncGCIdfohTj05YFXFIiUk6wkv6ZKoPLC2zS4uqvwMEpKXWq
Hf7rLxbeFKFsRyt1IeJIbmJzI8++zZvE7N198/cA2R6IBNmdyQq5vIxb4HgU5MHXXiNC6TWbJtKc
xdwuFFnGwv1I8J2ccZq9inbnfhJs1GA0e2A0c/asn4XEcuz9mSqMI+CSXRTyoisrEB/KDi52mlXF
Sr8Yb6X4IL0a30qDJygwcejQS7OS39/5D38RU9rFtCnSyLne6L8zSQnOShTAE+EmLdPadeQytfyv
VufxC1nfrDXhC74/fR17hQuu9IUlrVHtK3XyywCPUioDUGGyROjV7vbaiDO15OhoXmksrklK1a+r
9Yp1yuGMV/CaBBICNULvbWhBL38lnnvaF3+gD+TlVK8u9p7mjyHg6c5iJGTMmPfYjhY4Cxiv45O3
/a5YFNiPQxx1cfa8fPw8Mt8RQ1bAaMXq+Thpkgcv+Fs0gWmJDGckwfVKogs/DWDWW1elMxGltfOv
4infNAsaURKknnKZIn2TmaSMbJVWXlNFf3dfUvXwzHKjZf6Ejt+91nKG8sI1Am7Y3weyso5WhvxA
N2yCcn/3gK3emDZX9fSxhmTpuh0wCWP+p48P2W4QYCBmgGnA3ZhTFf1QkpxYL9aKS+1TlHNIrfTY
LT1N4qLDdLvPqar+V1yL1Dl/VDhNF7wacfKZrbCEvuNG5TydZ8fQOXl7ZAxSJmifpX+RfAKCOamv
ugR+6NOZYgJKWO/d6USYlC8n8nfHco8V3OSnZbw8g7TG6DpbhvZtn/Ee7t7Dxtlsq2EY6smvvRSW
iCwRz0u0/BHvDgIVeIpiC89cj5LBwmPEW4o6lzCCOkpivv+TsLAVxtsXr9CLt7R0oRZR0nwt+jmL
XzOFn9KB/fjWw+zxhJfJP4WcJe3VURRQPUMV1AumdA3istXNAX8dSKpJszQbH7mpwkkbBFAIme/D
yyEW9LU7k+KiNh07SimEBUqHPlkonlvXwOEg22dxm9ZwAaLdEdVyXjc8Z5eqvHz77DWHuxS8aqFf
uar1Qjzv0wiYuF5kevzLGacvVe3BqRPZWIet0mmBVlujkqM71uaafy96QIqCEEk/VxnYnTcr+isH
IEVUHBDa96se8tzknd92AjvrTFD3MCMz2M2PnYynPnNOQvvQvnaScJSVn0tNkIMTFMZsQU2lWFr8
Rka15vlmHWxWexKk+3IJCLwSfApUTsH6EUEN1ZFIlGUnAIT1TO37VY211N+JtV/P4VIRkdUax5QL
suPOkIFv4UYCThQoRPcJOmOk/Pk6nMN1TyJ6q7ydgPFjh6c5eKRKGrRkQpwUTsFgut1Q/vkSvVsB
bX/gMcyVl5yTH3HwUp6uzobGtvPlZt4zUXWQ562gEtgh8kqToKTQeyO6m69WzxqolIFDRS9C7Tzq
ixv73yx7Hk8ELLQRk0lLtruHaewBs0su2xIqBulC0RCtmxSj6Wn4ABB1kh+V1c9qFY0C87x5szEj
HSKi2K/v3qswO2MHmeUnJRWilsDS/ZyeUcZK3Jm+5j2wMFxEyIhQIzAs6LTuzjcmxjKb+t2IwtUV
L7Tgkr4IQHVWXmnKwmGHiSFM+MdlYtoFT56DplaRa374n76JU2xAqPJmlptMp7NzsH6kapxfCdva
6I6wnSN9O5aNpkhTuzGB4hthky2lPe58KJ5DuBJmHXnLQaScB9HgBUG7O00IRUQcV78TBDfu8l54
DTz4DNsOy+EZ0W5mPQ7lKUM1e9BFL43eQ/glk/S2gaOmiGS1eANZTZ5tIncXwNNPRNYWF3JSrWSR
t51yz/6IMbDNDtS2xE90DwzqXJNhwT6HNcElRWfjSG014URkA/dOtBEsMBRNgVwOipjOnrW2f++f
Ufqjn3UtYz2fnwA5VTaMQNzKshXRJSqa4QPMYdfJqJYc/Qr3jWJmt3Z/+iFNAqW4kCQ4kUpv0lY8
cSSLOsiywoYE0Ss9TO2wsYeBYw9ksvdig28NBH9ucQQ+6yApAyvqDxpR3+tfhtnMJp1JcE6HhuIF
E6uImDewczffkr57hb9He9jRBJvKIuWh0/aQOprvD5YF67wvJOfnrYB7xmbyi/BS0JuIHWAsDN3H
/jc2RzR9AEWGTj1VSfMEHVVQyGtHB3JmAjAzJGkQ/UeAjMRJKDl8gAbM9R8yIzXsBUFKjO7wiDDw
LjTD/1DkwuubPlssiEPZG8eXHXGE8B5ww7TLTImGdoCSi5Px7uhkRLSGabI4reqCwC2VXvHQx5T2
GFO6aJZfssS0gRUCfedmRRf6U7jk5+AlGz44X7HiNn1FHVWAA1qfIlSXy9DeTXL0+XSxcijfdJqa
zdvBAy3FA/wWLm6d2cUNCnp3TGhiTey4aaj00yikwcBbBKdhzlfB4a+7KntvO1yn9eXZkA5ptDOU
rsikaMF4esx3w9I39e1bbFWDuT8v3+5dh1ezeWM+4RTcPcn0P6yIjpGmLyz1hUHykmSbtISSqOkR
cxN0fe5gSKmaZhefqCLu/gklICvYpANT8r/1QNDXoy8aZZiBfZ18617vt6ZvWEy+O1bp0pCD0wcs
CnH7lL5J3NOS69Cb2tW2N/NhhApLeHOiutkG1540A2QdgHS9BFIjsk+ZvL6u4iftsytX0nWXJxei
12yVwPG5kq8qnAJc4jO1TA0ZWWMwmxAo8LWUjQzBjFk3p3bxJNsfc7z8bP/inDCupJpFveQrxBiW
ViTKj7gj7Ssm2lDko3dlQ019o8rOftwK8F5PqLRnwRFjXisWTm68Ayd7hTcXPQZlT5qDBLYqe6LX
J8hU84PJfhXflxEtSVP0GxEDILgxj5vH3/S5W4pr0nEyVvMTuSSNW0jSXty0heUczg7o8b5gPQbO
caQ3p+Y+2gHXlMKzYbsQmjsCl3CYVYcQ9WwPH4tP3mNxmTwJUuEgwYX4CJDE5pbPRw+ZoXaCcjUv
XDFDb2guSry4d5UcNekujeMlWxGwlCSKi3OyKpFKSph5Y0otw61zUgna50cKPo4Ah3KbhEcVt1uJ
xAo++nIEQ/LlvE2KVLnYj4qIsDwRemN3v/pe+b/MaioJw+46k1PPeqsiKUp0NO0aQdvwmxuKAKGR
F+IMQ1tE1dpK4UWRTPNisdT8HGW/Ux87aAPKB06R7gUBmW70xyoqIipY3N6ex/fzlKr6g38cbZPK
hsF2leScYstk7rffb5hSsSl7/Wv1dm7YNs0XZUUZIc2TkLlxXTrAKwctgbSY4eHmYTLk/hH0au29
W73FNgNf9Go0JlA3dso5U9KvrAJr4/iyqUjBU7CKiDFglOpla+0ubrq9lOb/2H/TDeaA5mxZ43zs
HXtxkt0lIGOzuIXbXwj7uOnfIvbW5Le+2oR4cdBbUFUOZ8Fw3oQKe9ZqKtOBYnVFnbfsGI3lXhw1
NtIBx4Fn0332YTpWnKMjwvTyGJvdG5T1ea4m8FrGuB5ipTySLI0qVtD1hRWbmV6mFPhMPCuwXupx
rLXo0j6yblxYcTKRyt0vi1slVURmMXmezI9kmxodqkz6Mu6tBjfX90hJnZroN8HO+nk9dz74OzA0
MCo32k6owKnj6oVPEv6D2qxpPMCytJ2fZEY/ufQlcu1I5BNVS8s8KqCLWm6P/OZDN7P6wlSIsP/1
CRShz9wla7DlXeD/wBKwAxOlvLG6oxffRXxe+ILL8a5ohUsyMH5l+fjgJT9GhCNCp+X5AnpE3Kyn
SO+DaSH2cRzyQi+QzPu/z4FDbcCMDAmD4eF9wTYTetKwtbiEDqzAkG+w0cRMhsguXcQk44wNOERE
hRkrAkvKRZ3onYkpIpZFZUCGbYmZOd/xNKhScGhhTsoVk6jNkVOfzAdQzhYtRkgVNf7oxFjmwwh1
WfN82Hx39m5o0sZ0gqRHMHgEYOdlj2RHMBtqLond5ERFjQdK/L5Fo3k1QcgrruOfeiOmFR3cWz6H
YedAs51wy9jW7X92c1TrjZVAPthvSnuUhTdVZrmQlZy8V2aRQmGRvdrelSVVXOSffj7WsXaYtqXq
knUlQG5Y4zYOQ7MDGYuBAMzVE9/N6gSy+WA4fTdxmWUc8tcNEJ9FhdkiEUozZsUejCryhyNNZbTF
ebuO9174sFTKiRGf4g6qy2K37UggyByu63zLvxbmgMmUL28IrzFlWYmmUihzjjUuG/t8WB01b/NH
khkb5L+PyV+I7KljK1XeMwUIKMY7EMSyqmU0mDSYjgnrSG42goV6FfRkp/2tp5Zi6FxSFpvN0IRX
hL3qdDpZJ3uRA4xy3TY2oYMWw2UdV3IHR4vDdELgcbfwO//qqCrgNjpSkVyS+0NhM0JkxHOzeD1N
kZYRhfUgkNR1nR42VTP4cDdmkSLkO2PBhJs4oYzL+4+c4/1dtda7BAiHIl4tquYsl5sJJpn7p/Uy
F73q6Xmm81EUNZKGzBhEEQWmB4z+hycLJXD2/+au0FxhpqE989sTMdOmhxNq2hmzEV1AW9gq+z4o
6UabXZwHREok4EZT+9vqBUJcY3+pb2qYBBKklYErSH9UsswqNOcLTJMAko/fIyNaiJHrRd8s1Adx
wfHaYC0j5/NxxgSAiE7L+frf25rVdXijTgCixgeOfWsykrQW5M26a6eX+nbnzOqre/SpIaEhQW6o
K7fDL7j2eoL5gc1YQsNmbkgM2IH0otIXCHFlPmubkqk3mEteZbFL6CFcN+XijYx4JJqJi0C5ePdo
pK+MefJkxt2RZfxFRE9Gs3/plRAwv1hQ2vmkb1up/MidJz1Z8EQK9jEX9KbjnXPpRzFKvdY10q/t
2mS2Et6ugXsHCX011y5LIBUT6WVONkN5SGD6wLttOrT4+kuI0t7db67lm2WF3E8/24psTCNFCoc3
cBmdhxeZqVuV4tIcqQyUweRANRVOf3PtowAA/uMH0z4P0t0u4tmRne0hYIFGE69ycmiHMAkTF+l/
hYcp7/uxSdxJF1F4C+MxgVgBIGPfFgWMwWgR7kwc7x1L4rTGjPBLUx/kaBFx3/ZpNJahgyefSbGt
DyAN8aTaxokaGSpi9mmo7ARrXhTM9TtMMrAb6x8ztb9wNRW+Tp35VRNmkSykUc7I14Yu0FuzKoV0
/ZN3W7tgL8TMaDGTMST5n1Rni3UK9pif5L8iNlEXltYpNkHJMLV6WwsCujaevHJrkk94RrPHqda6
cb9KI4UB1RAiwDM02cnNxDjwYC3BVNDgihfLfqKtUfhuKQYFwlEJ3yFzDFm5OZdorvuPVnFwSVG/
/aMjxU5k61k15/8vqM2uC33H/NRpziqnkj3aHHw6xZWZsSTtp6wb01lG5wwxQoRW21/xmUX1IEB+
O4PDQvh+ybFYVY/WVOS6V84fYVKE3IGBaXNT8/DO5NSZVZctHtCNnPRNsFIyOIVeEDWwtoBgR3Bx
T1qGdk37ZWoD9/wTLvuFL/J5cQpZkHLnUNs37RAOksgzyE4Z6ysMirZ09eNN+tMkt5MDDVliGrDA
uL1EmA/8PmmRKUqHxw40KNFEuSQckz6PbLffuDu1mIgv52/ceD5erSh8gkLqbExc09tPK9+rQ+P8
4i9btwwrAdP+itXvwsWrbgYOaZBcveQeluLOrMBGYmFSaDGDihZjqjGP7jeQP1QuVHyuSIhkPhiT
hNlk3MjOvYkFicT8BA6UtDepfnsQOslvGLdOgWNeW9rJwzUTuVjJTc/TIhwhzAbjKeLmVXVex6Tz
v5Y1FPClNrJ3PrDeLf224apZnwLEKMTiF3obVu4QBJavN1JU+pGteWs5p65Az0hHTHnLLFSQWABW
AzI81iJPgpa3ZM2PUmC2IqsHtizb+UO21o6RgkFUsvlxN4gfOao1dZUoX6irMkbUqaZbsOz5mpNQ
iaqCfLB330Df4Blgoh6E0BsA1BknY/VI3NgE0LTyLeu/xNMD2DL1FfRVOixqOuFFOnl58ryVvqYf
XkEKkL/n+uP6XDKWw1nW/VWELmoYYqb/5mLtQ9vM5H6PZt/2mvw82bYLoRVWTWviJv6uWqB8ZhDd
lZaGjVXFhc2iewivL+W11XRZJhJpbBj986oChCDLWXhBmG308ZtRkTqHehTI5gF3mjdkS8Gu76/i
QBG92yyppTvS5X9aRDprVMeiEESGlevpF2M/+QC4irl0K3cCj8pOlImQAFNjPexWs3Ru3VIdeFk2
8Z+8oS/JynskFIzYIf3JBtW6AWa+czBSJzeUllTlccYMkUyf4BWBjkjPgwF/5cvxkaqLqORCJFa4
YfpczT4fpTU6peMEoBIIqM81vwoPdv+CxJuabPJZKkvGtZ0XyJ1hYGWzSaguedJCET0FL9/4Xt/i
ugl9bF913Z13toKyTdET0A5m6GzCP14e/wguWOIvPNIZCMf9Aj8YJ+PxqWKmseJ7FxxZAP4RmMCm
6nBZjqAL+53k+J5HLzUabD9GLY8kDTWk4Yz3imtW6y3fseRhWotKfS8ui3kJrjVJuBDqAfiQU4Uk
5/WLExeUx6gHmBF2TFtReyA9fkz+HfLAVUJuuSULZelkUJwDCrQD72TDY7YlJ65vlJ4vleqmTWYb
pEltUYS92rKtu+lYvNPGLsTLKGd1jXRz3M7kxdK4Q7X9z+BBnaZQEFEyvnvtBrtyeWaoTQNKF+m9
yXEeUY9y2tj4s2o7b5w8Aeb+cQldyvkqvddRor9S7iW/Yja1yxsTtUAgRFfk/qTa23Jdmv/pzVeR
X1BeXNjXClgHCtAFohVtZYbDJFKz/mdMZzJ45C4rQY+LgagvSgr+Ri2P/WYDitRIt5PkInrVWOp0
Mox+kNZd+QPqwnRs0GCpth2rTduiOOm6CCeu1p6SXv021rqdouv3wRD63ALnuoNg3AP1CYL9wuLE
qmgUHd6GSHKzh7x97OfDuvPI5Xkzk0NCS7H2emVh715wi82Fl92H2873A54yF39lvTEwwuDuMFSa
3GBLrApYVQPhX9bhzVHOX4rR3JB0Ks5fKfC5AtZzTe4ml2dVTKgFMkXPYsm2eRd2pc+RcClrpDmE
rjbKrzc7kh5O0Og4nGkUxvrlmIg+MeGrhY0WR6Pub+afW8b84HBlqK/HmECGZz6hS07dFB9Lyhnf
hzcM8vQ+gI8/wELnUZqXNlfqCy+jNwXp0zWtguyCwlsp8jXaucZWDGqRD8wKu9v1og4u4TJlYfTS
/OsX4Xkea49/Gxds6G4Inmz51dbmMABq8YK9UZnTbkrCBD00abyhcOm0c28SeC7dTK0u++xdHj56
FVj4W5eHtDEWw+l8eD0SR6PSVcuAEo8AEZaep3o2l9vhmaTLftAP9OkQ59jSTBOyd2j+LCWDRBXM
3p8ahsJCJY0oLDeKDluL+E6ZEi1tr59SqqicfeDaWLAfsDiWciqU2fJN9LB99dq6Og4MZEEKgZNj
urfag7IQXhPSf9bqvHoj39DJ/OARL+T58z4eb6za36acIpJ+e1a82bErh+5uXIqfQaQsP8QMJwol
8aQGwnzg6tXcyVhcSZnlNKCmU3G7Vz17SttkoktktE+Iy98oYtpQ++jEarAsXCM9jp2FJLd24KuC
6U/U7XSxF8V92JYSIFHwurpEodVWZ1bfee7fYgM7KkVRldOWS8B9zXKBk4X2cZM0Lb3Cg2BUVXV8
A0vTrz+18Nr15ARLQwL1Z7Gat41tIphjD7tfDCrwlFczrqgTy24q1BxueP63ykyOC1puLjEX+QAJ
c8I48ctEon6HUK/YtjzeJ0P/J14XtjQj1CWksVJxfU6aWigr52GXZyAVORBBdTwgB8nWYOM1kKo3
iNrY9h9aKJypIAdsZJ2WlTN+YpiMZdFyO2QuT2mHKeDvxnF8/pVPi/06fwnntp6edWQ/d7SozU6U
UqVwpNKqzXSF3pLV7WomO5eJH7FJUltTE8AfusNMgy118j+0USdTTGzY8jImMMftfDEmP1xdSOVO
LEkQVUMHs0kWXxUvBx+z99xxruWV0X+RTPfH++61oV4tUnTCED+a2f+qtX1y+RN20TAGf3806EB9
h/HrAiu/506C6d4oGZmTjwIFNOD9JQQfoBJ/m1nR7gz9snVseBPWEio5UHEDXtBrDyX+YhcI9E9n
Mc2Yb49guOt9trbAiicVSA/fRv4C40LDd4rnHz8G+qWvuq/Dx6/Q7SEYskoGXDFc8CfRAZF3GiRk
BEzZCbAK39Gsq3AX9dvfgu3NSSujPYG0ByGGli9awQ45fE5s+Yb4OitpDIdKAbt0QlONo/iWxoX4
fbT+T/lFe9gpJ8F5ssh0ZkhfS/ckqyo/IFBfVopqEbsEL24NDkR2T21N/aKQpAUJjCV3GgAYd4V0
OpveF3roHQp6TTm9jf/nVVA3le3ENy8t9jTNDAh/vnrA19kZDaagH1BGJJzSzmGTAVoNDOGAdn2D
xwABsxaQmamupBf8wJGZQXRhlkfvQeKbheQbc/B7c70ayAtHXlFMwLnuseC6d9VTztdOm3nwUAuz
UzaTpBOTb7szsGG9s4xyurIY5DZxTvTYVbariJLSV+ukykh7zs0T4XS/Amc/u6Unv0Mxjb/Pvhn0
3OM5HE8M8CyVseuUl//OAclxVgZr+BsFpLEMS42DwS4FK6FqH4Zpgl4lw6PueWSkApmuvFaN+qay
nGD5FLZVs2PajEYn+ecaQQ+NyhxxZsBb3l2dnbLN6PNt9Q02B52XbLBJWTu2Q8Mcj3gCIWEaAmjk
Mdoc8h71dRHUSTRMFMaQwMQt59n1GPXTevs2P/mJEDicoScUnvTwmtpPNmTxgAnRqlrDFvLDAc0C
ftF7sgJ8I46ZTrONP7rLPjl22PpVRidnZCkpuiUp4LnaGqtaWLa7dmgVYRjxaUluAtp52mKjTKZW
JQY2OHREjlD48Pz5i9ENPxbSMhaa/DouQd7aoibErvykVfQX6Hr2q5e+ZyFLDVod/r3TA71dXnWd
YjLX/MIUORvLgvJB+T+8wpuicSgjXajEQl+5Ad5ettB7nyHC7Mt1Kk578XBQ9DkIio6vmudxUmXZ
UvKpipmRUoK7SagnXQb6qiIZqaYax2ONk+kangq3YQjewcS2AfLJeF+d17DhC7DKcIyPPpVEL5h9
95C4cUtUd+BAN59ny7J9NxFRG79dzBx0sAzCmpO0QfLoNVWamWPojANfiSmEjSsny8MezmtJ+SSy
c67AhtxeecE3LsW+nm1P3lTKJmLNxLGqeKm8NSSGFnxGLt3QKxNHTUpvTVel4pPmOYVOR7T/lGiF
hXtcc2l5/+9HtswiKtBKYPtE9loCNNaRqM94edSn0H6euSWhDSr60gLiIOl0QxiseDx8fNEOfAnR
auGKE45FSYR++pWi4vCvGUShyI/5+0JvYqq29NUg7xZqMQkRvw9BNDOTwe7y5iLtnzgvQLEg+5n/
/sq1ruYEY8ylTOnWl8aZEy2pe3aKCmr/6joSQdyPLDB0/GTaakd4sLSS3zGU/Y7lxJsQJ1IOWWLq
sNgDrGmwInlnL9yWhcrT/Fp7DKclXLKSE4Yi8lXxsfsf5qn23qVelV3Bj0Z/Yn5q7Q7nuYJs+dCY
eXwcFEbJ9iigRTWNw3Gg6j6s4bb3YdFf5LP6QN+Sb2878dgY3MlYS4iigvWldcn4Iqub4NbBMpWd
dDZJJ+0+EgvHDdXwt9Vf466Y1cBR2PougsEYcRHhKYR2wo9eVHS0Irh7zDDuFDXJrF3z9lFuDvqq
koYBljkEUqL05kMkSrb/yNUAlLvCXBJeanOgPtn5YEyA2Mhlo3Aohc0TcrWMecTrarzMmKgNryE6
4onKsBZ3OWBYNyLFCUbTylFgMVjfiSwsm0bSZ00gXE515kjpCsEaZ9eKu+tW8VFxRLwh7dcn3NyW
JpPKnh9iKjThxdOAN7xhsg5ubeyQKVUJIrsKAjXMlGflNkQsgzb/yFU1OjkVMO0yL8znv76ZgPaN
ONxSRK30joqBNZ2IJb3vKFS8RWsURDyDINI750KsLuFIO/18RMwzjuGT6jKMNI+IdGjwPPKtJNGk
N23ZiK0TwYqZGS2uWlX088syLBTsvDYtlImzwk0vpX/Xc/s28/RhUp9yV8ICvncJPGaSuhfn4xfa
G6QI/PvhJNpTU1i7iRcSZoDrY8gvzZC9FC+NmW1vpVVehn10i8K8EmHcgNNMvXE+P8aZDxfsriS9
5sEVisSM4TrIgs5WQ+cg1rZl2ynb6W+FcsxMUX5HR+HElHKl0hNXoarGE7dZyKjUA/hpvqWnXrGo
3KyJ0foV4Fi0YHdRSgYlFFxtN2oTVtHvSgpMp51JSY7iksUu6R4ONsNYGHQtu9I/K94X5mVubYMA
6Wnq4wWPTZHRdsf6bMGfTBPWSLoEyBsbdjEmr0XnynPXWuNCWeJ2S2HuWWJ75aXnPmKn5vZAlPi7
JVfjJU+eIX+OiP3IkiJ/RyhLkM3/K7xaXI8C0E74ItvnhQlikUsy81BpR9O8rlf/INky824SSZUB
gI7dOSWVk9gYthadSuoSqI1ToNoism/ilKyPTp+Q64SSTirKKgxkYFSNBgcuVYXhOblOgy2X/RmT
4VRyC8u6DN2kcgZvtgT7dIynJQmpLqrUKu52SgBbbWtD5SN9ZO/UzInTw1KhDgQI+HEcYSBwJS05
1hroQNUGMgjFvQ7YsPShSizyIa/Qxo01QH/X1ZvrTvRAN0HkhojdjkO1VFQtS3WhmSgWEdt78w4y
kyNn4OtdzRIcaJBLOg5PfwddIoDIC0lgPx/Ey+xjvifWzmHzPjUyesEUp/gVYtNjBVWRTFG+i17q
qI1QQxqWmAhC/XQB1XZC21Ztb4SpkuNm0NFxYYjNfAbsLpzERxoroE1Qz6MyPGFka0dDxcq3YPdr
C6flGCD4tttCoouBCmYJjTiS5HNF98SuheTez7PWhq7ood/pWhLmw4b5apx4lC3Df/WeAULV3jOt
UObKT5OJahFEZy285KWGEii9ICP42OC015W0nruOhubZXXer+xpLvamYqjLcFlndX+hFmqdlmbHR
vW1kMCdo+dXXv15DOAUvQbOCHE3ydmRX5evyXNxoCtAgzgb6Omgkr9ByItBda2Ge1Q1WSubl6r5i
mvScMo5+ADNuJ9Ir3Nf8WbG3jGoNZKZnxit7OV/rW2MVDJwD3j/JihQ08mhik60t/nmVG9Bf0FhW
2ZdwZTp4Qrgh3hLLG8Hih8+2IpMrQwswYeIN98VAFA0TEfG5S62zLcWTvttWTXsFhBmplBc3fv8+
iipBhDPpwASQRRGwNDA6Bh/yuoCOk0WQnS9XuwMnvjfo+gkeWreSR356xwvPbsvvX1QjEoFsqohp
q5K+1rArdpYU7aIO53qC6nCKFXlf2iSoxmAsvD+d65dg3jgrYLJlgfMUcm+6BB+Av8mpeGu+1QuX
BoQMONVghd6nN1KLyD665QLcJRkF9SAvhTMM4cfvhMgb3/Lf6vea3jCZLxlxAAJiJN3X/9EjHEPR
34sf8WXJciZBoiX+6G4cf9S30racb77VQQXRp2DoBDHLTh37vy3jIw+kqoXVMrUpchU6CiYNyYz0
OUhIgI9qFYkfGIlh1qFYMBBzF6BGL4gt9vN/jBIYCPKX+gtismo5O4Pb7qrd/C146y6TbFH272ml
QtoCQNkw5C40UB92D5O5GMocNEOAEz4sKkfMR2xDCZx6zzcZLAAlrsNQ2yVdQ4oH3LIZPAeEqbph
jInxnduBrcJ/POpXwzOLrZmK9n3ffeap8ve82iqWxkZeVARn9dQRVayHdrl4nzaSctPiEuIDKKVD
dlnow0OQJMnRmyYfzSWDMfQcVdY5w/WKSfJxPV26o2HDpXJFEMzJB3zts5MDh0hQfN6WeXDrAoW6
WqenQBQw90hADqBCb3CHYfcqWqtsDrFODBjbXuFGq1tINSmHnTIw0b5q/50q/30cGNk99QmlzvTA
a/NpYsaVy4AF9kft0QL364RorpzHOPXkV0wOCly0GT1q0A6rqzBoz/y/y53Y2zIe09obv7wqJqL6
DDTlai/+5spkzzxd50fmQCnYDmHzwDEJvhFMm5w7EsM7/OkXXPJ67yxPaPQVUROKiE+h1Dg/vHV6
VtwPD0oJxdE+iBRtMf276n5r5h6o2pJ4AXwyfMnyhr5W3yXmIcMKyHK2ZE1nzFwpZ1RM5nzorD69
PJ+sjkjdB8Rul6EjVQ4ncOZvP3CAWjcB5YzAfnlbjlbPhI7jxlGUCUQrHJZICWtTHUmGrqRdx7wt
Z5ugQ9AmUZ52yUsKfWtRugGLQ3FGhIef3keDJfvi127fd6uPMbgTa6Gdw13T6S4PhmO92qZGHvbg
50BNoEEiEgG5wAcPZ8r3LoSK1Vtj6UpKpz02Rcf77LjhjYKX4oaFy7fHVj3f92ind+LtCaBxBetk
IBqug2bD/6D84rY1X6eZaolrn7b5kKBsTDtMYM+VC8gagQLltGHFfPDRVoDQ0U1ojdxFJg1on+ba
ClQE5oxBIkeEXRnsdFAtW5nuhMRkiw/23bTMoZIxThsEnv0NaEZns/y222Fnjcw7BjzyDkie9BY+
rNTh/NzhB6zJwSPaoFxW39oSKai0+t8H8wnVNnLl30LmXuMzT/tJafuegGqMRKfGEylw7NyWgAS2
1SJGp+vv/zQ05CYXGCeAa2/xowbco84jhtmQvPiE2JiCCBHuCjPLVxCHC3MjFko9ROvZhsDQ9nV+
oFYFVJkxfz4Ufi1ozC7tqF3Zqpblp/1qy5rtx5xGBevJyAREeeIwPMYb/9AArlo+XYb2kncqIp6O
Ljm05E2wecqEH2NtUhRdmrCvVh9ey+lZklIW1sHwBf2j5k0gsg9zItaOFpMGKtqHXgtYe4Xva4VL
WwePtR+ybTFtkajaGageltwRy2n+joNKcgmzxHSJvuZggPVvz35YUSdyMEzxlx9A8ynitMutrGEo
dr40S6IbFnNTqtkdlxCDjHH94h7xe1gAXoylVr5Rb3iCiM0cEtf8bXIgJ5tlWzGPsprqnG1xlrFr
Zb0GzGGFC0xSDmwhpWO8dFUSzPD4Pf5EceZnTMW5oWHkYWne6vG8EHTxtoqlG1A7FJO4sTnAZ3sr
9Ca5x67W8fpggrO5NbpWB1ej/viUHNIQMnKGZCVRxI8a14NE6b0s5rYa/+rJznaYCee9FSUrApFW
pZW4kGHgEodmPr4iby8e1n4u6mzjDPMgRclQvImbfa4PcEVSfr4hezPrH2dBgxnshFVq9ddAvXDg
c8Tns5FBwIXM7pwWGstzftJt5WY2t6mqbHwcrhv6d4RfpxzKzAwueAgM0oVC4WOZivrJ6v/ZSVvS
wcds1KIm9sCMblMh9a5wtorHipTUP2svL8VGThE190KZp8o9VL59AdDWOWcVH8yN29Bzo9feUY+e
COntlHwJmGKFPS0hJkeSNjlD866R77Zruy/263LTPX5h1eqcxKIWz5UZB6pMgXzP6dAr+wCIj9BA
MDh385d2badihdcldiJC2eAPiNRqJBkAO6VrbfuEGy29IdkxCXqZIgHD7vkn4jVEz3hGjmqBN4u4
YDcO8+eXkGpjlzriLCS/gVMpOEgzcR2HaH5xDjjeaB1qGhF9hTI3DSKV2C1UbA/32WKDM92bSVPm
gotuRjuDDrnhYJAHU0iYxRI18wSfupHBOt9F7+mzljrehTNo3hpCFJOSNQKKo6z3/4OftyZkVpwU
ZeyTHJZuZyDC933PpsRYdaw10QpAucbRU+Hwx+Sg6TYhtY/yIZBt0uVqFxIYmXn/SiH0DFhqDtaz
B3rlAiKrOYafYlERYERoTrUBswwjecH+Y94xmnBMnSQgkUIESopdoBsgQ1oVKlWWsjSGDlvEysIY
osX77RkgeRqngWWMAF9RyAqp4NQ1RLKdrI960uY80kdLPZiERjY94gw85BlWgfpKox96CXkp9PC+
ydroZgWPhYiHyWDtvXLYSKmewnU2aYJ2H0UNiLOEwdQsLpevJPj/3OAkiONnA2fwSkdF93cx89Ry
M7XocFRs+woeNRigbD55x9QW5nCrPGodk+YOeiS++SUrNv0rE8ZU34sR+cgLVUeoDW4S8UqORVOE
miGicX3q0dduTID4JO3BQCqMym0FvWRRnBLsJrgOYMp/qL6BjWARGe8eMb8aZlOfRHqQVGJOJRWQ
PH/9yTOoozqo077RLbQM+dydvHYK5nAN0HXagLKjjqHX/4u/5t8UzUVuXTClU2/7Vq16wOwZZRzY
BSvek0zgMaQJHZglh8EVgy5igW2b8mOyNO8WVKO51GC4W8oDIuxq/r6dKWgVHuX55eNZF9lEiGgL
lu7J0X0t+GKODrQk8WCE3i+S4DrNJeTF8MX2KBFwMNwmbIfb0EiFF/5snSUv4Oz7UkALnw+TRG4p
8RhWgLjkC90ZCcR4AzwhEG/ucLPdnJrDzwbpgxPSD6L7Hyu/OIXnp2ARLNv5n7p+lFPk8BiXJexf
54KaK1qkcphC9U3kpgcW4136UlE3kUH+HUFyuSx4a3+7sIQ5T33+nhmGrmq7PPkthFb9Rp21/tMD
KkN6Die7FSvvwbaK6QQ2atiXLjiC55xCRdKGvWWAxvhlYyynmjPdmT+y5nxP0htxBFyiboaofJYY
En5FJ1GsW7T2N3Dm8ACEoD9DY7rnskOYj8JfvZaFlPXjTmTw9x0PbDugLbWI7pwSaSxArBERzh3T
+hozPj+TeKtbj+YcXrUKvXo63mzB9AUmpRPeQFk1jvd7j3UUjCHvGCXDzGdbfbJpzDaQAvWDwZIN
vg4BW8l4ino7Th61Itc3LrrypLq+s0uHLznPiNJzpyqWL31Ovs36Jwka0rGg7HBI4t1AEyPAgcMk
loy+X01Rt4Fl7pwsQv8ksdYJvmOyJ9OpIifDt5zOtNEfoqvm1Wx1Q+ydxSYfP5VgZ3R5HJEPtFMg
dvriW4NcoK3rUtsK+PmluwUjfrgQJjuVf+1QFfIOaSQBaR4BqjFNSUgGLfl2V6WRwGpdYTUMKUjj
lkrYoDn42EgXJbzJ3KVoDnBL4a3XO1+774u8Xvc6R6skE8eKMiQ1ONYXhgGUcFHx3ubI9tOcMnkE
3cuu6notzfSEAkxGpiXSyNY/LYsjgeWEQ0lGXaZHTL4lkKoAemOY/FgZs9bzoQlrr98FnpN2tEE1
/dCT/mNnISWD7zsPSx5Fr61tPxZhEaBob0GCSONBTqFRy7dJZNgtQ8NHoh5ZS9psH25Rbq1sVdlp
LKaU3pW1OK1P5l19h1n27YWJe/stQSoYbSMKlQUB3DmaSvk5UDQKvt2sW+Y4txxi4ySKVds93hix
HEMP8tkpRy5F4DPvDSukL6vQJc6HLl/GzPC0z8FPO2FrMyEYFT3UkSDCbzkQIejTqXIh43M+cTCs
ZisI9sHDf7dQtbYxS43yGxDLZWNR0A3PxGV4uMEsDJ8x4LgUyWSmIDLvDH5C3v1bsuMTz1mBu9E4
msVpAAKzTEYiKUZxn/NthdelgPJX1icCv95LMk5BniXEPDMy850MKrc8lJv12t3wOmLyLSexfSwi
grSEXx0FSzSPSXai96onaUM7u/KTeWbjzNwe1/qlu06ZNwFRwb85xgpAxarBNwgBEy6/vieQ/ypC
klFxlx+9u0qSKQhUtulB5HYE+lQimQraNOSZuNVzjb+OFdEhy34s/vtU67VesWUvq817WMyIpi+H
VSi3RUhssHRXRuz5DuBkELcJhvWdeBX+h0w0bEd6pSawMp5Xfcuc2mZ0sUxfSiyc3FDI9Nw3SR+Y
CvmYlW25QX6MojyLLgdXq85r5XpMbhMY+O+cRgQdwVg2anyk+BpBDGKy8PDNNFerHj93Z5Z6eGTA
4gCPv6bPipcUPTcUJ3iM2dxPVexAxC+RXTl0kOfU/JFIxtMN/NSpco7C7/dRoSgrfqVg/y8uTrpY
fhODTwO45VkP8EbkRzgqeBAYo4yX8sztJDcBc5zH4jxyaksdTfx2dri650bNWYUtWWlo1WG5gitX
gLqtrCnhFdprZH/TYgU8+7d1aQkvbPlEW11FSbRrHWhUTZHlWmJrYaTDi3CxPU4dyN9TPLlbhRFf
qb+y/qs2g/A+LCHVHTbI5q1hO7UdbbuLcoFc7L8OMsc6LcEtFh5P0bwIOSp5uiaEO+tga3j/CvIl
4Y+pex9U74cw1ZJU2I6c/B8CanrzI8t4a1SR2rUFZA8zo1kB1ZtB/nivX4fSL2fLUKHEcXyhfHyk
AjveDyr9qV1tE1ahpuFeNx3E94MUxBUA8YN6mdwZoyzQsYgeB59GgAgORK1tdNSMSyVbRLvdjDrA
8QOZQJrfaehv4egtD4VqZKawI51AVwleWgn2+Utm3oDSIoy6Dg6AB715x+SEvCetIDxWzxolsAIQ
VNApHvMKrIfeHLAdqFsatjqIDddEvSEyL+aPjLTd5NpM3WoWnWdekdRTmg2Fujn8QVyGbHAF2s+2
p3JpHrWDS549oq5M4YoUvBAIEAhFDn9plh96E18Fh039Jezis01caN6QUS6zsRHodxTmnDhqSq1u
I6F3f0Fp5gFm9zMe1A0PFqLn34IfCbaIrBXbv+8fwFjckuAputYtu4af6U1ragdsTqW69haiXSHU
g644YIZRN99YKnLPNpGuMOIbveIgb0v2g4xnk1m0771cXcbVs7lTTGMlRAeQbvsldEf9aIoDdjcR
1E5L6lBMEG5bV1LaIlWhgkAh092L0qHF/unS9xm8HYMZpSrvfRiGPljn0m37c7vVKetHOemhCAwm
tuiix+mhoytzrnyYluk5BuEGZuoWeCmXir0M1t6+oEKWoq9ntcNIfM93DS5s6V7DQhQroTQ9QqEP
IzT5cnlRwqMzFzpRz1lLiO93V/eqSP3romfQETibF1exC8fFN3LSMfGnqoRd3oJKjw9I4tBsoNtW
yP0BSi6aCsv8Q3vaG79DU8gnycCWsWaTMXa9++t+3a+H/7YIFQEQL2rvAOtdpRns5M7iD2a90QUC
sz4aHqT4oylLkRfYEME/crkUir5Qd3Ez8tbN0r3I3GfyHJR7YUq6SUlc14IKJ4fReTbEhicpynrZ
1mM0iOhiLiaci5hp/KVZ9XdDrhAk4/+DId9c7JKRdErcFbIjeLLhhQnAdt6HQHfleyKiX7Ov5Ybf
T+JBXRnICIS/xbmnoFpCtI3OqpzQMbOmAjrwYzK/8vOeqMKFoPoeoxoCZSNjZvt3vQKEs1Ka6ZsK
iOpPE292xNQEHvLTf/iVuTtPVkzJy0sJ6S4pj1TDY+9hi3sSZKPCcOTDEw+mm5fW42+XxB/ramca
GNX7x5X1cU+wVoUTkTOk5UoR0ctxgPpHVxGaRQhkDKay5u5CVnsRbeKH7pFF61ZB5W3d7h1pmyCn
V5JF5VXZp553b4d63XzhSZ4BgYP45MzOu9kg6QJoNehPiHn6E/Pyc7kDhefwwpN6qX79WC5ahuVp
M28n14OgZZHLcmTr9BIX5ytEY9tXTN4JF3ScxIX20RhXxrhTL8F63pOYs1sXQ4y0iEoHV4/MukX+
dDw/vKIUM88PeH5XMFC2VFyJn6pR/+h9IuQax1TueBhpB+e6LfZqiAfBRjLihM18nrdlx/9+TXyM
ozOpCuJIOny+YFw/LBumnPo/IsoHSttzmpOdCXwsaqb10hVDiwF4NIUDUTy1jDIWRNpOemb1VEzd
i04tumr3Ea21VrwQa+nZf5uyxYVfaaN4BG+VYLrR8tR1AWBEFpNghJp/FS29C+/jBT3v5d2B/3dq
0vhhXo+a4im6lxa/rhk2jT8FhFJKO0N5lnSF2vCIbTW3llYLiyQ632U10ul3XObTyu1xSbNt1OXe
S3EkvU1ZITPMCzwsfVj0YdzhmKqwAPk6rlXLXOluz5JpHDM84j1A1/svPawrImuQKkrqnNN11BTc
/rchY9Xx+Kp7Sm5AZoBCkVdM5xEnfifRxoWVV9lYskcEBlElfxuhfN8UW3WdCPaVYgv4IvuZm9mV
XzfGbaP9MVt/+VPeONC0WJZ5Tni7ogNUvFrg3QAmm67gw7kZMX38iVpurmin2YwVFwsE9V/ZRInl
kW3NVVkRQOwgW5mMg/KIZlHewOLaZ/+D87MFu7HTDRRbgu/Fvqz9VoJM4r9lqDkb/MKk8C6K6/O4
7ki0xRITRbfAhW1jmMWat0+GZSGLW6dHqCZfcecP1AwJ4Hcuqk2DQWtRUM7XzgNmAaY0TzYlWTJk
5l+m/LTuTCmmNkCv59QJLoL7Cmyyv1QygxDQtZeqhGWr4CIpCPmq4pZF2owjhEXD2uBTft2NZijB
6j1P16+8GAPc6D+ZxUyyY+igLiLHETMXrknl6G3WcSAE7DwZSTYrr8z+qv56eGKku1T3JgYnqJ1I
7IasG3sAbHTQteBLtJDIqIt82cWRPiKTCWE5nom00CufnUFqmumYD7ewaSuhMys6IBH6M9/Ns+gy
Uu3QRBksTK/OsRjz0KM5HbwhfiMdfrv8oWFNmGz7UIGziupAanCy5kAZAFNGjZtLU8J3NqOQeB2Y
NuPqqTxnPzGdU+qLSzv0Jf+wfPqbboTwdfV3AgTHrnOV6Y3EqFG84gchCX+1zcYcsJ9+TKVKILnY
uAi+awZturOhvTKd2V7LhxruQTiEJmAPt8giCIpnzwSV8+p7N5aznY+YsFx+W+lLaEBa7673VDyT
Ha2S6obHyKAcDRpCV4KYXfmeG57+pIBlZK7U9vS8mOun1B7V2YkNz1DLk4Sjt65kbdM20WeyFgRU
Hr3aD581tdR/+rkYTlVIvvLiDZCVgJgrGVID9QFuC/3mwiRVPSj9KU3NrcWqckLlR5/dxmWYjsoa
c22M7mkkG1KwvloIoeEVSOrZYtfCOo/rB1iu3YQDOeOMLmDXSpdfl8tB7qCA+eMKmkZKcoTS4BG8
m0KbIbYKrAWyo9IPhvgU44uokwitb6AbklDyLBdf0op1N3yCJlcdHuXXjDwT2jmkbtZYXcGkvCeZ
UXOol8TNgg34uLXNAT5CtjnaszmyvRKnYjlcUeux9/v8Mx+IZz+3qF9v0EbNCO11/bfaGovsHvyg
jw7OjGDFUB9N6V911AJkQtkciAV3JhkW8bxY0TgDjCF/l0toDPaUDYX339Q3hat/KaDrK88fISR5
6e9d+a1YoOCF+vNOxijD+T/kiEXEq9IRniT00IDNm7N1u2L3DNEvsxywIqCXR/USYi0WMrSb1MYT
L2JoTu2zWXU78anZdUBgW5tTJRd5ooB/GqGPn9whHivNS80vZZk/Rn+xkTOma0KSdUnbNo9mXSKU
7NaBM5/pAmU4U0bw1lT5S8zh239/n+tO15lntD80pdnTz8RrPkGnPXEOlRvja+ZeUYngzYDj7lhG
v1g2C7f4ZP9EnQ5lP93QB/WwceyJ0ljWTvyoYwBwLSHk2XfGCH6NGVLuF6wgptcqIOcysIRnYoS4
Mrj/AO799z1gk85a80NU/A3W73tOfEh1xLgmj6COjBS+S/bdnSmSbY7D85smrQyXCnKNKy82KOdc
MY2JPtFdoKnmHsQq3MQzUhZpZvDh34Qp/w6lpOYbijLcZBMnCGIMmv7SrWrsbuj9a/SCHm8W5aBH
QVgl/5khmyZHAG8GzCNpliAqX2BYFfMRM4oo2AJXf8iQrljJUSjrsmiLVo0muTYeEOZ2/Hf2bSz8
m+JU1eLG8wdLNqW2qA+It9CCLZ8eQizUCKOxM20HSREXZ9Xvtv4IpB9QmvSI4Wv7Jn3tdwdngzgd
MTlOS1hmdyVkLAguSemDrQhbQo5cxgz64GR6hnReoeZhsZ5rgHLDZX0gOmPLNV/vRpgZy4Zn8aXe
rovgf/9MK99rLfFQ4IXwXZMJCQBcCU+fa18xeNHrFL+Duvo2R0oepOV8QJZnipEVevu85ApyJdRJ
jJfgcszfJHTrHaSk0c/qs7uo8j9sJP5E/DzzitCNLQsBbwgmPkQPxx4gkwjAI44drs6k4+BxFIov
ukIuKgi5j4kedPxl3SHBKizlMvjKLhouyFqil/+5lnlhG62vyEBtXv3DnbMO6aQ8b9f0I26TXSJB
WC0kA5GHKuKAGtPcXcjiH0OT5Acfvi/GQOc85YzYDst0IXp8yThfHTsIaGLuvOIqEYWLe4IOJICo
MTt7cER91dsJxVWCMG1Qgz4SYS+gFCCjoIHuZknK8GVTxDlcq7Mz+z40Xet5kWAwhx2jD5+i4Nuv
PMzG17cz13fwHkyNIWPiZ3tzjtzqB5MbAMqdL8WWi3fZnHSKEc/yblN02fTqKhJO/sVM3pK3xFXS
R0iyoMmFTVA39+xo8SOGTVT9RhhSuXPjkXoZ+clysU5GJ6OjkMwZIoK4euAbqA/aAsQkvbVNz1NE
b0UJrfI5CzwLB1p8an9MVSKg14kJuOZXjiyzUQ0qMbK1AjQqtphMvCtFy268o2kksynUzsvvMD1N
fLuViIIL/DkZ0HQH2GQ0cUPoBTlnbsGlwX/gv/8y11aiKtftyLDQV+4bNBIe2jVrO5ttcLlMBnpH
TZZSJzVZaOUJ3epbSmcfK6hNS1Di8Q7u2YeUFHn2E8VvST55PwU4elGRv6ozQAMAtbs37k7qFEkH
NIccEmGyEH/uQ2zDQ+BTcNZCEG5bCAXGntAgKExdhsoi53teDccMKelo6dXlC5phky4JSOOTYWZx
832Gsk+e9oeOMWv1r2w4UYz9kq9ouKQ8kh+WabALTJfpTySCt157XIOA4w9Pb3pn8qhiLPJTMGNy
tGrUuB17GkPUGDW2XnV5t0Fotg7Gk0ZYv9bQsvOllQrTx4nBIRda9kg1fKonwGqVGX1z8Mh63uGu
WgZrfOcfLixT67vSKzA+w/e5l2amfV9DBKurZrjFcrviXgd3k9Uk+JkZjFXdNYs404J3lolacBuB
KzgikgF+3g5MvwLzRwZErDMPjwtBFh+vbP1o3SQcchFlEFUufB9um1xzUit0hGREkaYccpHNOqaG
hfZQClvC69Xe8K2HUdzLpR+gaV9y2Xfc/gbEbbEJval6qcrTdfvq2HCsBv8xP5C68RWWRhyZnu8N
ShxYfCve0eeYFJAH5vNsu0H9Ewx+rAZbmc56Pjp/5n0Mw8+B4K4p3g0Jx3H6fckh7nkMFn6DhMVs
2Gp4TpZkdhD5U5INgnhD0bDCB8LHuf8UcVuZ/3cjHi3R1+F7NzezQvvDvnbgO7EN5eUY4D1XYNNO
tmdNda9c9yVWa+GtFBiIWPoxKYhWK8ADsKqMiJMBlKII9uF1evrrc7iCs5apW1HDIVpsGW7uRGL2
KlRg+2cAwTSMiahc1wDjwNCqYL+c7w0Da2pAzz9HzQqr70aI2oYeuRbGcZv6xeGB7SZ1S7VZ+bZS
41qOuNGT5AsbT4mCqO9ay+SOHxbU5qoDbsDq/HuJW6gTirCqyw56uzXW/DYi3Cz4R6QNeRkZXUwn
Rvn3jiFvUq96E3kK5+dURPWuO4RJJ8rvkZuckbT6Ofq9cyXHKVRd81IticnjeUUsfz+tHK0giym5
A39WjFOCLYprNBHXEva6lyUTaEtEMvXB93dRCwoYpRpU1KV9V3lVD4F6lU+KbFL+n/PzW3vcm4IY
YV75bn1xroddxJVoIFvsuryZiM+x9YRHel8N/lSbHClUtHa2zyPEHAwZOXdjsesdbvCRbQtRX+Oz
C4jgEox8Om9Qlj0IfVLCj4ajypWzIZITmNPNT5Vq7T8xld9O9mTXL9+Q+nhXH5GaLseGdL6qw8sr
EBa2bKo6FufFzSstzBAUThz/NoblSKYHE5Gk/rXZYOElDO9cAdH22EOqj7ggbXkPDylvp9OETZxw
F1ESmLH2SZ5Q8Yj3oJdH6c/DNEQ+1PQDYzNPd3TCYEJTQ1wV+VF4K8FoWqmiHZoR/WVA/8mCkppL
llXH6SVtL2YB7FROb4+gu6Ycc43auTiY+3PnGliDIZ7dTeUHs9AsYYpdjMb+3lgVv5yU+sEqpfDl
IPlYh0yQJsJz5xIDtux4rzT44X9HG7vcmvxShNRdumxfTggx2LLKmnqRlD68m/jn1XbU+xaqJ+E4
yu3FIAdiVnftcHhPz6d2tpPQl1JZXiniyHMXcAd7mnnk3euSwa6pyF9MHNU3wAv+lrXQD+UDo4M1
AXYWte/6Cuk0oGCcikqWQfOr4+grjEk2AMcCAMflAuC9ZEqoYVpZ+3kVCguyAUSQJqaMYLenc8s+
ttuFLKGx8rjD9oQsFLIYVjXvnZN3kewXjqSW2nM4FdPFc26Crjip7qiS0JEXbqDSMpzAms2ZSNej
Q3Fq5uAas4BSEax6C+8Nc528OqqXRPqjtbQpeAs07k91PniHCs8lReaMSTybSUozBAU8oLGzgVH3
VUixmFHNp5lYcsb7m5x6CSdL7fygHMnXrlrDPd8QQ9ELU+vyT6YfjlxQ0H9XzfGyKyo0L5kzlQAW
tjRv/Ip+ILATGzlIVC+5jUv1dZES9tE9AHEJ6gUqfATgdq3Yvhi9wjNsSKYmS4+xVjGqL16gjGeL
pvlADS1kl6VWBSr2xFn7a2f7vc3vfgtUy3HmBh+gyhY5Zf3M49fLdJekiMwJhvmSzwgn9+ZI6dmm
LMgjF+on4Clzis+lmMYr51P5DHhrnfXwpbmOUNqzarTxlFrT886lGqW7zM5+Gm1RLGUn4u/4pKzO
rtoAisHS7qdrC1dGPW86qtROSU6ImYNdYREVobXNdPoVAfV/Vp0EDDjiXCqBNN3ct2bpNkzFAndh
U+DV/PfTQ9jp+qloToWmLlx+psYW6+yldt/JaLmeFYJQLfLS8w1BPeZgOMrObemVjsY+sErnxq0l
dBU1G1CvPl7SvwRiuU2gN/YzgxsTUBmlp9e+Lg/CGb0kqwCBxPa0l8fcX/pd0uctI7uB5Lrr/4f9
so+4HuzGE+NWRA+eWHqQKT84zT2oWDgC9iTYQAlS9hzUUEcu99Wcs8o7y/mrZ+7hbmVo2AeAWcdK
D+SW+CfY8LZCW7IOGT/fZbB2EE/e2nHHAsuLg8UZyr04rrl6w3SQ0S93y9JLwVF+mK+FFJwyGJnB
YwNvQW1BAaFfNlFHldjbP+RMqewqW7dOJR7RABTAE0WETZeju3NfCBcaY4CvxM/m2lHSZ3kqx10T
XmrUhugwy6mDxZZK4TY80plVxlcduWlpaTwG7Zuy9+OJBZXD2ikOKE70eocSsOeIAkQ5zh7+i6W8
2kAY266pZvH/lE6jvxtQUjR5B9NApwXgW/ac1rhvVxIyQHlH2wuqfi5nLsEH8MM7emCSbeCzFigu
5yR6Qm/Muz+O2PahpJf46UtplxVtrcPYKXjw09FCf/vp9j9A56pmcKvObkD8+rcOAS52WhjNMMWI
SuEgJRML9VPE+6jJ/i8YA6DniWYdkrLF2PNTHI9CgfC233wJ+Ovu0U4SPhnpFFdAB/niw7ZPLUTP
wePBEERjs6a5XqxkXSG9AvaGXbwtvvfIg4C24PnL5QjyVvNckGLC1+nqayOwQ0FwZYXmKKJgtqFK
UIhICYgTBKMbsyIth9vQyrHKdFH3lhPfxH5lCTmszY4JFP6liagDqDqt9wguOFeiU11ZN6++mFc2
I0FmF8SQGcoxYW4A6AeiSLC8xWpIWWiKDAfEW/QF4NE5ZGqgQc6/6Z6rnzcsSkUbepRg7j6t5w3d
/1wvqOzgYADVcs6avh11mEmnx7MLNyYgkWEy2iJFN9gROFZ0jkpogfvnaXpybCLcs51zkvJilAFO
ADSD7m+TuRsVE4eCMb1/YKS3wyLcERuWXXksQ5iORzrlKK7ozdrYKizlljEsi4NxfpBjNCYHYn1e
VoCr/ciU7ThLQ/7nGMDXetcnIAmaeA6hTHjx72aTR4pzLi4t920dfc80OAhtWf6e9d+AwCdvnQlo
f2KhvX539iM88ql8iLp11JzFCrjnLlQuaigq2O6aaYd5wWJv0tbi8tguHsj52NlpvbWklYP2mayu
mVIPbiMCflI7McdlzwjVck+o6LT4xOIqjNr7i4BBLPInte8FALJRCrd6TD03UAH/cs97A/kidcYi
FjsjzWqWzWNhadOhSNcJgyG2a1y0YTGVVT1XQAfTL5JgEOaEuJ5HhoUPeXbk9VNSM5PkQ4JytoxI
yDwCsZF9cPsk0VgH0PlBiV9/vvKlVb5j6BLFkYUKM9RS7ipmba6CPAUraDRu1eouGYNFIgRtkXtB
MzTInLK+1ATPr8roDNvEKplFBr8HZOGdVzt6SeVQ5Ce8Y+/0o4Wr48OnL6RBEYUQpC2YTJIEgmfG
mM78PtBSWkAatMbWRxViqVyFCJ6RD+TS1LaYKYoFDoj4iclQ1GrzN2KDLaxMK7vwGvyCrDRoJ3BF
0v9hhJyjhnUTF2QttUPDSfTNhebLjTTHcRBZq+eI4vXwBtsu387UFGEriG4kFoBkoiPgzAhlMN1F
xV29UdZphTknPnCe2UYRF8JAc2HGX9oaCzrFS5rIBfv0Z6b+U/AEwUn3puztBWYsBlC8ezSKo+DP
2CutOGbTgE4m1Rlb232WXbkLN5M1+jaEQkz+UX/CJLwcrZyOIUKuQnh6aexbJ154VZuAyoeKxZ3T
RsMhJV43L291bYgCqVOXoBUTGgi2w/Eh0S/Nq07es+M36A+tVcwFmGzCXRFKhgpojCrGvYo/xvMt
w+KKfCJT3qzthbCTLp+qc0VSjLwBJfMP5JoAi1w2/EPjxD0wDATSaqOCrMxlbAmclqVDPd3X8/qO
zbZBjUeRG3E96H3i6Z4cYGEKhshDb6GWUl7H9bz2SAFrDR5KTHBzTPfdtA6M7SB57vicBLzFEGdf
NECLLh1a1w8aqZiMANkzejVLaC7xwE93MTvXWuxaQcCagCLmA/+cIZxrGgc9afDeaXgLxVNE2ufr
Eh9xVwrc+LdRYWk4bQ5tEr0GlYVMWlOF6j0Kb7wYOmjLsLBkq2rebW+mloj4MP71k0Wxkkjtkygw
kpstuSbE8k8LaokUhUYMsNVxZggRhUop+tUmLy23NKCO0V4JQSnihEoJ/owxJZawmjJ7QBrexmYJ
i8NdS/B+P2bFdMXYazHscJd2Sl6q3rg/NlBucgc+NPG2ptcN37IV5tnkTMtjmp7T8XdzOBHRZ0JO
Eldj4lcVBvGcrU2KTuFtP4Q4H2LVNxHeWgvG60zEQHVm0i/d8qCZFUjzHolnNOsLA+yYRdBTVMvW
idotxl4go97twzkK2ruWS7evc36sx+V7+NCYb6BRfE25OBz1kci2HGgolkTtgA6CCkoUQGEx05U6
nYC2v3tKinkQM4+sed+c0Kx7uaP/fMvhOr3pUl596Tc0Ob9dIiy7LIQbUFK54bTLJDswG5EOtd+f
f3G8UGLvT5SS1gauG+y3xQ5tfOcF2bQgJT3cPljTmVq+fIbxUNqGe5djz7KjF9sRVfxCpe3xLGJc
PHAqdh2JqeoHH9/sriMzs5GOI/C4KPt8iZASSpCuqYhxxglwfigwbxPI3TijrNcPYFLzCpvmOVBk
ouVzm6ALAh+fqhVt5IyVfBEK34UPIMWnDfgL5h6IA9y0N1d3DAsnvYzbOvH7KdiOpBhRLn0jcGMf
XqdlFtaYA6YM49DqbedeqVyh/fKwVLqw9wY2/rClSjm+6J/OAHgR0Oq22s7MHOMCaeEliSHGHVfA
jvNaH2JTv+JGhNIk6fECIyJ3ieBaAagK0hJ4chEGGV8mattlfxocKlED0cXWCWb4apzGZDX6bhPO
kzTjv67uplWeVuYd8jf/aUa5237sIw4Pp77sxjYHtsFEzRLV46vyffyILqnGdPHGOPML3DNxuE20
0XtbeP7jQ9JW0XiLGYvtpqsKhV2mREa7BeA8BqHdRAWJq1Gu7is2cOoMoVXfoCCnO7DfqICKxHB7
0b+J78Q9z5WUY+BCdp/62MoCt7JTDTMwf9/JdTL2ITNsMeX10RVQBrsmrOuo8ER1MW9a68wTFt2l
etBMmyCakzH96yNeSmCef/U0rydqxwNqbOrjnn19PtMybfyLCsz/gOi5KLasvET1Ni1GxXP6F76k
SOQz4NKthOkbB1KLEGCGbmWdyTYARf6udbuWBBcSwN1VQHFWnB5AZWjaRZ/G9HrSM2D+nOz33xFK
yWl2t2w/xRWV4b9TU1CFwJC1K/Aig6YsxLDDGT9w06RkKdKfviyG4fty/DJf9IocvKnBGeOb2gwO
uFTiHaUQ7f4RLejRk4Vw8mYAHXkrue8fePg56+xI7+6cRjSId+OPBgUxGsHey3+krbYVw2t6LPv8
drN2fYRggBnvsZejdDcgbk516mRAGP76wF/20WV79Ml3dx2llx1Si2E4YkMjJoQUEm0Ve/8TvZyQ
d5EM8nPb/3t2QN/I8h+DXS3ifNUbkWTJjb5iRxl730YZsEf3rPBJniOOOYe23wVPPaagN7RcNO9F
QfQ/U3v3TEuV6MBVVrkMNAP25cceBYFeV2zhGzEc/dvRm92ZnycIPeKNVRUTDgo3tk08JLrTj4nv
oaF0B/3/C0nDwXImAzlO36i5PxtZ81mB+ghdteXNjPIBRQmPBNv/NZ221mEE9AfOXQD+aoYAy5GT
AkEjLNfXv1eGhRCpiEAj1l9DCwPyikl3ypuxzlhFI+OKlSQa3R1wxZWnp71LmeHJT+Qf3lnNl8w9
lYnXopR+RGFrkwWE9EplX6r+ynSEoimIpOv14+Xpf7yWIij5y5yJ8hh/OL1ia7wpj0lQb12ehDZ6
VKPUWuojJm3F/TiJJgn5e3i/d/nO+AmufmKQULFTi8vWbdgz7yWN3DZ4di1UNGT2HmYAt+Eoja7N
JyM9gGFYbzL0ejcWpnAiP58Bxy/m9Xgs/YIF1g6pU87wYonopLUeFA3d6m4geym8BJfN0kxdxcUP
iUGzwv0rzDdRlk6PegtnNVELkxACydBvDXwOiwrAogACJ7t+m7lAmWnDw3xRCUiMpxt1EM3CDICL
3M2sGEGh97XYwSRAyTwxlM1F4Rsp+9dGxMtx1nSX7p5oj//yMOq3zQg1Okd96XEfYIkaw2CcQkzV
ogfSEcFBB9FG0WdsoDE1t2j4GDHCvwzk/kfHDnW45xBjQqG7pr5TUsbyBIpkssx5BpTiA3u/W+I1
g7zjsVJI5sZt8DvkkXTIIdLsSAueZDd+jCCwQGvX9XnAxX9SeNyh1r1/QL8yh1utq1Pb1FDX3jJo
U2zhMSZNUM8W3wXLyNhtrnDCf7yfHnskAXGiVOmZJFRkM+1c2Ca10gey45gpXY/WbK/BWy688xG3
T5qQWs/jISjVY28GlxOGlPYquUESpGxuupWp9GTd9QwuwY7I7orHsQn/EWBdnroQFsOmj9XieYOq
5e1ZXrA3UTHT2bUOJZhgL9qxC3lOMOCV28DjhDY/U5I5dvjpenQVV4GJ6SjIjkom4trx3MKZcn+o
yoxB3LktKO+Cag7xfDa13w6XLd3IvoP6hpSP2m271jX/G5Act7Jke/UHKEvrvcAQXk+RkccLRn5B
LVq0HoMiF4FSxQJA4fX6NIfEe0R8CLMvhR+rl69MvZuuWddkcLCibGgBF46ysrv/fRDz/d6k2Nv0
A2gQyWJ28riHVWMvB7rN0mb6ckX2T38zmemcCD3o9cPNi2RxHbzgart8acfdq+1drUFbO2hLsQJx
jEOKbkpBEEeOUj2jY3rz0x49TZZfojBba9KQDkzdxeqN3sGpFjdC4ZVc0xzD7CdLkIA8jGLpm3uq
uZOAwTjV8d1vtIXGE3H9qYIGYy/aef9+bI6OSRHQSPHKHVgVUYe40uVL6W2Ye4gD2YmJh7BBb+Xi
8B03Um+owmzV9tPdT6jBjw4HNDdFIQbIEZOd4hSDy0PWZmsRYb7lTv9xHSS7szHSUMLco8NC+w6y
+3b9zJ4O9fNHPixP1p/LfghOYTIPaNEqj+gcxRxgtmbSFAFdAJho36c5EUL4VZCsMtc55p5zYoPN
cjtGZBTeUxOZ4Hf3W4eT2edSbFHiSR+mQ0/mPhfFFoEyb64cvXP1h/mTcZD8goGOKNqbDt42+OFt
3ilnDPhPkSubbOs0vFDM8b8s6ClE2B34jLkslK7kFLOSLkskKoewCBm5cE3AXa4OUU8zu2qwEaBu
yukecjp7AYbDxUv9du28prZSJ+9uyb67h2EV7U8pPC5OfcIE7DIJQZn0ilM6rUWrhJTLWJOuayYh
7U5v+4prNTlLYpVuVNFrNqRWdgOufmrrCXDeBWL+2oHi5fBN2AIX+gYFm1V1rZGGr8tweNfqdDra
OGsOE4jdovo0oJLkKNes1x8WBP6ZsPU9oGDUvSaF2uIPkodlijt1ir/52Xe+OVf3Ur/ZAU2NVV7n
0VYNOIh7wzH9oiQwHFIAtZpZmFE2srnEBoBTj8ChipXyNvdhEo9/uGfsmz4PkZPFKMVTiohZ4Nir
JH64zeeYaTnI6XwpDkndr+A/U9Oswt/IPjdT4pGIxbDoqJNiz9Bl0F7xYiZ8jrgSg42UfR7EZU7V
h+scAbgv1m0NJYUWrS4lEbHIIMQJB/auElJ7zUQUutq1/XvpfXDeNWhdh9S/6qr81CCBrbZOOFdO
GxfR4ehJDEcB8i9E9MNFii75TZQ3eze3Ocd2bCA2F723r5vrJCyQWGUEryeTDxInv38nmSdW2NIq
kazOM7XgQ6LK0Am6Ny2VBMINkaiaIT47J+u05ZOENega0vKA7paYlabmgAvR6RFMCGegOBo7lzr+
q/8my5g6Jkd5i3AtH7PQ8UxyZ5aGjjJBTAOeQTc+7y6jJ4NAqZlASNlzq2R+g9lmakB1aB+xBAOc
c544FcO+V0CBXZ6MBRUfgPQlKLw64MfL9urr+VfujN506aV5TvfRE2tXT4cNQj6Vx2LmAThJ8jhs
sFvWNqP1Xs2xEezHsArj+hQ8CyDJlRAuzLrFmloTt4lEXWUkXVZZnUQx4pFPHZYFCaJLRMnrtgYr
4HZ/EewdOaaaSoUAKt1RGp+N82r2AiDD/+3uDGCKngzbtWKrWkhmCVUfMKydkT8+rbsd7hilBhzr
CPR6imXkw3lsFyMWZt01auUImxJR1MGxMcOF4XSq51EtqeYBjjqBYfU0dl5YHKYoUyaDcTDUwwhU
9TyPzHF0HK4R3AxFOThkHUiCvMPKUA21izzzZcagpy7LcXnSUFvNZwJTW0ojK4vWHT2rpMLLBeF7
dwLWBM1REfLykzozYk1JYjzRx+5gQt9rSULVa4pIDiEReMsqTiXhMsYIHygXl6UhMC4bLIV8KN6m
5owiCJJsnqjOklgH6w2fBc6VFNfmdbt3L1UO0pqRojHS3YO0GHaoCKwAW7JmpLWlOFgbhY1ERVsC
eWFICLfOMt+p5X3r0Xf0QKtTdPT9h3xOGHSDcnDXPYEpvG+7tVz/YG7iurFEs7BKzOSTd7pkGChK
Olq4/wDVly/bP0k1C1ZEjdIVDQk/VlL6IDbuuXQoA+4mS/Gvd8EXFY8Hb8t9VzETxhlzBxGEB+pc
B6hvp68hOSeA4qggqTS0Ppl8+irzRUUXkvV9bVZA36YKwrXtJy6Qoj63bfOPsAehS80TAqzjznx9
aEz0+qklTM4GYuMzuwHcq6Lekkej+Dg4vN3PYwT7uX1LaCrRp+wZpPv7ZlYqb+0I2dML1nHmzDim
MmcyeMW0+QyBrGiLDTvDv6BOTuC/+550yYC7E6zBKbloRcAjvraSw86i+g7pKesnKT6ermLCnPk5
Al8NnZoIxj/8tqCRbHRgSrS7KoKlmLYIFs/+xpjAveduN2HuwHEUdGmhW63IrTY9oSULUVjoF+IA
+iDw9LhMtBNrVAC7xJ4FxsWWk5pqoJMO3zpleic4x0KsKRO4TUuDy1xLFhpgLAGnTo/Jv6b6VORj
E8UpKm9OWkRFQdI3MFGXQ0uuQ41K+aTHtHAe0VLVcJnkq6Rbby0LsZy/Goc3JejTNxT1xIDTcqjM
l3yuaBJ7CebaMXQVFurs8GIRSTcpdVrj+g23BnV0zVUEvv6uGh2SZAmBdS9KVpIDezp4QGk+LvzK
sxLRCbWMFJVVcAeS2PAhcHxYRPGWBSJ3b72lmCMB8ff5i3bLARSFKiF52+gwqy2lz2ghVAxpmEoU
snr2UBGNB6Is5IJysnTxSAV7ieHNmBzK1d9wPHKfLYl3KmGGi9rpIDP/5MR1fnFh5/uqgtMfzkXP
L7ux9HF4Ur0rW/igNeESF8ctPFv2xsbu7/QtReU1b6Tv2cqKZv+9PtIq4ZjzEMqsH/BPsnOh6Y67
6I6HUpjDQE36kpwpiubYj7n56QXwY9wR0EWgIP8HE0OFtqtb2UCiCe9wgC5SJEQKtqnzqHAUJZxs
KYUqF+UoKCA3fAaw558ZFbQlQAVbEgFsEaU9klPsNFlJAOl+EQzzPZVGcj1Y3hbwkhgz7xYTQju4
zd7lZQOPP1BZtSUnmuBFSDb2Mklc3Ghwnl1HbAzXCxYCUrp5pIN1+HFEn8pHw0lCzF6RDVeoSAuh
UfN95Bbu7tToyWbH8bjVsqeD3TUW2/EcnSZ3g/uSQ7Yj9ml/VEu6Ivj91mrkF96a6ZxZMO5cowkW
d2+3Cjkm8CGcD+mmB1n/Fj4dlkhN67SNeUzmCDZ9Q2qSY0+nwkFtdHwQd9CFMJKdFpD/8yEVgDoK
V+9X+rqvODdblRxjLQZ7hyqhNQPmBRiklVSykknWK/hbceYeHQCnTaALrZ+F8e+LI1kHKl95K/dm
+5HX2YV7jP1C/hrQVALA0BIK8sYoUDK0GzegW9AH3b33I4JJfKJJW/aaDabwovp8wHtvf6bQ79WY
YhupIat9eV06skd0YwQyaY0LXbW9BZQAb/yfltMqK9mKRZgND+w6dWYqnYkFEG/xpgmAORIGiB7w
MGAESlNdWL/cdxB0zfF3REinQFHotAZ+Z6eJ2bI4XGeajQwU82UcBgNw00jAW2/QOukzCAlQKYKV
3U4BQgbiq1Akx+QhwRg8d2y0R6P2GiNi78nfduoNaZks4Fw+zhWqhujs4Vh3g1k/0htd///lIiX0
ci/71+d3If0sRfv9bIpzq0fF8gErz+AX+MhGl36EKOKaCiefMtgduDKgTHUKXy6hnv0hMOuvi86k
ZeBDhJ6ZPyYAXNfScRh7GLIwpxzk6M2l87RSGszHInGQh99C9jkDJm3Bns+zx8NoI+xKxyHYA+gV
+0TZClT3Vq/z+YWiCCDNlaHwhzGp6gqhKE558vVfZGeMNWC1PdTTm/pWd3a2DzHVx/MDm1pojn1M
9mH5lD/6A+JwijZj89BCCCHjFQq5rcNXLjF3aTTiF4g+o/agiuCBAUbiQhGjvQ7UVGiEH8lsIvBu
aAgWeJsYFkagGCxH02mjc/j0JTXwv0t71SmNKi0uIY5ukdMrRSKeZyl4rXElv6bu/xUt9qXQ3k5m
F5/kK3F2f9Mu3m7JVnQtL1Nsy22fE35x6cE6Vrp05xbXC921sMAinh5y7rz5jrFBpZVq90ZMtFyk
M/0bDIZPYwGQzYbZvf4esf5IAq/Y/t46y050UrqJUha/z1n61wtpiFX1LTfU5a+iQ+ceGO2Vrgvf
kd1igUJUpdz0KD1SdbcjBTK2QCQ5QV0duQLvrb2eBgXZdl49MTrADgcLbrxYQalpze6bzr6Iya7L
EOO4wLMSWJdG2TUrBDixaYnwdat5g/pRLZOIsSmPgkqZDWgUF9kzv2lmYyz2JRfHoLPpisrsvVy3
AngMdsjLDMBApMMUAgyxT1ZJA2YGhxlrJkQtnb63jnNroav+WMz3vqKO9KraGiKYE8ZVrg/I+Ne2
Do5B3J1MINDMVuThoKanGTqNagL2quzxJ7JdM/yvg/1nWZepHG7gxvxca862hscTSQhTxhBx2Rlv
AC0PpDoJURJ9LtjCZj+BEX1vj7zF4pOX6W6RMkM7mXQ1HJ2Z+KiZIpziKoNxqDpN6K66kOmSy35S
+2cRs9Gt6XeSm75RX6AxWNdq2ThnCQCkpf7dZJDAr4ck9ILtbJqdtlSA2Nk5XWlTU8PBJx4J9938
xPBdwI2q92aaOfpN0GrQlVkCGvd6uaJqbMrYRgxtxe0nb5srxf5YAyofYy1bYcAcc4YD7RaROdsz
bgjHaNy9ZMBSnMxeL17exuBuwSUHDZvCD3NlgX9opZmWzT2Axwadh+Jskhsi7KOLXRvZgpNup00l
i4D1FOjm7udetUC9mgy0vM1YXH/wGe2Qnf8FD7LEbTpeHLCFWDMrq1D/F1xxKnzPkQEbLTdr92m9
xBW/OhsVX6eVA5U5m76mhpqlLjynWYG83O4z2KA2/ypC+5yeNJLpckCGQ0RmZ5xHdNkILFivjo83
qBg0KLcq4DMABbpOy6yHuixVGlIHarYl3cEVWaS7vGsgYBSXdbmir1VxY/Jpyf+pPvfCqi/Zwzvk
YlzE4Tt3bOFjbjED0B8a1TAgeVIYVPO8908Qn2+7ud1tXfBnEcf06YwZ71wsW4fc2nbgokLvRHI1
IxcJ2JcCkq+5ksIM1zJwnpr0UOgPD7hLEo0nUfuL8IWiHHml26J4pk2uEI53Y2V/3w6ceXPlhTKK
014MHbZesoq5Kd4eYV5ZeR824OAFCpsDgk8piT2eYDSfSRTChR6fZgfpzhcx3tE3IiXiaO3zoWSA
aNDonN/HjLdw/1WlrT5t8+X/x9xgjMAUeZIjq8FlMAfTZV2GTIQRGuieNiV1Avj1iHbqnVDsIwDf
sYrTjDsdDDfLU76QBEdv/GC6nsmG6igCizAXgASf3eQ+BWtGMIUjG23FiqCV1I1mijIDh6Tt5KpF
Q8acE9yiEQ+MWX3OBw2OWnHqC15bdehMrZPBxFnTwaSLLGzC9GtWFKepbLqTWmztF/DPBB/PrLQB
bZYmx+x2TN/42Z7mzh0NG52CyPrb3iWxnBMdrW0TcP8KwmMTNF08vRas9BE1U3Z7LvMd+A/hMO8a
cFI0UaqvGaGPB+tOgDlrJiwZOHueiZLJ8NHc6cX6rfljc9BX4ATCPD0sPVbWKuxUEpkHTYxEh4hb
JDTPqP8G6g+kNKVV6hGauMQrQWmV9MYxanoRhlRO+4LffY3H56c1CeBh0rcnQfLlAbQ0UTrKkwNU
zrVg2yrANfDaK5DFHv6r/AJmQAQskmcfjgxKUJS97eyXDddZsT3WHahzWmP+4QnF3fFQcMyB/JoP
gBrBy00FK0eXBt9xNzNMuHLp6FYe23Ykogq+85ubOTSaPxea7QVPSZbUAHaMCeU0h7bCUQNAVsh/
Qu87npRMgR1TMSohkZvmupDVgjCO2gRpO35BV8N1oCs8f9oFlTTkT7jrGUvEzDtJ5OiM+dxeXVz6
PuXVWtmcs3jrl4GCJpELCZSYJHjunYZJ6mDs8SYh7Pv/E7LjWnbjJfgqoXMILrffdX9TnOy2FtQT
RZHueVYedww6Yr94QFIskpJSXZIEe0kqroXkTnzOhQRcyTOZzsE2z9VV4BgMO1l4LUyFBDtY8z4w
XPN/hY+pZK4pnhmtrbZdMACrvel6FiICGQQeasTI5o1MekPIulH68sbYI4QSacFCXHGmHrkTqdIg
7HiApkgs4CkY6Bb86qO31vlYuVM0+HQzZdA8vpigKzCVRdtTxlVia/SQq85zVkfer1nFyP78UdhD
3AZH2AcC7DnQ3ZMcDgsSdZK6QXsNfKHx9l9Cey+9RYn64szst4JVhZxhodNRiHJ5sYccIe8gggOU
hJ4uRCa1Xmz6uwO5tZPNiB1miBBL25GpjCaUT/pv4433YdP3mTaC1LpMVouOHE0kCSEKe9dr6UKl
dJ1GQ5h0jhiGFCW4KoU3I75/p/webh0L3uAsGCLgOm72fcyBriXviBkWiDQeDz86U+6KGFP2k3cx
zp3gOs+L1tTlo4cSdurM8Meshtep5jxO1cf9zjdgO5N0teBUuIhCCx/2n2eQj5YIkN25iAth1lW3
P62lOo+Gl/SxlDZekf9Nnmq/DekSMEedJCcKViMjvL8XNL5KP0yZz3QsP2H/kzHxDh9FQ1W0vnGU
PaOunFi1sAW1h7IGGpsrV9xbfT+rvudEmXWm155+mwdQG5uzNCcy2vHdbVtN5OVbcOAnCxdqDWuI
MuMCtUhD41ZHcXVuOX5h+e5OZ+zcSGP8978ienJpoxhoJVi/B0HwlqpYgdrKmVn2elDloGDj73q5
SarNRI2FEbRYja1blMcN07FCUAUDnsCImc+L2OQbakvNUIcZULe1geViZ9I3JryrEsV3Eto+fxKf
76frGG0Or+9Ah/8RwqIgwqluYsn/I6XggPGZdiWxi5M+ZkxSJS0+ePw4zaCDoWWjFO2YphtB4EI+
B2Y4TlQz2fr3A0xBUZRKvSCidT1C2Z61E5IB9l2fk0MnBqF417gtUeN7KiPLuGqf3c4L+EDgAQSP
Ia4II85DrtMDzc91bmjxbDmsR8FXEZCupzUyZj5WW9Tai9uF4SpwCO/n7TUyVuko4+q4R0qAaJ6t
xRx4ALFUGIa5LsEwwGWv8+E594KU/GzLN/d1S2TKYOA9NExQNpSAh1o3Z6OrHqVvDu5EhZMB4EpU
1mEUJy+CcECHg4KBQLFrMUrBx105QS6ejxyNYvbcV3cMop8OTAzccxhgwnjdFRh8TzSQot00A9Zj
6SCUX3FhhUgKluS7bqUWRtPg1K+yvoiQH3RIrN4YlPnz74d0M2r9At8DgPbcJsYlkbO5VjUQdmVu
EerXKQrwqglAnL/P9Zkqdq2o7JaOZ8e7EgShGZ7HQuTRYkqZA9vCEPN7MW/GeA8Ft/TyAg0m44XB
jr7Xps0uqhYewEzSgjyhS9vOQITbZzqqyJcdsWgFxkmSOADUg4vh2fs5ZDnyickZUlF678Hqwv8S
0NliwByYCaHMN3gKAhYHcVJ3+bU2FsWzNp9/t/zao2IMHOLjCCaihFbcj72KflDPZr6aSgIZph9T
GbZsBzRQdPXMv1P+s5mW/9jXyHdBGY6qGcrPCNwwTJPtCG0B4/GZt6+1jkTo3UMu+vzmI6hjwyaZ
HlIeNTF6q+/dt5SEYmthj6y5jdnW8Z2auogk37pUewNrfit+9jXLXVUEnhoRAI0FiEwaZmuXTc6I
aBY3wb6b+DPyCg+vzPPyRRurROYAQlaoE669c9wOv2V7QdbM/yyhjtcT1gZ8UczorgSWGXCW28Nd
w5lPlvEUE1cod+3VwqP9zezXb16jsovTQ4g1tp5Vo+tq1ynNfY2CqKzJ0r+dOpSB+gV6rIHA/H57
crGcQoSvjhEM2oTzVnEoKaPMbiMHTfZ1/eYgiBr24DhrCmRSXLBg3IHXdeVvJbrwrAONc40EJd2m
vAIN1wrToeEwGxwsAq8l53Y47n2ELTMUQDJqteiE9rcFOpoOvq1rt4r1ExLaZUKBh2I/Sqlerk9Z
o5Z0P1CtKkRxrBtiJBF0tr2Iec3+petmhyi0FEM+hThZ3/EphTH+Gj+XR+vPlhR9hO51jTvk8MIu
uvTdymOKY/+2yaQb/LGMURdFhxZ5BKoVH/S3D546whp3pYxvevNM0sQmFBYzdbeoDmGrzqWa6QEX
b/Rp0sLnKD9meWPQUexZ3192hM7McLJow2p76Z8sJqbfxMTCcmy/OcoOjxqDpg5W1Pzw2cBwYrUL
7GZ3tiRLW/xpniQvMSP8GGKTWrnMqOftLWzUMJ+WrbJZ301eLMUYItmTj5ksGwbh535FaIz/x4jV
fCPcOiToYRkKdA8qrQazV80R5iZp0r/E6OM/lLO9wKAGsXORk5VThh+Zhz3InIcliNqK4+J/vR8O
9RTKWnPApwIOToGE/iLOWPuGLVhoGW2cIn1YZ/4AnDe7M50tWpCOslQhaa+qf+gmmrUnuzl6eLFa
lOPF9Qc/vn4pnBtEqsXTjT9OBowbIbgfiaFJbgPo/qPbkQWzWUN3tUaGf3WRfRGThjYD5d5yDbsR
42DmLaYERUlDYD2VvljFDUlSGXupYFL1od0a7geK5gUDdRwRwOgKCu5SqMx9r1VokExNkFp7dsrM
Kn74CWawftGeYeBQKdMV9MXHRg/+RAytWrOKAVFTX7AdvfirzeWZ8/UMLXka6P09yJBGBnM6iFGr
LX1fh5AtXXzpqWswFRFTjjquKlTuHr91M8f3lymokPnNw2LOBW2Ksdx8Fp2t25xybUpq0/W2A+AC
0UiD3koP9jkbgrDn57wlfmIq3Yawj2KotxMq2Ndxp0RilFx0rF0/AwIB606n0KsDE+54Nyc4f6iZ
MHrORmmIRVad8YcNYnzcc6HZWbnAv7RwNIZbRvUABuIhN70BQLqWVjAxzF77AEXSDnMfIciWoA86
VPWUMWEPLU3hyRlblT4XpOdJ2WZgv8gifb+7OowAYIy7welHxseEfEphBZb0ba109XhrchXRxixy
iOnRYqV2116CqXlxhhBDmxE+CT8FhR9BBi3QdbAPoO8nLLrOeFH9MtU/Gw7juhSsGNWnqKob9Uwn
tvqSKLEgxLvndFXyHfG6+aec7sOq41LIT9OMxqj0+Tn6RZ9I5Vuw/AiUQy9HkY48AhnXj1eTfTiu
oQzjhTIKibJveRz88FI8/17ncL/9/w1m1n5p4XhCkXaTiO4yNxbvcPtHa2vUIyCnEzDaIgK9Bnzm
uR9Su2pjirajZL6U/SgOPVFIYRlybofiLskgcKQ8WpuTeLDHXczo84+B9klSVr9BsNDBUrACWa0Z
rjUi0ySisWrdUPUWoC9wSF/idyYlruv6E7qM34BHaUJSNZjxCJj5G7JuV9hlPIy/YbqxWp7ZArpF
+3U6BgyMtRaE2u2mTKxGDvHPtNRBQqk0ZOeHaxrFZps0+/Sy3iUOcgWfWyvAJxPFBamwLn7Ce4EO
txihX8TlddasgbW4yDQgxbNs0Y3R6uNywtvNDRjUJaBKOfdGUS3Wg9/c8aJlUj78pGzqFlxVQg9q
DovN6NXbpHkDdBDsaEHFpUMeJ2tGXqLfad9b6vjdKBNAaVGRNsWAmW/PGWBPlEjRGXjntLPhjPMO
LRtcQ0BGUofIR1hGcSrhrK8egtzhRCgRtpidIs4mZRFeYaCIBQrcZWzwB7KrktleNj6OdNY7zUvs
+LmCEg/MYWIQVEe6vWwGN7REG3gF4YnHHnyX2IlKn+RWp0KeezLBeKo7lNE5QwlHvPBePDFQxFtC
bsAUlJDSg07RDbhC286ufWdUvqfGpqh8Lwd7Bkg6lAJcJFq3Hjz2NT0Iji3Hp0N2JwCmK+T2D0Sw
UJ3+S0TsFc6Rx/O0pw+noj5bmJ6VKhUc1rRSRsvXL+9EjgAgFURFBtRg3inq/GLCPpKuuTgPoo9p
xjv49uiSqpyDOKFj//yz/NvZZXfKELAZZic4vEvH/m4FYcUp7lg6yCzHiXBJ1B0g/cCOIxpfNF9b
Cig7rVMuNhju5LOVc6Y3qyI7gjS3dvEYSJkLWQNS5tcVorj2TcXwRcs9XLhXcZSKc/f7om5PfJJ6
gsYlmIpkErPuQ04QAO2MkU921kZct1S9jNzEbFV6mMJbo+aWaEptPAYX/KxRrzgqzCMq6AT3yatk
6MKRIUEpPsg+Hdgdr9L9yhTBd91Wpth05AZvjLSkaoGzyn/ieROWaI95zb+/YRInIWYvJ+BZVLuW
PqCny1jVwnvozEByhkrg2fQf+g9xpRGkdjwgovDs9E7BxMdkc2Tz9swnKtQNV96o2JQoMayy6OgR
l8s0ntUOmEEcHWeO7uQPjjms7BVTb/dyNMeHFo0HXZDMoIMp3k6vCf2yHyH88dJADgeV4ezCE1ya
IVFaaeFDAi9ulQ1r3fE25B2EKojO+7GESWE0jk5dlbOINXRCeSEVrEC3Ki9rta3+ORSfYwBis7dh
Kp8E7WqtVGsKSfQE+jORpbYaiYL9VD0rvsRI08T6yPW+92MDVJZ097AE5m7QkxKDQdDT6UueMXC5
BRrqL9giM/6QiiuMv1tLTOEqESNvbv3ItA5P/CcrfiXGfw/RgPFn8g6yJ0WEQoyQkEULeKcur3CK
fyw7+zT96Arn6tX3EDhaWaPGkUu1v9a0k7ofH64bin594S2dPHOisqJ/1B7YpbkIudJM98/pxx0R
4cY/Q6FfIgZU79wS3E/Sh3CnZ7XysvPZPBBBfkcFptU4qZlIJfpStk3+GOjDDMtmIE4XiHFHivDT
r+0+YJ95FBI3eMSxWV+Nhr43+A1JC2eHKJpy4WGm7wGvsnXo4LOc6KNvoSn/5hu6z2QGPSgF9zgA
V4MSINL7+NZDZi8AbfQuvj9oCMVkQpV/5iH63CK+EOYEcJtbpY+/XkvKzXnk98Ll8Td7l0K0Ky/1
Pl2YBn8j3oE8P962Bliqmn3F9fg23lKWEpfyQuF6A4liu3RRazr8XvxwqTmYjobbzI00v1DIN8d4
ETP+4r7xpwqQ0G6U5RX6Qh50HC3VGlOhndl8CIDECQWcKQZq43DVctnIp5kAOJ00og7btESUdSri
s2QVU92HrxHxi/ilSoWhlmdkkIxHRpB6fEM9WMpZBWg6nERSembn2jFUfHO+Y9E5drZa/kKUzRXQ
NKlatyzGLZ0IUPO+IGdTsQJKcmP4paeSAdGv+8OcrpUtyK5EQzVA6wIVRmr7g9a+cLEiAGE3iF5V
+SXvx79NG/7VjFUIsyhkQ5ClUZ8Wkv34JqwnmnpTfJgdLPIggJQkddHTQFSZjvbHVXwtyZt9yJul
b45TUGCIeapdIr78b2g/EFTGEk/YlWiUDkCKfqHZX1/Zn96O3ZhYLd5jHcK0Jpln7s7isGANJsrZ
jgXoaTPY5tkq+ntAtS0I/iY5kAd0zb5BY+zhFqEoKt5XFMx1t9Xq1stAGwmb2/55RpH8szQaXdNE
wajA9RYiQNZ5KCnQQ2BdEAK00QTgwXNzOtvGtlJObAVxu1YNEpG3dsJnuQ4YUCi/g9Zh4opnLvUT
SvLWnLl9FGzYU8nMvNAgdILmKt4gEEQ1EFoXy7sZmddwpBYgZ5ikrnatnp4/4ZYmc8jv6D4P9D2n
wml51bNnNjAWclDLOM3orQ8oOBC87cQH4PMDTErk11Jy29PwvTVaal4qM8qjJVhLZHI6BrnxaXA8
t8nKsuHLh/H0ZVl4/B6fkx3lUTtCE5/gpA+TtEi+qG9qjKfRBbFI+JsJl26i3SPO3vZXQCYWOtNv
WiE/IO/l76JYsPQtleSOLUaMEuugMHnieucfQXmJoPED+IZ7/H23HM5S1hbjHD/5rS5yWyhyHoDE
9fyfVkd4Ym0Qdje6yjVxhzaTfq9GfTTFbZi7XBsLEdtZ+AxUeU8O+RbJH/+YHRLN+zTIQBfJ6hqb
PdHAFGKf5oZ67nY//nloT/lTYVPeoFED1An4F9CBAwjrnEzJwgfygfwj9YSYeTfVMZ/3byrcBsHa
dnha+LkaAICtV0TEhX0AjPupXZuFPq8d7tDw0z68D2/h4L1nD4B0YwkSpEc5sSUA6vn5N7wEftQD
w6dNFjavqk5DjGEk0ku+TAY4cqeaRkDnmRpljrhgLARcOd3stDYMPzc2abgRpKqUtbU30dH+9bFf
MfEO4D+XEx6A2DFKDsNYM8QSlzk6ECacM8oMWbL4uRJywfr/MeVRIato6ntqVEyOdCWqGioAXYvK
fqT0iY9Ok3eggkZY3pXr/6bhYwkcbGl9XRwh2Ssohjiu42dej2hA1/Ok9BH+GybKVoOF/mIMBHe+
mO5LaTu6TvGXqMHGydTwUao+OIbwbZLMSBCwHLcPTZLFDaKdAyPkexzL+6U0a9Tr+ILesgjLudSG
/wWU72aWWnjNWgMaUmsASgaqx/O8sdAWoDsmxvcexN2+YOSn6Gx9wej6M92HssRV3L8YSxs6mA56
laKL7LheU5y0zBvXf+pYv5emPaWOYBGrlYlS+b6by+U94tbwhiaKKcken0trsKkvDUUsOKKEozZO
3eiRAb4IiSRalfBFZjnSph/212UWupOzFL9EESc04yqUvFSJvTgRQYUsFVyLVLBpI62zPQ8JmnGf
sv6CCzZu7MePFAw/F0Xx8toejPSpi1/q7XEUs45PmvIUsv7ZGQ6wsdl6fgDWrPOKodVPxKsMofGJ
qwFrky1zukGe9KTruc/A4wcXmQ49eTpu9hlJm1bwnjJThnFIQvWOBcq52XU/Usz9kZmzPW5UrHCC
jy/RgYErNKvWftSni/7Mu4kpoaIPRsJl/7OViVZTHrS8C2tinEC6l2PyCSZ/t1RAsFX8wOMOEil2
Rt1lawot0QHXjLIc6/azjRFseKqNB+pKF1pD/djm+LCXMCbH/0ZG+hGGlM4AQcdNW++316dutk/G
ZwKWZg0CiTk8aFIcCm7YoWjAUnBWF3qX5g1uAB9fI/cac8ks/Hapd9thodLpJc4rOE97By9K5qG2
u23VyY4etFbBznSBXW4p3rGUl3aPClvjkyteiDCzr0kMA5UZUh0AC6qP0zc/Gm5eon4uEIKBKgsL
S92klw+bHeID5a29HCv5TBYm5NeCz+MmoDFggySNg0idlqJYbmtE53r1Ig4stTntDrfz0nJ7QTCf
VG9+02IBRRXPo/NkI4y8P+ompXLcQl4XzTPfmBBeX8GV6bsGObR/w2KniED4wo/reJFQyVgFlrnk
CFmht9UXfa9WZQOlHOj6P4a5Fs1n0eF/MrHJcL63exWhK03Bkd5Oub6rpkyqJ36Zdck9PmNu3ImO
lfZePNlLmduqUjq6BxWtKMH/B+sRBBAdZWYeKNH8UJMdmmB24dkZQTNz4T+fdJYUHXmA6EHUHCqG
wZbO9P2pDYhbHtOT/Za+g0ejOzNZ1RKwcFds66xKpHGkrLkt6OpbGh8xsSKl66hol1qncxoCIdWe
L7t1MS0fkDUq9+ZtnNZOfPUJlbQspU8zJusCdSyUSfUHYVx0FlloZMx0ZLYBx4htffeSfFZQQiam
HAHLOkOrGW/ARgm8qL7+NKfPMsqrmRn1A21qEV60mC9uBJYEvUx4EO6PGcuyHfejjMW2CyDzZUjR
zSFjCyCjtH/NcJVZdez6eh4aSnZ5LbYT7gVnonBfpUxW+ITMHU8gU60WAfH125E20XDSMhT8orTE
aRJSmSUTpvLS3EkzFC+hrnW8JCGBtLorIg2B4fVAw0HbTjjTGHwyI1S2vZ5+20U1wOLTRK7AY4jK
rZUd3Hju+q7kKCkRPczMC3SZpqszptDAfGmuTYJMT7hyQes4cz1tpULddekUIfmOmW5oymqz/9Di
nmC2/dEnG5reSjwlbEtV431IOTweXa3aLxrz91Dw4Vh4BBUiNVLk1YlL4+srnvTQLEbg0V8dlVVz
B3uR+2HPWXXXRDGQTaSR0DbuJKeZVwcq4qC0l2BQ41OMe1o+vCDXwelvIfKIT8SejEW+ObgvBKZk
5mU1sF0vj8KtIV3Tdxenvy0p2TP3Of5UtjpzIJI7668cYfthlCATq07gMLvv4ZfYlb36LR79bYL2
A4RQOWPWBYmlSCyuiKUxxn9jGTBCyFbePYev5c9Uz0GWhANkpd8iB0cqonu7wmBVk6vk2UFaKlGb
O1Zp1tiWyqfJvce2mevvkphxyWWYl5TKwil/xOBc3bECU4D/zqvHkuBKX+tCt6rEHgjpfdYkmNoY
2U/EepmSvm+lTjkdDz/g8SZH0BSV01ZOJ7M/he3cWJibVAK+HKd6SYRv4mvd9s+u5g+eFaRmnv4y
iJy9XIcE/O5fGVl7gD5EHRidvpfGQ5Hx5Fko/9djFVLZS0jycwiqUsx7MFaPCePBSQTWRAqHdqCI
Dl+zbgnlOdVlZyJia/lWyIGgMYL9kRhvhol2yJaObbDk/U0Qb2txTzLWcZzkXyy9UZ4zZ+eWPFDC
TsOddLD1nP69vmBZOg3xUryH1mTGTvVEc3Y6rgl1cTwvacbctoibouf/4VbzjWyfL/a5MFfnkZTw
2HicfD5l0lD6uBe2+QkLoiJWPzwYAdlzettTnzCsKFFXKZ1mvkSk6TizaRrGQHi3QaezGvJreN0K
bWDrCwGp7V2TkN5j2fry9e3v15dgzyW/a3WgIyyEvTG5tp6kQSjSHA5RDmHP7OIstYyRLkDc78vw
/m3jbBL9htPCx1YSFyfyPpJaCkm+ba3L9yXYpO8DeKyPWpqoaQN4fKCTkY6jKZpYiizIbdP0LmpR
ijPA6hITsXAmXp6OVkqsWuz+9Yn9qpEWWY9qPQXbZWDyXe7pE4gUEJcug4kkN9WBtDwqDDz+LCCy
38E6gG9HQgjaNsUqAlmXExDIlQ7Rp4NEYbx4hr90nXTL8UeGa4BRuUc8uZSwABg2BYonMSqxWosz
YL9gEmFiFNhrRWYy5p9YCz9InIjGFF33/dp74RoXCbdlTkG30PnMA8X0oAZPFCpU0iHNdmWDUOeN
AtB7vmMwStbej1t2JalPgPY+u1Z7J+MoAhVlQwY3am0wv76jREcGXwLDNEVqa04qK14MUM1gXb/N
eLrH7CtuHIONiaw2O9IA/yfZZD4RQYm28CbLeaY7N0IJEbrUG4FNoYytu80A76Kw1PUdDyUURVxx
h2ZJZ6k0d8GNA57WXUQYEc8EX2StuYYm84J2SNm76y8jEjAG6pM6EZyihFgQGI4U8mWYFTuj6ULs
cOM3cHgd6NlsIEidhAmuYXpM1BRVjHZmVUv9kr5HNWEpC8eLH1zWRGwEzzdylBgIv1mlq+28tii7
rVaiQoexbMTWIFcRqQWEAq/B4KI8xR5rhWKMj613g3d8qK+ffqbe2BeNkTuQnlVlgJSYrCY6PkoW
1/D+ekoCilw0jHQio25Qr9ojgsyUB1ypl30YjHd5dQiyxsCiAwzHc7Vs49TUinN9cTVJq1MgFW3C
RikKF2U3tcJPE9XawqJSSAtc84P8YR+J4JPpLjuienhK2cMFnodUnCloqV/LGy8vWZOVb9qSE9aJ
bfF5kRTcoOyDkVNfcUg+rLL5dkpkYaAXD79Y7DCq1xDyzkx27Wh7lo/fu6tojVnTKV/02HyXqhaU
O1Yg4hW0XCTX9VX1Xl4jtxQWaLQIZ5Gm4sUioziY+L0/UleS4293tEAklD1MA6oPWxwxrgxICcKX
j7Aav3YHGx/uLF73HDnjclkWKfTtns2fi7BprHuezROt8q8w5TdeYbhpSoWa44RzyQh8kPL1xLEd
4QiTGN9QUMF/IVgvjoHQNosv0yehC77OQ9O/Ic3D1O7dvB8Pl/gnTtHvJCoth0AIuXwQrcsk9qdl
dxcz9TBg9cnDtkIMDXz+YYgZpZpp7fIU6OILeWdF7l0/xj4ZtUGyD9bqSa6uLNGW4dCwluaRV5tU
SP6lZUUfC5iSFgwlICN7Mmin0JhZtf/V1AO34jop7p5lpdlbyWHe2U08EA283H2Ir8FMPMbrZ42i
rA2HgO42DyQe5NsHEfDDsS3o5s5Bye+qal84Z7b/v+8OzhMq+TgfB1Rs5UHC7BGkwlxXEFOpAmhn
K2RhZT7s0BmwHtUIHmAm8wv1ytdor4CRYaElRpKOoNs6PyOqgIeTW/m7FrOw7qrKmaq6YQD0AWa9
3whbW/mQI1isGBa9nzZnHgj5x3kYcOI5nr8MFXrILSSoOjRz4g2IpZTRRzTKjfameIcsArngQcaD
Rh02rLosDagWnnNlz6XDnBHvZoTgVXkoK2c0Usvl/GK5jP/n6tqBtVUVYojfodIz94PFeJS0PaN4
fLnoU6+SVaziRh23sTjcg+4xs8rbubompe7xpt+Bgn/RWvUZoFgQYAXmYudOTJKk61gMOWWoK4rN
pm/TWCgu+uIzcgyeruze+8wTFoKVpuW3eoboYllrxVcjSQwFdo/SEBfgjZrFU+SgsHV2dfqTBWJ0
AVUC+VTNt5/wdUgo7dy3oS8dnCXnx7IYBoXPm/ihLhPy5rvI7dDN3KoSp8/FHdh9TCsV4YYWVJZj
6Dq+2GGsO+Nem0lZG/Vhey6Ynt0tmm46EsPPPZ/rcTj0sbk4vKLKHaZWdR9zZf6CWEpitkvhMElV
tdK6vDEsU8AapUE1TiSz9ntCo/KMlfm7Nyrojft6I/m7HqjxDzkudxQxNz/Xt55tYk1346mtXwtZ
GGCoU8F8aAPqguvpQFTqSguL4F7ph0kdi1cyjQUJkY+Kmy+XyYpcsvel4HXb0RmNeBWv9UoMFuGo
8nNTDvvR27CwOXEsPIRL5RJeZCUuBSIz21+2o0glFN7p+mMQ/U9M/woP/Ma9vJT2zw5RWXvCYVS/
F89TznUXc4TZdUHjqdNI6N96dt3Ar8niDuuHAS+fKfCY9tEoCTMFByOT61n8vq1m9UH9epPKK75K
ppeB8TOklVicDe6p/SNH2cekINi8E15bv/eVTEyyOdjE1W32aPL89AT6UdaciMW6T3rJoUXXN7Es
dZITffG10HPwa4FYyqigbAxW+IP/oxJknirB+Dt3x9mf74/rCngkdRnIB8iZfrIt3dEjuauOxxB0
BRJpVdLZ7n/rVYx79jdL/QipltjROtKek4V2oLCAsioULJSlBHRfocNnrrHiX4NTlScA795LVFd4
ibquXeKqYLTfqsUaaJ73gAAYerWkQLGvjeP7MHdZX7iHkM9EmlyZv3pmm8BYoDPDa4yHwix69wH/
IlDrkmgd2i+RL1r13gjZn2A4soyFe60lAGlVz0RgVSnPlcBvfyJLjDQiMYAU3inAd8Cf6V/dXyQ5
O0an+sbqiJde766lGFVf4mOPDjqFgT402YHdAZDHIzeEIXV7Gf66PYC7YlFEwbH1aFm5A3UYhWl8
oEvx9f3qoLc6j1jCVnZoXRA6+DR8ERzQDoVhVB0cSZ6/Zc1ptG7YfM8GZ1h9I0hWyRG8LmuhEmE1
UQ311iuF1NYE/6WFsQiJBscvtsr54EopxfUAeKPsGWeJaTvDHJsHOsoRZZ6EFb7gnlaTZaVwwvWz
DCwwDhotb8yIkAOnMic2OXoTvMOnpuXTZuL944DTJ+OecdolKEQoU6D1tt1gDxW1zpTd/tq2DloJ
ix4t9VrY+inQ8rZhq00ZcXyIqC71qaXdZ5Fy7XPv0Ank3DZVeY6LyXKa/yKPOx9k4oIffyiR2tBz
d6+aKI4vK6ueerE7a77U7bPn2rEy6ZTOBMKuKjj9Z8waXy0/DbFctsHulFA4adoxE69jQ6xf02vu
nirG5i5H+WQKEzWxupmPszSDoI3d0iLXTXP+030PseJitfpSdJn5FZeGbiLE54TlZ9TT0myLqY4H
pdQAHxEbFWcx7++xynrllG0KFgHEDjkM6wJNnm4v+kHz9TJ0zVVkB+48LIwhwSAuEHjl67ckUb+Q
4de8R6HLVoEG0dohzZ+3eqi9ZOcj/PNy2nSw43+o1EONMtsTU3cMRoinUgnYnm1lg86TgxadzCzT
dCaxge1vSWH+xmadhVP098+cazeGbiTjFJ7WnTppoSBixxYV7kH3XqkJ1MsLSxpxjBCojnS11iQB
BhngAhO//lKSGFqIPxsGIj7965G1Ck980evfFVTmHMksOuOic7GHFLwpxMLI9wT2SDJVvJJakAXE
Abap+7eRBwXG0MUnI1Otkk5kP8qn46qUnurdEpkXCUMZZbUg2snnEZF6EqaVPT/lnwGnLU9Y0TQ5
GIW1+xWWrOT+oi7ai7U4Q49cOwWsXJceD6FKpc21rRA0EJahhrv8oRZlBBP99ehgw4r1OhpfdTij
4KgPtjSOye9k5PG1pLIxeRriv9rbPfQPBXbIg+1bnIBEkwkRbeTsWNpcmvIwyo1Vfv5pgv1SNJ1W
8o1coFtXbyYBJ09eKtf/8sJBQQIfKCvyC9st/mZ2YgpwqAmp9mgV+NEZ3RD4Ljd0iHRe8sxoH8ct
f36M+wXNdPHVw+SFPw3W9nsmTVbNS4Z05v16sVMecxHT7AY7Ond1ZbZqehsM6ev229wwwDNLtXR3
yjQAwTHUVvuYyAskoJK2Tn2YJJYM9+NsZgb8YQpKBV18QbT8yvIrp9p/54C4MZUIUC654R9jpeER
pD6EReeVFZP0zwmmAt3F+JyShqw6ahpUx9A1ASacmdbzkVYO9x4PLyKJ4Qs4xyKi5604R6+Av2k2
VROpbXP/ClEGTgf+1oZpcmeeE7Sl8eSrLXnIv7wA/icaljLfSHzYQ+icuLNkFGe91HM7x/Ge6ua2
KDo78xMNJ1aiCAhYRTw2PO3oAPmd0smYc8W1DUdyXvkgsjAq1byiTejuqSrZkprSq8/01g6jv1zO
EG3AuAJEl0ysvputlaQtLpunXPypMC5RrCXcCO5w0d5iOAY/v4YgA5x1A9YADDT2U8tDiJk1KWQP
uzVWQ4c1siZZ79K0xCeVk/55/k3db1NKr1ooMxBIRa8CJ+5VJTaxZkhE2RbUpqlYJR6srSt3S/CM
kI8nQEjKtBOJ9sQxZ/qMmgaNdKWvHL8NsHSquvH35lOvbTBsrucjOZ8iKABvCqOO4z3VHVY3GE2y
KE7xD+mZJtxzqEoY9K9URbiNIV5ZXlxrJeVMLCyGB7oHPnx4dA2j5BPnbIiFyyz+kcSHiazQ+w4y
gOgRqugwAKebpdU4Z7QhYCJv/MYWCjgCYJL5FUt7zC2zXNYBu3r/HmTCK9YLFCodV8UuopKZ2t4c
iZO+h9g1W+ktQmco/gzAeMhQJcBOSzJRD1SZ8WxAus95uONwAJG3x4hvZ+11V0Fi4gp2FxvBsl1N
XmXs9OYvP7i+5952FnO0r21nrCQtXBewL9W1ta0KEA+9Arml+FfyLGAZdwG7GM4biD+kjf2qlc/I
nJEi5mRZdPo5Gtrae+X4E7oUWKDzItiEI6b1LRANaIKXrcPEJC92PFPSpd0Ark9Up6G8C9l2w6P1
tYisjsc9iG0slxhkZZw4QSbY94/N1HNrms4MzdHgeNJe+Ks2wTh9DbHSnqmwctkkvRVmheWwVBj7
zw7ls5/UXsU1vrhvoM0oxg73qBODX7ttIlaw9TPFrNf9WPtl8PWK2UJSxTR/lv0B9o2YeQHt4l3W
rfqx9EsjTgurhPwx1F2SByAJD4M6SGonPDIA4AdEjw69JLYlK/fgFkLs5MPLc6KJ+sE8NX3VbUOc
A8TaHORKWVBXOkmg+lL33H16wNl3X2fANheIXcwmVaaJoumCMPGVoCTPCz7EmFOOdeX985hvROSK
BCIUFttFWItlzI5AThNNp0YsVGBphUQx9V/vN9zYZXjKZEK/8Tu4DD/w/UzSngK/KecUax+NR/ZN
Ez1IKMhEM1/uVfN7BxJmDdG6OemG0RAyNP6ZQmuA5fSfv8Iw/rKjdqc4RU8Ky53TbBZcX31g0esZ
izLXXsPLxMPXLuFMjF2eYSegKfEQtgMPUKYGqM9rEpERNSL4fRwj3yEFSeENiOHqhOW9OfxDGXv7
x2PwQ0/YwUaRRKA6XKrXPuVNh1e1x/BUCizRu97RuWXQiaLZ2WX6XXNGW182SZ3Yt5K6D298MER7
CfPCfEWQxszf4NKZseGQvE7flXSeer9WcV4dTsPADLmOZSCzv3upM5OrnX+VflUnLMw05mDWn8gs
ISW3KdNphd+MzAmnwjvEkXiNGeej8bE4GFqvtc81Ik0J34Kyr+mdFtmlc9JiMF+f1TCQvT/EYbo6
1sYL8vfLLAFr9cdq2vrWjCfnKFfQk8RLbYctoXYee7qI7EkUDE7o0DieDT5Fsmen1hqAcvB9DxCU
r5vaUukTskOCbHjEa3C5MCMM67qYfOXPfn+VTE4Cdht5Y9gg3lqsbbAjzExITQLK8fXoVBDFVqKI
Tmy1JnrBxsXy98wky0iaWwssGQLByUwOpCzumQTe9VMyVuwZMWHR2guYVF+O1qYKAoAgkNg8zc/e
RsYr3dJTCL7VfAlyx0NlcttNEQ2AmoqiVqKeCaryHuj9rVUdkobSTswKqSW5wiw25EbqDH5h9wUH
scJnUUOARpOZ/45ZcoqtHwzbz1HrCIrporqQba/o1uwG7x4IQyXkjyRFumsCQ3zpSnG8lpDcHD69
wg1Wgwy/gFHtXsUG4xrMewHbUvbCfNEP5QKePzGjIIHgtVL1j4RFGN1RMRvbpGA6Ql/47P/LM/43
dHiexnkp406cDKxLLb7KoHoE66uvDjZE3qN/OO34T9s1X6Nc97mZV2DJiqSm5Qn54JO71vW8Z2pw
b4zrTt63LSsjbIhmeiIJ6DHk/VMjrsdIy3pL3cN5CzJ0bGg6LNV6DzJ8REIMyRTtBO5YeXMrUSU7
3ZGOuAjfdK7neNmsSC8pkTDR945NdD76SRFG0YAGe3yySHshqlWe0UCyq0jbDA1XXfubn+chkyoR
cAkShhByyGDOdO+5y4tJaKT6be/diwqOKw4YF6ouNyMbaijoEYfHVpFJ4/GjfDGqGPw1G7iGPCnK
jZ5TNJ4HOSU0uLobZCr3qkNelsc7UzIUQHOXs/yCd1SSfw3lCMdY9WQN54e3z4M6uP4J47optgi9
3EqzwWLnC8TAbdAph8DBy04tbE3MFdDHmj5qq+/uvlL6XYMXh68rkAg9SIK8idXdRDpiOUDcWldB
BRVHHZrD0/MMu48kplYoT+nWfWVdF/j5ZSK/2j2C4Rdx8bQShs1KLyq8LuilMFhw3dWMyxdeRPmC
/JwUI9bR65jWAoMl4lEshQyX1St9CMaxmLMEvqpo0LTgGvAum4D/GdbEOG/vvpGd6p4cl4mJHStW
+Y1Gn5olucMBATKBQTHhmLxkyvGOnf20BK8/X5tPZ0FL5X7oYtjBiHDV+kr3FQeOswVfZh/8E40q
gWKmoW6OxxdEObLm/sicNh24nCsLCIriIlszM3rDHSRRbZapIkKBDGEcbTUo9FO4rf2Oae67J3x+
kkoNH8V/H7it390A/XTHmtZLVOEH8Koq1qNr2VbiigJEB6LQD4THTD3uPStFTb+ffhRVTn3TtJD+
dLar+timXR53n1+1QoyRlR0RYsYTFg+NPkHu1D7Jc8OjfGUMm9o8rRLDC6hSbf6c6H7M0893mV6S
Baeh0CNRUKoYRHWAtlyUzqYwxWQj+lxD6jFrlpNoSeSJcSC/lhq/nGsdHz1xKrYm0ubkVtctUwFL
ID9PB6En6qg5M8g4rKnKZ9Ou3mkeTSw1ERGk08jb8k/8OesrX6PAE1m+QbFYiug7mlZ79aOEEjdC
zGGyulRNz0GPfsbpwmMUvqoLJHDTvsyiDqfQJwVjfBKrgfKxvoK3MQxss4nuWpbYnY+lkscGL6a5
Qw3n/5tv15amN33M6Prn9A2d1F64R3bpbU50mq1Xq591dsSjj9Dso1TtpdTomgaMOV5e7hC6BGIh
lufExMG6/nRFcqJ7Kq+d5NX96SnaM64iFn3eFmoig5+JkTLtwIMlU8eDXjkX6swXyr9bbs3lQdxG
ud6ztM9KVTbbd/ueWi8dS5zjVmXNylO/CmXvsT3vxzLRVGu6q6L6pPk/DJ46SK8kyDFOplj4T80M
eTnDhjDNUtt5B3B+R4dlsTLLb4I2N0q6fVXXlEeZNlRCRNtyukORkf91Fbm7IWAyiMHidhrVdeIs
GneweNgOQBxszIl/ZE/X3pMnm8b0eBXhcIgidE9ZPmWyobJK5nbJOPmVNZES8aRSYtujpv0n+boW
p5yC1oAKyC+EjNKekKWaAX2zguCdJmAjgdzPVLcYHMGInkxJMaQiK3O2bqGuu3gubrWaKhFbEZ++
Dvz1/uLoF3BKbhx2kJ9iogndi/AnXNRG8C73JOckOEmFJScQ0CWy04Ts/Hz+p8Ge2eCuwU2U2eEh
TWMDE9fADXU3UeuAmQbWhHParLcvJ2UfrtAfUKVplBFs4iBmEGddes1zYW7G1TdyLRPQbU1kgSHm
zrG4nN+Dqn2HywuhLbdm32otakgFa7g7DMZ8USxryxC5NODxXHnPESQqcIUZS4vWowNTSlj942tf
Q7Lp8t+6SRfFM6jzVhK++3pkKsbDC/Hjj+e5KZN9PThFa4Rwua1UJ5rJX3eHBQGmiRQ5VAUIku4A
gbb/1dONC8Ni6DfseKEtSUBoA5htF/sOZdiP1koaiS740YnOGkDyrtS8EQLBx/dpaSJZu5zfg3n2
5t+V5Ku71p2I6RxO3CQSr+7O9PW+TWMTihmuI+aix9L4P762biFRDGImF62vX/imFtSd7qMFI6or
18MiTWZ8CMfkUUPRf3RXOwCpqIA9XLQuyQ3tk3uIV99Zs3PTXvC6Lv5cRmSBE2+rjY6n5NLoefx6
j1nETII3ivArN1Xb2CqK9OTdaUiyeuKS/vks7jKEkom1yV7cri54se3i88M2ch4p9AUG2ytZ6hJL
zCoDOCdUtOb6q+oOhm8Jo4Jw3rD+5GsgBjj5la8RwsNqQsUdAndra4bbEWY1tjg69cxLaiJ3eCo0
mZxvEFMFVhr6fHjcfrDXwRTl9THKcN+evqeJUrYqm3tbyDeXPreh5vaXUu9j3B8lr39PSsRXDvfM
97c6tk0SMhTZzaVKRvSmgjNi24VH83ngFcR2j1NozPNYwPGmsqZPLQFa6GiQaMpYHM2c/jfv6pdb
U9azP0gbtF3yQ8L5SbSBfDGuJKSXUiay9m3jzK2uQwp5ltCGteTXaJBBr2+MIctnrQmjep6rjjbE
+Lo0ls6cRXxy/zc40UWrxlglTMBAmfbbgpWNGGNmTnsS/l0h+1CXPIst8gN/pXlEQjoCl0XVH7z2
wTM60Ik1T8qdxpUm27Mo9es1BBE6At9seQzK6Dx1Fv0KO2F1t9/W+hokdiRB1oBBrj9N5VnZBY4G
E+QSZ3g6AmWZAdmgXMSHceVS/g6C+HAv0V31C54M4udDLRzdv1iAs3wirij+oNesD4w9qTlRSKCn
hyB017ZSJ5XLkJtg4EUfW3TZX+25BH4Qp3tPpipYGS1Q1mCEzuS6vXnnVUrb/aTpkwcbygMDMJFm
x6jN87ffYPT8tETrUGl9Nm3tvC/ZN1PhcjhSlD4OsNb00kFiQixfkw8nfClz3bjPxiU+ykazr0db
XVgJw01N5JAoFUkGDx3LvCDrsfCPLEUe78HySVPhoZFQBlIx8fbHXRv2EWRU70tCGX56IXGxjH3F
rCBtp/vZsbHgRGYCePY+dk1+tOGkSMDyWCN8hkTuIeogChPjOC9JLMV7ZscPyyrBR293iY8XlvDZ
LSY069Tsw/RuBvmDrYuHnLGyftuShNUNGZksbqxHX2poMHm6gisbM05osC/mi4rTJ7EoC9pm0/0J
al92AzUZNzPI1y3cRkrKclauaqXjkBEbsDnW2ClCzascsiJKm4SSVln8HpZIW1YA2A4cgEsKldGn
y83FBYlXEIZphbpREwD9gQBFH7GD/EerjO50P1eOOYrANRVXDp6IROg4UdY8SHEskQZ4Osrl9SYO
wmWNs286G2SCllyayXq/s1ayF1quyH9HsHPe5ibIAadGbUvKDCwNy43s9zcbE1XTWGReGylXQsiY
R4XyQlLt4sJsoSmBOUF1LHD0uTQmXwDP2klKFE0KyE17fQmBeR3i12179kKMXtaz0HhJUoO8iINF
cAcVMfmIai7/r3yEYYzDW8hsHc6WqXxYu4CZzH9jiEMtAW009SXkcS25We1fQplx4qcboNn+oKOx
hj+1mcegqBxdmklTIdqbYqzZs9b6EdiE/nfdnOazroPfG9GhLP5AB43zOhZlOfj5a8Uh/k7lYH2h
gv9s1W6/kSsLxCtJENrB9tCry4HrPDDNnjWron8pFPONPWYxMQBRpiiwESz/f3oihjPTnYl1jkUe
D6XOCkcRiBqMj1zlaxWhe5Jv2ppd5AKIa0/vXqxDQG84V6XdtRbw3Xm1OuF5xqW1kIS/rp/WpFQS
MJz5MbXyLGUm5DWGoGWKnDLMS3GXyeAZcqsfoGsiImse/1DsWLZwjeRAwCh/hxdXglNrNRqJ2pWm
VpNhtJIJrQ4rO3NVbPkxQqhsd2NHBstIJniMd7PoKBiDdgSzsUTHpHvRseTGcaj8xji4Dlq1UBm5
xL5io6Ci+52WLZLod8qveXe+u7DSGDWYa2wDUpQHlV38l6fWEGhuhQIFb4CfX4tJddBCz335Mvm1
fV0GBpucmwu4BhJJKru5xjqe6wGtqjlGg6OZhU9UrIBAVRy2cJ1YZixTXrguqI0WWMyev+TZgHd3
0lpVtTRGkDfeP7u5Y/23Eq8TzQAxq65TLsbGIc96+8bLhWNnbpRJK289hOisrYHpgAVdANPRsx4M
5T9nYLhqTUPwZIBdB5BAN5GyWTgwr8qACBRhsz/Wmbu93PNAUMrjqynNFfGXZq3QjKAhdW1R3UfQ
DW0fx07SvaF4BD1dmDg+zyADV2xVlIrKt7tLrwxXL8e6etizKVKYskSOfC0JT7dr/8xXL9udeNpo
tLHwfwAx46PARsCT781BIBpyx+6U2qUqk7QrBLh4XlTDvCqqe9xjrNyWjsGUJVgv7t/eJPATfDoX
AhYSxkKKAF2cYLJWQvTNtUdto/KIAZQwUKJI6MW3PTMqzbXHbBsEVwGGPHJIH3mwl2t3Pck6UGlg
KBSmgRNfJMK1mwDbICym+freI/8VCpjdecAcuJgi/w+X5DPSxZLIYwKI4V1cLMJNhEus8TvsSa/2
7ZkoEbtW3XUsvd/JQY+CcSmhU3PRUSX9pVviObPk2GgWJfgzW9zKUgWnSM9yPPZRy7P0hHstrTWj
z5NJxZKy/AE0bEv9e/KfaVB3ZVpm8wHwYPe1qSSMOhmAnKUWBdznfitvbowLwn4w8BYy8Cooxvqf
y7kS515DBXcGwb8DaIOegDmbgb9t2qV3/b7lYTzUC18Hd9vToJSsnTkG31OTRRCz+wFnWXx6T5sT
ZQ/GrVXnecZcrIqzgSGPt7tZwR6idjkRqzfveapxqx5lnyRgYZWONfAlfQ0LQ3YLwb/rTMn0tGkw
GNS8gzo8zXetd4to9Dqoo5XmmychFgJWGoQuqnHlS8Ysc5Ox4wWZDv5bexR49v8Ulf1voVinYy61
n/zSVnyTTXwje3s3Evt9CjRsJZNhLRL23j/Yp9mOgwGutrwapkFJ8rJ33YqC46KMLd5bd8HeJxzw
E/tWzcSjfZCRfKIQCrEa0rxzcJvd9E22Lsqj+G7SEeuYDc0yvkcWFWhcLTfBAkTsVNi5pDPRUDkT
exk/Y5gZII6HP+xcgt1Al1B26vFLz3K48nPqec8HFkphnLcJKyGm/O9sS+5e2CYzhKqA+D1l8ng5
qOL5lA0vH4wBGKAloiEB1RpBeClgy8jHd2X1wn8hIVLQPmi/Q1gII++q7zNQOTikM+OOsVRTfDAU
XhNGmnYSm7oxeXiXQmNSN2WiWOG/FuBDNa9nIJzlJA/uvVvzTAj2LvV09khfcEpAY30DnklXp2on
2EWszp0XX4jd17LP94moNGQF1A5oXneivhiKT52hb9btufPSPr8gu9jvQrF4My0Xdpkbp7QUeovh
DshSLIf/dFS1lxGkVHMVwcAp2R9z20yvZS9TM1nb/A8Vm+dFEtZJNw40B4UbY3exaP+6oTTvinG4
U39uJOeHPozzMIFkVgbH2cn90QoXRWYYBtivJsEP4pG1Hdfw/SB3in8spiLbcoYa8tIDA0OOs5pX
xyQKe//wWeZFq19RTFnZGqjx2wkKseWUEcKq+6KUmGf2X2CVY1SKu4IAdPDhqoKf2MBQcU7RQ03k
8GyvC7F+jf5dkasd6/yLhu83CErqLnpehautLwFl/BXnLshU1dBsPaTt4qgyw4TZ/gM0OAzxXDw2
3sVS96lF2ad28i/riynVeff6cPmRYkoKHOzA1RH3Kk6aGlu7DRnesBSAf9NsOoUlDYqQvSWPZsJU
NLAUEsjWxCSCeahT/3ZkKueVeDIb4scjb9G5F/Yk2fWwMuFcg1VwRM0Mm6BREdMDwez9ZKeLzSXI
DtiAlUcSrCKuzSWKinfEeYF4X/UvoqhmiSbZvjAy9nBxiVxU9Rl+QoUsaxcOVIOfR2szRGt8CnaP
fH4PymIOmYA49HaE1i7Rno7LGoX2yjeOZoP1g6/C9IfUXMp+NSojbeR70Vo3wEzpeV+9hW4pTj3w
jYcJa4VKX6rxH+I+U0fO1dScK8rRDmZduDQvR0KXEf1mSLW+2RFVDoBcvsFWR4oN6o+ICtEFftEa
e5Pbuj7w8XWzSz2byY/fEvnpS5oe6KOoni3O5EhzzBkHlbpWtxHPCGwJHAF/J/cI2Zfnt1NSSo2T
idSTuwDhA2spImrOcJwZ866cLXQp/zzvREc0T6U0z3YE9wBdY4ns6nhiNmLN6+xvgn6wB2BkFrid
psy1M38Yo7sgNDwkDzSG4p8TV+zBSVYsrqBFwmOpe6WCe4pKXhtxTMpIol/HTKlTE5XmIpi1fat4
3JeODc/+SnbpKxPddAYtbwCP+wcrajjakt1Zcpd4LlocOA/raGKn6bBXO+WOG/BAolevh4luhHR8
ZfcqhzDsiFnZfPQqCbekHb+rpG/WMFUqXmWzi3Lq2TVsQ/W+iTTi88OSIBxUIDN23IAurHx39PB5
+Tx/ahK+zGHcri2NUyBnE8xyXyPaO76WBrLPLURvZbdaXf8GxnwaKwKDAOZPVxI8aIlF1yER4/m5
QaeKGlp7XSHk1XMBWYeOHTbC89xBmRE++VJl3Y5KbOg1NHtEsQbb7pUOhot17lzy2GMrRiXgVZBW
/2VqxV+RjaOIL5UhFFPV5htgcVXD9RIGlF0hCxkZjtLP/1Z+F0Hu3j3roK1Fc+nnWBCXhh2QMO7C
fGEfISm/itOuUl+/Bsyxo2+BAC9wFEhtX0n3Dp5Kbh5qpiCZTxYkR5+GHgNpzCGP6JR+NdftHPSb
DmkOLFOA3DSIVwhp3Ttc5dmYpFxnhG9ivqMs4v165KmOIKhqeFuoefe4YrsEG08FhH6wzm7K8S/0
q1wq8nc1626/s6sKmYy/dEGOuOSi6t3YCQ5/74Bafeu+CL/yZC6PRi6aHK+0YVc4JmxpoUN3FEIX
5UB+YmauzMa1Am1UrkpnYunMVmllYAb4CGc/SzRRTCzy0ES4yiM5PE0mJAY08OIU7h1Hk0udny2a
6AKwCJ51JKdjTFYwe78LeOPm4Fig/XdZaDA4QBAEEKQcOhvcyRZdTaeFcKofGUHmtgN/7rlNbrGO
+Ret16uaud0vlHqL9gdOhR9xu3tZlXii5sYYdvjzWc6tcE9KnB+deMgJxPZoFra2HrpuNrwsYGOT
zV/vhQIX5GJzIyAfAUFIZRPwQIC/h0aqY322viS57Y0bmZcYHvrg86qV/oyF6C+ih8ztPEod9hmb
6jmyQ3j1yPbZLA3SgNbsxK7VBEl+Lyco0ScnhwgVLGs1f/hRWCHECyqEyRqzOptXNCfNVMn+H4Bu
xtbXRm9GCxQd50RjDSsJg/yVz+A6eEzXECJr8IjqAp673EwuC5yhU1LKV/RZqqkKZdx53JlixtmA
jrd12di5ootFwd/YRP2VTgwCSSswyLt06kFBA2gh7DFr/CJYEHjjTHHSfXB/lba72UTXp4SW854k
onvxglJNvRPYbDseNwquE4BrKvCwCs2b+ynbTWVeBU6W5Q6TumlHKotoKw2GxXpd6moa1eEHiMtc
eyXBKgRQWYcYFCNEhvbOLnbT71k10XGwo5Y16BtTL3M9lQ59LUIx+k3rcFWroO2twtKQX6Bgorww
lVY6riEPEgrPB9c+nY0+sa8DkW8KuwK6T8nLNJ/IVauTso+IfhqpoSI0ksOfprgN8ODsoRsb2VXH
rcEgg83vyCXn6Pvyn3xeIXV17Gpdw6rWtJU8m1clZUXMGdBr59OP4wIHXhGWf02WyBD5R54V0GxP
NkF4K37w1Bbw3t0KC2FtTU3sdxfuhvU7kABX3aG9PTJieHtIcpyNMAKBa3wBUHuxtAL9Eu/z+tJn
Djvqq9UJDhWfy79oIJwkTWmoCzUdABrUNGWYpwC2556XJHZU9U0iStc3fNXHf3OZ4vS6/G5ZIel4
WfUtkHBdb9NHoG02t5CaSibNKqFo7ilzaVGJgwELUq5GIi80O8Kg/OSrxwQLJ9NZY1cs8CW/UF90
mA8Cyo+Tgz07ypoMHvaz6gCtqnY0i6YhxVe9REZkxFZlBjC+fJHOAbjTnvYtNvzOc/sp7aapfG9n
2xMthi+lljq0j/JtSGcFEhMzsDmISUDv/81E0quUnBv/MCYDhWSQ3ALXGBp5tpiPvM/ibjTfT7IS
USrlztH8kXd0iU4QB3VjepiZqVTEaQ1ZC1MvbwRCiYtdytGQw2JLgrGj+Z1CkJoCEAMVGfiaG37V
OGJhxh+mLSTS09V1w9C6+pdvH0eFx+FWAyGRdT7vu1M2hSXvH8IURwKqMGC36nDoYCOm6CTrphxe
AF8wOQGrxjH2HOyB0f4JvB3r2GPJf345hwrUwHt3ZtawOtBIevrMCdEJdzfmo40DczQVl/khK24W
N+t4DD5QgVFGLK++K6BVOJi56Fj+xSyUqDXAMqfVhfkPXcyHWLq2CnRTDd2D3xrl7O8wacDNWB4R
gCuLmGTtVDwkXWuCCnC8rWAbfraljAkNvT+HSyNrxnk4qBFJUqKg/3NFyTzNMv1t1nRRK6PzDsbI
FVePbPHOQAX06cttKwEsm03zMSooEQPKgN2T4LyamL8+7/3by2rdo3/ZKWz9z9zTA9swt25llulC
1ojoUWA4DpRSffWf5XE4sNNTcpLyCKYcKNmCjRa6PPBfjcPxL5JChlxQZYQO4Jaff1fJ/9YcI+/7
kVmvb1fddmkO8gtutIx6RjsZ+XAQvBDYtDksWeqPauXUmibz3mkbpSN/sJjvkvl307J8kCFFrvfw
WKQ8/zMwOFTXpAO8Y3Hwd7cXITSFUpXSpnymwbMFBlAj9jNULTVqyOXjLlodDk+kVFyYcebouyfk
dBUvMS/2cC4LZnmFNHuaQ73nWhqnTOKANyGA97imBbC1d2gn13wZZPnRrkIZojBCiKZ75xGV26yV
8hkG6+Mi3DF6PFyE/+/3uHIUjGN+WrA98uZsKaOJYWX5qDWkBqgBhfI1U2gHaocW2URRhi2UdB3d
v2Ur1P9feDQx0VdyM7nAGwNBrwpevmiLlQUAWH2ZJd7y/6pCIC12KMS3j+CgY7+npLvvfStx03ks
lY0paKZDQSwF4QUoszdcKI2g7xW9GsPbtOI4asI9vx76AvdqrJmI7YfOjsate8B7Q58VcyG0lgJF
bxUcQoRJ99xvaPl+n1HYNY7ljdJFUGTcWAj2uqtONiV+rnI37Wg+MTUws5hCsQ2GAWyyaBjli7OI
Txu3zmvVSw8MvbkBRZzAOK1g8KPvbKhzYHL6CZ1HdjiVRAqdEO9PANk567eBWbx0MgyS3mVWoluP
3hh2aJoXZSWzibZbJY8MfAUtf8ZfgKsRyPnUNK3VPIUkXf3/oZSd20ggihOsBsvh2opmHgoCZC3k
71G6PYOJ2Plx3W+HAKaWfwWLg0RhOxZ2SCYeYofRr7OJop3/KSMDmLVID6tvvVLqCzKic5Z/5mcL
3QC4I4jdpdVza2Eeq4iSXsDrwb0/uiMjL0tA09GNdbXHOSdxZWRLFbRXdIN74iJp7yTsyavrqUJ9
xHXl9iA0L9fD7ojV9ajgJOSRKfWOk2LD5kkTqVVd8YknvFZnjXnTCkQOOTmfqq1QXssApvM+1s8e
oBtRhIOLk7nW0/R9zyYNH68eBdNbQYdw6U3pWhiUqTQLjg+tryBWshNiF/XIuBk+A9HNqD6oN/DB
I36Eojlw7N7GD+jPla57mT+4wXpfWwkppuFUK+GOJXluUwVCJXF6W7ssbtqsPHZVkoKgTYZpLzwj
4HY/HWoGWlTdOQ58T8tCCWLLofXochK1d2wDZIXUFSKGxnkAVn1veL2nswjZe1MtmlloaW2kOq3v
3UNJMjcwsYV94hVzve2dekPmYIenN0owdStVOx9Ge8ciGSWTZDZWk0G612mAUuIz57OMvclgQYmY
w17B99M0ru0eeGxiIZzTlOuTA+FOg7Zph/e8UifMJR4KdT/5aZrAKxygE02CibsLPHe7PlW+t0iv
BIN6F3x+dPTjxASmbig3EhEj9UyAwYCSWWdQpXA6v0PTHHN5l6una7I5sRPMLSIWC3ldDsflGu8q
Cb6e5F7tVAQhzRqlnFOd0ZccnS2sjIix/RE5G1lUsAuqD8NVtnRKl6vHp5e1WlcvIwLWlP1yaMSJ
G/bak6OvbsVODDQiTT0vjeYQ5l9x6PcQjqo38lOs5ianFd3tY7Wt2eScuwe1QWu6p8GVIVkYkYj/
sJIk++ivejnX2dnBYMmECureepkOprdpmUM/vXak1I+7S9DVtj9mcMPC521ZJSMRb74+EVSxO3fK
eS5K97EijZ6+lefYV9GvyYFoiLxIVVBtCrU6RTJzNPxZLQnl83IqKrcf9BvETXzj2LMnobR1EX+q
+qbvrIhuq5m40ExGSsmCGn0XVSBPy1MNfvuriicjBWTEV7M1PE93Teyv2qB7JfBT1XZ2wXJQ3+fd
t8sFwsLyAuHL1Z+NNZYzTQoDYXDmMLy4mk0o0p4uBvrL/LCd8HjCKX7JNPpMMej2JoIY9K6rkMx/
eDMqTFQjFyJNXjWEno10EFtxISP4q5q1d4B1J2k2Rx9nXr3nVNnRP5wKI/tprE/HqzT0E/ZpnN5h
QcdwU8SoqMyFEM96f4sRQOhDcHykEsYfBC3+HfoOF04xq1RwRgIzxAbyc0wVRwfCJm9I9DFwyh7T
o+Gc7KLS4Fy7EOQIwEkS38Uhb0zeqTXiofNIEALTvzuAMB1W3ZL+H3L7LTy71UJe9dEu5rTg9pQB
VJTtyzB4TAU2mmQYp+VL7k9rzsim/fKEvRpa87+iw3F0LiBu+/CM+vE5TIMt/a8qP2KyqZSKqrLl
BPRq46aXRZtzv55uYKBJcz6tmQfXc5L99wftqFR5lrdyaxCOklrO5sHJcqdp2k2WQgxDrYsi8+sP
vDRCCXsCbOeqEByr7dpf4+Mmls7hYtf1+exl9EAhwMryRpUhURHcV/5wH2q3UVYbXOgV1zIkKI1a
5+aPQlPmKqzxjuzi4xR14h0z71nYgAwXvYBlHsljZ/1ihDqgtNLI59JwAgZ2zJTqfZcxT/h2O5Rm
CQnzr/+Fphadya2wuQbihL1vHdyRaR95V5eh7tNhAHQnj5zTqYtiFjBQTKZToSuQrGbH6lUQzAyn
0o9678dc3FSiMEaV1Uib9nfM7VaS7uYX7Gr5IpFiV+r8KxbKsWcdGR3WQ2t0ut544Tcucj50khFe
Q0GycJqSjW6VNNdYhypU8Q9UzcMOh3W6+2mRSyWS+w1zfyrTK4WNAppRL1dtZqzi3TvhIGqztEQ5
zObNBBzcUuoPUo2CAP6failDe1fYDRyDFvcrrU/cYIsMuq4UaQFmTDnF34zvV30rM6NCEtIc4u9S
oEnl+ZLEB6HnenXbjETyxMhE1TvRKtXHKm6cmIoQoxn9RfEJjAj/dNqj8xrfFXFgTZSjnmHtHoJ7
jW/jQBV0kHbYroiB8+GfX9O+ZOUtmW808oWVQOuyzYauG18B1L4+ZjkHNZe+HxiB9W36NPViiWzI
mqen3cP3TfxpLdkk19vx3gtP8oMPsNg3VQiPs7O+gKjenTlFM11JPR4E+dovYBNV9EAKQtbWrxNe
Pmb+YzptgXK94hNSax3UVW/vbodBSQBT/dEeXINYbtXUhxEjw1uEU9vQyH8xxMFyEo8I7uS7PZSv
gTnP5rcyHQ7IzOg84td26h/B3cTnq1g0KwSrEDBDLzepLir9BVJBgrlzsVzg6GbLD1PPS6uNBzrq
843co2WClulwTrwzjxVVOhTQzY7DW3e4zNVC1KyOemDkxvmnc27nMOOMUQvktOEgOaY/yC2rHMlh
glWhOAoGgjviLz/9AHnvvfQao6pj433Ep4VQm/HLqmFNl9Kq6jSf6OsBjkW12/p5IzbI/ylQCXF8
aH5YdZkv0Q2kXi2iECY5eJVnFXPM5JrECU96K4jX+cDO+EARdq9VT80gu40fx6nr3LGi3mCOuffu
eAOEAPSfO0R7fbQdLwogXQLbQYwYsOujnAvWYx6Jw1Wanhg+0w1cSiwSWK0GK4duXeAVgrg3FNNb
/r30PdY5o6LzH/uWi1OwNpiW72hHRwmIeaeVHpE8lDkqBUx7/gzOzeyVK9Ii/DcjxRw5L3+rPs32
zErkF/Rx+tEWORPWgNOe7lC07k3CVSdg4qH/y5Qj6jvdvzRVC3VHIGDMkGp7p0NDMoWfK55G5p+P
ciXo5ZI5ekhOWZhnoivtg4ZmSSktKit9Jk7FcvYrCdLdP4t55dSpb/HH9P+5El5wlB72b7jgKzB8
qlDp8sXBeLfIs593W/lup+v25Zqj8MQQZU5icYAB0NKPfR9LhTso2NZuhJqjUjIgfBFYUiXOBnif
Yat8mUdOFxhpDIU0ukzuP+TizV+iCv2b4MZrK3+nHZXbOlzlJxDYPVmHyTx1yKdgq0Sv9aFSnhWz
n2oXt6JhmFCHYMGwPmFbyz/tiarBdJq0RlicnbsjhjoFzY9jqvP5F1qFrYwjouthMuVTB0DO6/UE
MUQfAhxOOrkCBMAqg48N67XtrBaQqm9b7TWPWJorbVUTIXWEbGvP2UK5wcQxHckw7g0BudS/ohnl
qlhso+/Dkb8gBxal8Gyn/AkyvpLZ8x/zO8CVG0PHBTMvINamPxpAiLY7gZiChzUf4v81QaJ+Si39
UBstgw0DhD3MuUwKbKGWK5sCaANwBh2tmIvKx8xSobohhoELVdkA8XkQ6O9vZ9+oeNFZBeWMkGkU
h1NwKj9Zq/TELG/jb5ltyDOGPVf7EpWiptp+N3oPBvlA7ttkFi/gGDiyq/WZWXOaYPOdeO0OT4yc
QAvpttTUFzfZ6cXwa60Gord/UsF6COB9GNblfUS5ukz306TFl8YGbeMz1Slp8+6BjiT4LUB+JaWk
jyK8ZT64AcPZD8cp/s20gJUfI2O70N7eiyFVGXWPkaWe7XoTWQCuhMrv4mmB6f7Uc1W+jobREx9V
NWWo6KZbjCDn6eG6YwhAkXYOf+j6EZXpsJlLZ1SMNmhVTaKhYzZ9Du806ttq+jFwoDtjUx4QMCkd
YZsCTUiAQ9gVggFLMJayZiV8Pcw9o5xoMwiKYLjRI93IyvqanRFDO64T/ocq4e9wHQ2MwGoisOEj
+k5EXX+mkYaeU1LddXYjSyTKRhvDm73dCfJ8MNcGydgRvT6cA1fbc2GfQ6rhGRWWQIHW+fzg/z05
eSoLvcoL9k/A1MfEErYCWg7EMb6hZQgiq1kK9+QUBcFygDl7Q4nVU1RIrXjNf4LaOSJK5QYyAH8G
omu7iuHD8LbEzxfPcpvZfA2UNxX5CWkIe1Z9GxVswQO8Myto6xVBcUIcBUs9hwRHf7FP4Dxua824
naGGssXsto2gFXrD7vlpjOFQj8OYVprvH6PVj69eAzYi7OV0/tBlDpB0hRhjmbNZjiJL7GuwAlpr
dteXoTiU2ilz7mha5tONJJA043v+h2/rIXD2yhj+Vrgs+kdl2Ls4e1DxhUb0N9x6hJfHGA+OOTP8
5Wm1/VK8YmFo9EbYPJ1Mv/IUXs2xBuxC3K+ICzBNj0kPs/Qdsu2/dAU0ku75iyRv+zNA8Q19R0J/
MkZYx9SRi7/T1/FiJxiW3QlYMDr46d7Lh8939ERdRZS2qM5DlXpbr5Y9ybKz3PfUENXWjtuh1deR
GH+geXjQnm2BM1uUBrxolbYXfB6PCAQutsxGHjX90GDvkUFSH6+liLalBGehq9BflUxHHCdKvj87
6JIJo/R9I0iY4Oxb2I/0CTK0b7hwHcdbHYtpz4qX1X95JdbHlw03R+ciQVSqPQeCDIMmp/YlvRok
oxTUMz38amMqxXM2pqC5Oc64Cz56owITFSSI0ZBERuzL6j8e+5Qc15y3vuA/yr4880stdjdfVnx0
XSeimS6t1omXpJuc+Yl43+Iqfwyh/Hwu3de0T0l+iRfb9Uvdzg9d6jfltt7UNE0VoXRdB+blCCBr
W0az5UWleT1V3i8Sgg+Ie4BIJFoy0oaMRSZWDWqE5+12FDWfagPu1lWh770av7n3gIGmrUCmZM3q
IQv9I3Km3YDPxAbVlcmE639AuAS8IdABA+os4zSFNGHSVBOgA/2upJ9+cJpyD0jd1eiPZ4in+UZg
JOpBcHa8qh13od+wOLwB5CJLutt9dBa3vKfYh16npmxBzF6XGMlIQp5eimXIxqM1d6XCv5Jr/C8+
b5TJlVt3/VMplvFlK6lTWtWh/fpUQlk/3Mem/brgcYxSAXmwa2UemSu2ZNvzrVx0EppN2SNDJ1Pt
uXQT+Bl90n1hNcHBzO59bpKKpLUxjAX5Zf6loZ1d5u0JgQCSgX+QybYV8C4ZpRpdaO7JWDfuCnwq
aFmLWukSrXda9KMIoof9gdICCpxioc3T8ukvVEQm7Yy0zKkz3267+6/5i5HH6SWLGGXqYEJvW4mB
3DT4zTy6p2KIyg1UUCLPfBoaS5RUQ83P3uBCOPbABmRQ4ktcutAJl86q1T38YP441NZVZX3mA+Lb
9rauquA4ail74i1v40+cWsdYwcea6JO//lR8feGRbhUrLevDWmWgCIgtUuiJzT4UWQtajbyAzgGd
uV51Pd838eoMFnZHkd52iX3RbYIMCT+f8bpw9G8+SshaI+FS4Ax5rp3yYCza9j3JTRzJLE/Zb0NN
PGBfS9mYWVwlK33TiKtZK96qHmo8kiYodZDhErARH5RBAZmb1r+ZbCvouFhRJuc5xC0fW8LNMznq
Ln/zEijY8/LFNJTCFkesKKnf0SUW4LQfQmY3TSaRuPEzxs/titW5IAchBpfN4rTqK9AMOCbRGE8v
dmfWtDUWIGy0uwQ4z6gBvcBIaBevXC+h3oJss+1dUDUdgykKt3BZtkcCHG+531bBWa3mhrS6epnb
2c4+epAUOlrNCLxAC8CKT6IHFSuLg4Y0V1DQ7HiDZfUmszegTgk8uVJ8tGb8nlhLH8nSMVRqX0Vz
HCQounaDengeE8t5Tk1igSnUQEsd3JA057NAc9d9+9T8ohdjg35SRPokSLD7ebmrLaAi0xEArhXK
2POL31gVIEwyxQr+iP6qom5nvvZQhd8eUh0qXo7Ob7vc7ho1Ipc1MK24w/DaL+wIV7mjLcPFh+Os
GTAaWAJKVtB5GKBdrU7P0kvO8WGOPuc34C2xsNHpQkPH8rPb6X2d5U7VekDwczhQtubBfx2PJFE6
hHrtPJcqM8DZcvByCvb7poy6loyoaB/VSb+b5t+kHGRqTJHj+gMaPPjGrtHOXselr5iuDJ1jOuGl
Ke/Z9yeVmkk8GD0QOYHiU1LcPuVrpgjj0gjuOW1umw4SIRqIJoLlY9KhGuhDnes1PqH3xq9ZOxiK
1lbb9/Vm6Jf/E/Poo91ItrlCpn7nntE8ntGKQI9U7nDLZ8xY4g3EyjLePX0wKseuLM3W8glZtQaz
lH+rxZ2WHZ8b4qh45PNyQkyPe6gLKEBoXceDiOUh5SxYBe334sVgFeeVsbeGnMIF8sWilcL4Vfzu
mxBDOdNhhP43WQZZFlhyrwKPOL0134XLwFDNOKH+2CcOq5HomPFzMEx+jqefyflE3dQGvCgTTP4P
Erj57EQwB/L5YQfhacdtOmQBcI10KrBQmUijFkFiSUqGlqDmZIIhulZk9dMsrGceXsb+xgya5kgL
u1xVe+suotd4R8e4lYAnvDE4BPI0TjzaCZ+fV9q1JB8KpYDfVX+TXcatfzwfPKCCJMrEydlV2JuY
PMERwiRzbeBwF5q1xgAqGDtq0MNWAT+5AfJafrLdRiwu31+Y0PnGTbmTy9FaRjpvMeOdzPwuGo4H
w8l37kjvFjrhknjNX3QXp9nPLHt7cr1lHtHLDnoNAR04JKmziGAupXOuELTdBINdcJ7xT5QTgcUI
kpy7IRhAaXlgeIUooCUpPe12vQQMX1uiva9UObM7VcAx1oxhW5d+w+cX7nIDLDWBFyO8jj9b7r8t
TmsM85/eE2e4VK6iuWdtkFrxZaF+VxheS5c3cFCRKMqyWfKSG6k8r+jhK7RhBrqQsIRz7v9cZIkt
5Opv96lVxLU/YxgqQBA0Mwn8fLyqFI9HR5d8hPVOVykWl+NAHFdz+srja+snoUgPTzs9ZsGMf0Cw
NsxkdtK2Old43amV/ngh34rxb9oUdsKIJho80XubGxIPaOPshtgxroBEzY+pN/2WenGTj0gWn2lp
01GcJ9deMJLI9TLjTNc2vPI1LzZqp9tbirwfdn2MoL3CORg/fp+N5XvSdl25uf1rrAFKLxOXOKt9
3le0527OG2gYVKbYArQFYfSifo8s4Zm8OtVLd0iunEnCbeiUIPklrzLE+tl8odjqamNOK/SfkexP
sNDZSmHCZTVyhLQ5lTRMb0s1NoFNfLUlVDt/TVFPlCVRBzC2LCjztaEwBybS0cssFHshXAoXviy/
ssEkp3Mcme9AAO0oJNbjJNmYrcBriJXeGgstWHQLDAURwsRNYVkH938jAU0EOob0sh3kI4V3udYw
TPFBCOhlughJq52AnsBRbyGEwBRpeNAdtrpHsuY9502ZZSSc1/20BRsP8lWfgM/HyWSWqYMNCa4S
7y1+aF1uBHYDY3m/W3UH3/PRsu44TPQh8j0esXoq6QteWbpZWwmSjAxJrLyBaDXjwmTGExeQ6ePT
e7BjUIJekRfQGeAEPUK5kozeOlYj08LO+syt5W5vlKdolYfIc2gzoLOdW1aQ1tjeA4EtHndgyK4U
49id/3vgrMu35nwX6pdQ3+dF5Ec9Wd5WCEzTB0T/Y4jk/IuMZ5WjvIcnmppyfd8TBpFz2VewFfmh
A8hJiEJm3ws7nsBqC7iA5dEMlRN7fKHDLogXXFM1w3MDSHuDP8WhK/x7KWVgErVyeGuNNMkbp9Ke
M349mS5NtWKxVlNr4G6NnGISxOYDEX6RMMDIppR/HZHMozY5FZsLc9lhn+nWLKV/dsAMKjJzTZKQ
eAdi+WwF4fRxyu/QIVHy77mMVDs05BTii3N3XI/LCze15gKD19nQMvLYOrtDRxx6Zm50Rm+N1uHa
TchOn9cLZz58v08eqKk6uvyagMgoTQAdyKf52rlnKg0CVFKxv2UcpNWfo7dagB3VL7O441aKza+X
p9UVs46Im+q9PZl08cAMdVE03uRjMqJiFcubqC8HFKMf7BY2QuCwe6FyLqitvliWsXR18y3j4C3z
BDEH6aRB0kHSKe9RCCf0430lTjaaT9rtmwJHPy/+oWxqM3o2uLV/P7azzyuKX276S5eP7zGQRKnn
tRcXEMZW1hl4f31QaGOTEF7pwBE7ExPIULisup3gLDbHFnbpFeWGntUcq1cpYn3dU0YWpdac7rAB
GXjFmodT+eZisxh1faY0AtrpVMF7K26vkqJ6FQKjtyloJp572knSnLQlJf2UjD4waPNrlkb+5dLI
2dnXWcv9szp7WF6wx6enmVgkAKoOYuiHYscWYjMwyPX5Url+EouADzESdCsLs8UbMrIXRVHDQC5f
C6NAuIV60ssaCKvZKj4wruvEPDdSvyS1E2/Vzsj+1XfFrMpAFn7RkP5sufbc68oPkR/qRzZmuEyh
yXP9XvklJRBqecN4elY5mREeedVgD8QgbnTM6UBcbYoky5v/ThUG1uyXrtvp9LqWPXLVVGlqCwi0
NEmq7qSBodqLgaQ08NPA8p2/fT/ku5vcvk94CzisTjS8TwnrqEt62uAKYgvbxiK2EpsmTPDp4HCh
2fGW6FLfVZq69w0Iv2D7bJ/SXJEE3qOu/MBYFo4i0EpLseO9naFZve6yZ58tUhJauQPrPOtTtRqf
QO2BZHGiKLdIEdCfYlYdz1U/0u5AY91VixbMzGJpBkRSGmlfzW8j70HFXhPm0EgH+UWjeiNAa731
xVwWZWP/dnl1lI9rOgJlnDYZ5BCXq3aWmai9reLcipY5R2D1wfYKje3VwXZdACkq1ADCAgjCKpnc
EbYIiJ/zglMZu9v00+V+A/aJWxHWcflyjg1RS5o1k/qwgYm0Ht28m9tCugrjhoe9aQfGJNJ4fPcM
0HyXkRpKGTrFNZgbhtyMVlzcZOb6HwuEsyntszF7HZyzXyKbMoVPfoOtyIEGiDoZxNjV14T2vUrN
4wtt1yLiiiXs6EzAc+0REfmoMtMArjq1fuFZo05//TXUUcE5MPg4/6AZWPBSMdEPVXEs+ur12Hi5
a0O256UEP5n2szWyQ0wboItwIJEnINDh/IOf4PmZ8oDG4P8ftpZbbRsZKVq8JFaUxxioTu/0rThK
tTcQ0DE2yF6YsWlplzAovGalo7lOeXO/Yb0gFwOurOFOu+fNO4hc7H7qY8/uuBLDhHU9oyUZvLNO
pAFn+KEtO4Mt8EVI2/e68p9LvAoNLkVY8wlSLnvyzNagRsBdYnjy7VrApDTNteURb29QuIP/e9Iu
yI2jaz8T54M465P1zKekXykLZ3WhRe9i2o64E0DCW9uP43LeCLWbCzU9buiJmrNkdWU0L/tdwmf0
DJP6+hdnGsALcZGB9b12+aPnFWZAJ2fkvIJJrx7l3hduVeVTE38XdQBEaxliKlDifB5olJ6cGacV
TuM5XoQdw2MTCv/ip08PN72r+ofAhKo+Fh8xn0AfpNObSMdneeHDXkHYJJ5WdG4aP4b1V0Fyt9r3
EU/4R8SrmDQuX64gnF+x89cwS0nvbnkELKHZSy56USEuR11/FJrfKMi0pOjskRWBbgvsh5dpfOEk
Te/Y/tQAfTwRP7CVBjkK0YHFs/Dz0ahwNrk6kXEmyROnayGm2f4rkLJ5gvIn5iVv91WZyLnCM0Ms
vmQ31XPYwn1OfsfqvX6Q8gznr8dEEaRMS58INZqN3iBh57XwS7gGpEDNadEsfpTN04qkX4t/oPmS
g8QSiJz1+dCfillTrHHmk5rP0pLdeJOHW5pOWWci9PnB54+Hl/SDwleB/mECWa2MueE0k90UxRkz
uGMMXQxqLmIVK5/WccaFab6t9HJ2idUzeS8X8ohyjinqU7+R7jUNreY7eTm+jNnEKsFPgxytt6ml
jfn8hqJF/H1sSzvrl3nA3mEzvB5yzP5pGHmDGTe+J6Hayjb71sodPNlMjbdmy4881pWtRISuUomu
5fSvrbk7Q9PiZmUV9jXyI5sJp6aUC2z72UQHMvhEyf9/E/VdbabZt14D1a2i4U1iBRxOaybBjHM1
JKTohfNmL4WdxN/paU2KtWGulE/EoCmJ4/urMBmQYtXRjl5tuAbxu7aUzDGElEmtlQE2JIIHaCym
d35LIC9WymTwYwW5PEXKRKfKkmfw6p0dpn1DL3r8q++QIOyq1kvTix69L1UhDYd4Uy6xwsliLpPs
E5PvICq5QdcXjtD9C3QWeBPXYNSuJEAW3PFLeXMzarrkCcu1BXfuxgjprTzGSL/ievarzT1gopmd
hw5HRj44YXnbYItozj6cGZ4r0simgc8NEnvrU0oF4YXUhRUwPlgXERkL5LHg6RxDkQA+lalkYjjQ
7ETTDJsyf4K3i2E9IXju4GbtAJzNsjdig7J8uvEi+SXuT0cM/BAm6WtYGHQ/xyS6x1AMpo5MzQ1h
eEWhUqtFl2sVlXSZYFeF2nOU3GCGfN8YZVLQ+/g6/3cK2JmTRAjWVX6pv5B2inWYSl+z9W9c7hVn
2SDnGUf79C4rmFTdwnZKHTDTIoXJ+/NlkoNjW+PzLlLWDgi1PS0+67OWL0K+phI3cDd1jkucbJbw
bFfzCBTzUDrFCqyb47B5EYT0Kb7AGfFSB3zVjJX6m+o19DCkv/93/r1bcT1a8FReMuW9V8PRsLxA
o9rV+nFyHBeD9WlKWqefmX0V33rLEdeKl/Eafxk0DzjjqmP4I87GL9MpbGU0JC9/mppETR5eV6Y1
p7mCbc4qddM8X9bBuyCW+cS+mZQP7V5LhuTzuTRKwPwunlXfy3whzeTbiH/0KrCmDCCRk8VPiF6o
nzSXlV6p4zkFJ3bk8hmqAIfHsWY/dsAkRD1e3zIwzh/AnyyAG04YeUWI/cP7cQALA+vHBjw6V2FP
I0Rixw/LbKSHHEKjVNVfwe9vj02K7aT0jIi6AiVf4Sa8Jla1XZ/zHXb35Lv7kspoLYIr0BbtbKOa
gCkI9XLNQdhFHq5NY8th9vT1IfmIdLonATPe6gdJbcPROJaig+drj5T4NMr6pA3ofsfItTdGU9YI
QVFLLGhS6ML2cJvay+aWEj/Wc42EOvy84lsKMHjjConTOago6pM0HtwyBeDuvBBOXVpBXLUZMbsG
KkSbtIj7gyDCGCNKIGgV8Xq/s0ztrHYj50w4p8Xo/kLo/JpkmHjwxgl5z463/1I8kmYPnC4VpRGP
wPTnacchizCuYpluNTMe+emxfpGs+ghsGJygiGHLyuaIgsvpMjTkhNxOOJlsURUi0K7CFVhKj3zj
VA4PY6Xnb59z6YKlungjCdXSDcdDLRBf+VAj7NBc5I03AKB5L8D+ueTOhO1d6boRYyzJanUwbu4v
kLF7RWNLGQSOGHwTv3DgKuDvaypkziixCoV6IdGPvc6qO939fAsaUo02xoCZMKhpG9vNH5W6WIAd
18pZVu58UhqliCVNk/O3ya7ee45DEsyBNychTdMz4JkQ3yr7bN+Vih3POnHt2ZKzV7P0JqhXuKSu
uZz3p5w2aMQ5WkqclYhLiqTTJxLJcxabOV91OgLWD3bOOy4ek+AYv+SPNL4gCtOfuxGZ2Q66MC/A
ycSh1Wbje0JKNjl1T/zCZA6dU2yvrkNxYExhbrQXv874MA63dKIlzI/c2r/VRE0dQ+Z+ytRUw6A9
wlIkp8BiqRZ7bR0tEF3Y1tF5rQYdS+jDbc85h3CJLdfpI+XTVAHR7NmiYONBOBzjlAWRc4TuPnb0
CABCFIOUumg8enazmfjzATsRmnBKxq01XNBK/rvq3OzRgVhKpWQfJ49fv2Gs3XX/bmCSdkPdZ7r9
2cR8aSGgwfZh62jWxbfgoSi/wFU9MsVzh7fYC5GBQUSZtOqwpKPp7jxyP+1Qeix3lIttDDOWVFBl
YltMklJNt/Z4+WyiZEqBzmNY+30rX1TPxA0+O+8BqJ5Cvw6ATQ4KK8neWM7uYRcbEj4ytxuujNHV
CC3SSqEd2Yt9jW25VRwPi2kWWe4uAfSZa+6/7+kjrjiTpI+NpjiRxxwrKeoMyXY6Kt0e3JFLs98w
lBBmu3z+h8SnjW8q6rLMQ3TFqF+ggubw/udZoO0/3vvRoA/9iH/NhiGQQ7vriHFKkUPsPTXnmTje
LPclsxsNr8NTVKHS2mxx+zd7xjcWZKZKrypeLgbJGRMZJfYOZXZBYFY9e2J1W8QTlzKQM/BMWpOd
/xfkhYALK5gtHI/eFup1/HQoF3qMeaFd+DZGJkknV370Rc+e1yjWRxwGPknkHdb9RzhZPo0fC95u
CiqSrRmWo56bW/LElc9MI7jZegF7w5V+oBq2YL1t1ar4xYzQn9V2r8rVrI6o7D19MU7xeuqt3kwa
WUGVcmkhsWWCH2+jd9/8C0d3FhZ6XfA0RNfQyYssykP9B0VOogJSv8TG6iQuj4UmKxZ76G+1aXmr
og045o9DVYetnldSLcUeJcMGaAwsS3vVRUkmvaegIIQGlgdGm2OdNwFavcfxS5IRBXxuiguu+qm9
+7Bc4aMNeEAA4xBxug0sD9RApq8EM3ztqNeB+ALhOIoeSdCaypkzlBTWRWeuiFUVIpoiL4AtcqEV
dJ+DbkVs/Ei9KGprVovwZARpa8tueDPnPr7DZKwb6xgxPkza0nSdWMeqt4PubYNqX3HTaQCHT4vy
IPY6Isv4MMnyo6qAbLT6sCHSQ7VdfxdT1tgJNFEUjXhZRp6kHNrd3oUWYgDYGrkxObwAT3YyCB72
5prIEIRCXm0JEoG+v5jphvYvlytB3syfg/TiqVqXowwcRtIEbCSQMGhj8EisBMW9aiui7quwfjet
mIi/OVshdGNeR+QfAmoc0gG9baFYJ3DqPzCsqEHul8WkXfJZBnd8NSkHjpKn1IVx7hVbKbmUaNkZ
gt79UYiWH7LEzAzQ0yADn/PxmI9tJj0qR9qKe4GaMEpAfshIPNGkMGCgTpMBrbAh66V2j/VDCy+a
o/azdvGhqwlV//J45TV5m5+HZ8/4pQJTd9DOQUM5yW9o8XLG3L4pfKn5lO7s6J03wodvwsq9D/eh
2+/9+5vq48y5tiBuEgRunGAHJXL/5vVWigu5AELgyITt7YQKRMd0Qw94QGj8rORdXUTQi8F7pMXA
c3c1T6im9svS0gNYXQz9AnqUQuFs6X4PFQhAEkn4TGNpjnkTlZahu9pr187GPrxEYn8P19DOVEI+
hN8R3hMhiBTtK8DIhvWDvQKCDN7nY+73r7ifioQMn1a/sTuYxY2Cdtq7apooMp7bSD37Lo9MuhCi
mehZjBhuuByfFa43KXZToE9XskwBPrs3CqTiKG12G5UeFVId7o54GYueZXSLvL7dvWHq+rDpFQ5u
zbIvu8L00VTFLx1kNatthQL8fjnkLE1MrjPilWC9EfA4SlGlmynZdADZ1HvY2v1C9JcoJz75RjKl
4nCiXPiEqwvfXsKy3acl/9GDvZpWNG7nkn85zMmvy/VCsleDHyWxT1//fqALhEKkyycF+N+YEOyF
I19YuxoE3jajlo0m8bhv3okVW/Ed0LpSWYYTuv8+Doensea9sWMt0FcNFCG5Ikdkm8l7FSvzmTaB
iFygY53b7jrgDepf4hqzt8/l1ZblZOmWVO1ML5u257ihGKHDfuNaPZcwQhpG0Veyi7kIPEruQGQi
eA7dFgtsy/TJ6H+ILQpP4qoBn396ed+iMVSkambH15WkzOccWpba9xfM0/KwDTOMxhWiUONA5Rs1
f2K2x8L8wnAez6hDnjNKbbS9ETEMLTCAkfV1XXHPlvSBun6lMkAB3IyeGnBgb2L90U6rbCKbkA9r
dEHqzvtXjTq5jHIAczPFjigvVh0v00Q8i2Ec4z+Vle1Hg1kYNOCJE3s4SDqmWSkHOf0xW248vf7A
WkCjIOarGF4GBTwICyNJ2rOd/1c7nTN3vTPsnDb5i7FdVsvV2K9RM4liGPdb5BoN0M3AQFJPXYkO
0pIDWcfQEYY0RpuG0gxnNQZoxZ0wi6AQgpQHD5cjB9WVa8knAjxGdU41F8JQI5aks+dw86tx/Bzf
M4haUfszi+AZF3uijSd5+kdeNU7dZ6oSA6V+52lzZyMSJQeqQSveMv0JKO89zKdXoQrfFEz70xDf
U70Ittc5yC6x0IokyMpxzFu009qFuxh87OrSwaNuX6nIvQHATnZRzoVVqsfGPwPiR+zg/ppHgk/7
jmljUrpAjpw01yddyHUQBd+j+8yJgbwhwTNKCbNlyBfYMzbUsJ2khe+X4YdTzrhr6mU7XMLAaq6T
IlBwE0yJQ+9sdQ4YRF3EbqfW/ZW5ObFSb+tW1GS04tSl44QIEjyf5uuHHFCDRzax1MlLf6LeBSDg
a7zUiyhc0jCEms4WwQSCAyYmWvyk/s7Q6WPAm6tlQjzn+HgBKcql3z4r+kBOboOkVJ451xFAdLJo
ezQ0an2HxzP8p/BCyj72tQIfH1zkYPZswqNuJ3BqpZiFwOXK3v3hsaW7W3AdpUhOCroHVgEbHHJh
gIhOEN05cSMuaU3JEKtNvt2Voo9eTqliyvY6w17VU40qNKKf18gsgDOG7LfFuanCOheJ+65ukzui
YIKDilzIFUP0OM1mZQf4OTzB5fRk45Nlfw1eKPFR0hjIkjOifsz2HFiQahpJK23CDN4TRsoBC5r1
/CxNs8oTcuKEBwx/RlNPefJNHfhECUCp52nF7OXfLia+4FWRug65O+cQKy0yXcpEJKwwQ9Vc0DeG
h3sgqpca1xBvq5KFwCKihA6067a0ceK/K9PY6nUcrZqu2zLhFbloMtCDRztXphq/wAadbn0lDAeC
liS9hoRUmM8VabLzE2+a1QMavGGZInLinvxpcbPMTeLOUrVGPP4zuJz4s1Py0QmLrHY76T+RGF/J
zPuNT9U5nf+sXsU4w+VYofepl0xed1bh7BIEYptuE0xagKbvvt/KSI2JYhQNJZ7of3cg1Du++SuN
PB7e07iu+lEb/rSK1IqjZ8rlNf/ULruYBujICByPOU4kf/iCUFPaHzz5LIhGMij7EgXEExvb30Sp
6axc9fxpW8ivviNzw79S6Jf1XdHrIkIsZzqHBK2QaFT3FS/oVcKyrQCTB7Kuf5bD8hbhMQCNKNJz
N4iklgDCcr6Y3t1o1IAVkl5+8Td5OO/auO0hI8TroPZQXm0SiuTl/KDaMPlblii6z0Y1mIu8spdB
uiH90ZpeXjsQNYFPlqzhp9xnRefoJ24uGpW8iUCu9aKAgzWK4YNgrqExPMjqDwKlhpwe1u293PQj
Iq8zPfTRoA+eTuQp4GfqshOfO6ZgzLchl1PyHSBeYrenoQH0zuFFRY3aX71B6d8gM4ImL0g0oIfa
5FbAJQ6hYx6d+HvfugU7ErfFulFYdEDBSenO9o5Is4tUHQVSBixuBKIdpO6B3rincCTVeWqmCDU0
LTXHNMSUbMEVzAvjrGAbfF0Br9Cj0WOrgNPbmvEuethLordL/cIEfeFZO/u2eZooMUkB+yQEoogK
vgRivpBPZ98XQfuOG9Di9lLhhqoypZMHjnUiX/GsP+P4juHaPfQjFj4PjnpefmOCVM2n8W0ZQqdT
4zX9xkltceQihDxC4ZUe2f4L0a8TyC8j6XrFF0Q+Ebb66sdVKyp6VZWXQfnaU291ZGqv8/JkCk3u
Npi+J1olfIAshi7vDiZy6pd/z0ATYI7zUhcm5YQPtBW2aF/uaJJP018s8CAczhXwKLihRgu2s0U5
3btJaUd6u6MWKKlikuB9hjfnBE8jULpkB2OSpPzfjFzmD7ASAqMIkLNQjjimIzQar4r1SDglbjMb
FzPE2yKzRCy1wQsmZArSmo4MGjWL/CHVBXIL6O1QFCoEEksF68t9vDvrkc2PQNS1U8QuO5CuLZ21
MjyGM/XWCEYBD8QEisKC2om4xVo2ppvY03rlc+eeIp5Zu9A+A9GrAgquNSi0s6G5EJNLsIRlbsuo
xOUE+L//udijWNCAGShjoBa9izNtV4vLFWFDXKy6MTvem87qK/JZdWt/wwt2US7DgXh+nE6x8lzn
2upPkzN99Bq75gx0KLb7Lu3R0aBU0IUisFeDEnOflHxnhEGRGAKwLxJPq0jmjnkGubGT9ZyHOPvk
LzqOonF3ye6R+Bl4zup7OKE+/ofjzl/Au5YbkfeIhHyL4VH8sYqwPbO8ztmeR9AMteoSw5eNymps
WwfumNG9KUOfygazjhw14tQkdiXgWuzuZL+YGo0xkwbejRNkP+QFj3G2jH1sIrJ13ryDrBlNAjoJ
FRhtZQntiqIQ+5qCKM5Hi2/o6v9QwkOPbousTqrNYmtDJ+XzcZOHqzC5K6K25f3ovigw8cOLH8go
8TNl0dZYpH1qKiyo17T8yQ9WDE54JGUwBnOAj5iEfRxYBRilEqgt9TZbgZiE2Qpu+OJ4nKRSuaVL
DJ+oKk1ENhzvhKzM5+yjroK9pRj2dlf8JQOwCfzMtph5yEGjXfSy4Pkd2yub7ObsHzw9x4HIKeLB
pKF10xgg692QjcGslohXxhatXhqvCCa7t9hS5CYtgmE8xaeBeCYHwaSf5R/MiZR03G/qkaMmJWtz
8hfva5FKYrA6vq15h47kOo426o9adH9qHB1IKCCi5OTZeZ2ffFBOcOF+n63vikWDIpctTRamP8II
vH3cN/1lVJR1w80rlbYV3WyWqVhUK4y1li8rVNFdrFvA4aeWv8+lIgXdvuSFF89X0F5aCaoZxdkm
ZttJGTmKjPzW9MCUJazUuJMglQ5rBoDHTW0Hj4Or4EwUpCRNEpYIaMfQb6xK1PANh26W++/MvyRb
un3g1zoXUL2nU8DekrRA0eApAIYaT5bXzSvtJKZoP69lyuNORobfTqgVdIfbToqRupag4UDbooLn
egTSGdxx/tDxGm+O3ZGvgJGG/Ccp1WfFOFHLF23f/IspszMx83gTa1yuDJ3xrUqRylr9Yxkb1LVf
8zbqohYguaqXoAPPZtq8Uy5AnrJjgvgBIxy6xxwIKJjYjACaOP0kpxVDhIVvnW6GmKUQiAn8a+Lx
Lud4GljrLYqv9trvmMIv9sI9cnX6fAd1cczwREySZvejoby5eLpPmEi7mRtZnOM/Ijs8lTHQJi9k
bh61iggGOIf7ZZXK9eqO7u2dsGe+wlg/a/36WtghePQNrZ3j2RpCFGySvZhgNrsoqxYqcNXxBtkD
uDpNsHg0OzDbC5bS5N/YkkkMa6KZiawkxrwoD2xrxvh+k8jDQ/S21IRLNnN6lBnZcMLr+QWETfFJ
v5Q/rRCxHmde5S63XHHDoVR/4b72KbsaB6s+Kxzj9srbCWE3XUIfEeqEX5SaM6cpckUvvIg4rFDo
or9uZRsNG5dTRPhePYPbuOhl5YIF3vixMbQy/gA+DGqAe4UkXXcufhDHWFsOivKA/wpJ34j/WPvQ
4x72ZjZLDrzRscKdcgcIRfP30WDHddEMhYekprwI7MzEw1ySe9BjDFDstBmoSOApNzep9aWm1NK3
czlIWESPkiSp2M3HMQmQgvyW9xKJkYt/HAb2uKmGCE70cG/wtnt2XBga4CKb+1q3fdYjVqUUk0me
MF32p8COMXkTzrBtPQo3ApNuIe8mJ1BfIYoJLvqt1byJZhNTAENG+3W7+8PL1dg05+KRMR7U4jbF
VUFp/G2XwKD7SmI7A6FjjRdXBrEROJyYUe5+h++j2Ts3tXJP0X94h6RGlxhSi19a2QGuM5xHsMJq
fO0DfARKJsXbiU/P9AO0KgPz2AqdPufWOoXf6itE2jB8tbZxv3siExPwg+M+NU3DjkOwYLwbokqn
pZN3/4DDcZEn+/a2FaQ5UPVkMdQZ3V2ZtCeaJAE1Oa3B3mzjxc5YSKKDMWoj7C7maVtYxOHDJqeo
LO4OJlgIfU4EIAspwotRkJfSyem99KK1emn/2Eic+eTdVUkn3rqwtTSh4AtYDVqL+LQYVWMv+imW
AW4uzdmrpPV7rMkFjz76B10aGLcMmZNc1MDDAzGa23OESl2cM/0eylyjR5vecfkqhah6hd4hCxaU
aoxnclswZLVJIQJekPMs84imEaznqqc/D6dRdnIWhu3mllB23iwm8EO/UhI+uYs/6En8JyD8hHd0
20VGyx8sY4cLXOycI4MFwvmmffqxCB+9UIH1ef2LsOsnSja04ejz56Kay5NGeRTRMSe0GVxs9R+e
l3D7MJ3RrsJOe1dzew5sTT7rziQrqZWLtLyptA7DkQHckCD8pELTBXPGEKaGy/+WEn6cOzSM2lJ4
O4gN1eqnmM/gp2rxGgRnzWg5LqR7ktDT/0R+gCRMFuOfaXQy+19j/ISHTb1fnqjO/v5dIqsUarWT
6UUbibBEWiW8usX7b7E0gRqZzuWHiCbzd81nGn+gXuKCEMNl/y2cQmRdrs3gJVS4XoXtpjDm4VRd
PtoQQJ/ixW6HsZmYViem+lH2fcA+k0IKtewVrDXpYbkumgOZDD5lHLse7H/ki3oose5zYhvpnsrJ
BUeGHc99pZPe0xZNTwA6O+WZb/fkOs10nlO4IWMajIbA2lHvIVeNum4zZBjdqs4AS1Y2HezrXjLG
oKGr7HZjilzkgKikryhzyeu+IfzJZ58JdXrdGqjF0+EpyxSNSI4+fnNNNgxQDLXt/n70hQ/aEzuC
992SQw+BY75KXPP7FNJaqZ7u10hU2vITnNan+k59to+eT5YtTj7z++jx5HCU9D0sAeQOp6DgG97d
nz4VErRJEgfkgMyhlHFZLX+bCQYaX6wllkZQE9UIZ3Vn/+mh/Clh3W02yzjfsSGN1J6oBZHCZc7a
2RBAJo3ZsUhEhTIF6LH9j3RL8zTh0UHAzApx8QrFKSakYt14gWKvDpLcicygVZ2EOyJsWo3ovU0W
bckH12yJFqW7nPrFQCKm/pR4Ubu7hm4b5m/175ksb5Gr3SarkudhwhAVqLSqGxzDskYTRzKfNGZY
O6SXdnhHE4KtXLB6YzWIPkeAczuxTAUYXgaQ6Diw2JuLhII6L2TmPlP+ACT5hVLEflJ3JyqyVYXQ
PjrB77V3NWlTB2c3doWsMCkMLu7E73pfpEDzhwDGo4tOcqX2vS8Z1/nO71ybsPUstv40sT2MIDJA
nLqKXTQDmvuQ0P2KvHXwHJCAO3GgHAN7olXzMtmFhEI3Y2SmSq4IGLYW+Q7kgE4Wn6aUOW19+8M2
aoZu/nayhp00RKRDppqfpaaCjIeXRv2I0FmRCNXP5vNiGCQcc0izs4tnwf9p4lzAzqN/hDqtnfEj
mSyGsO7e2Ueey/47YG+H+2CEflrKe2ofYjYZaJDv9LJI0FmXZ0f6I09+7POes3zeworHVpEZeiEc
f2dJKV52f7Y9WWt3NoiaWGTFbcEDtlFF5ikt6HvZ8yY0fvNKSSTk12MJ8pq1/3hILG5EaI4igDU6
+9kNfz3T4Q0D0CZ+WOg/F0SzDoQNWCh+XHdbNaUfxEz9xCMNq5ou2g+cUSQo9n+cdtnQZ1ocjHNk
UC4CHvO+lPnMDFqAwIYBcnZpuV3MJz2SRjqVIQ2v2iuKa/3U4CEp6W4iVG9Zs/rvY3/d3MhQFnFp
QdTmRCIIjqcCGMYgoL5uy6mYzIfP/OnSpFlxndKfquKINqWSCq94FisQTQ+Wkxg3MSXeWTt2RdYD
RZzVThd8bpJLo+aaDi57TluUFF1I9QfF8SEa32HTqiI9JCWEn/b5loYw6W+mnqEpYIttSWuIpKKn
lET/6dGOp2B5QsIRromO3E1aahuo2igcCMz+KauWVrHh5dzk79k4RSgnqRE06iC64r8dDfhoHSVj
YP3fRNN269nJAgci8snl4/puSrpjPJHxIJCcHlhBGKHXL0adsx7l4zz4B7UZCc/T6MPp5hHJ6vLj
C8BXZBWB6/fwGq62CKdtKzY7P0MiDlbET0qhBs6aiBNuZsxBCt3LF9duca95HxPVrrcDkJtpp2/P
mrQkf2aFaHyWWijoJAh1z7KuQNgc/oBcA/nneoiFGJgbTK2hVJQoGI3R7wU5+LTkSxD+pkae54ra
DOr6iioG8BmSdDjTRKjaaMV20PclMXDowcxffcMvVkdB0Brh0Gux0exwDDiCyhxsU+4OILRZPVKb
h3whehtT1fwW+E2qoceA3JNHyTDGaSrMBpUqfnHrGyldJ7ayq3UElsz4b1CRXoXssnYrpNTp5Q5C
HUmat6fOpxzAPRYCMOLBVr9laU76kjFFRRUC1f1lK19Foc6QZ6gfLNqmncrP7F1vga7qQ7EH6EaJ
x75DpLxeB3L6uIL3u8Tcxsmuuwwh1Dtp0MsAzEERtY5TDDgpE0IkgF+A8NjnpTdjwSvXLX29P+tc
No1CWHqZ0V9QQgYwSkMend3hyJUzDZMj1mTWZvt6PRSIuR5s6Ez80u+jofBNNvxU1egsLCWkD2jD
qOU1hNg+uXXJX7/hxCI92soLcM2PQp35MqgUTXKzhsSGDPEpoo9Ad4U66ZfgSNTdid72K5+5b/7d
sE53RLdjWLyzylpsCqxefI6nyctBHm7ODZmDGJ6S/f201xL2Muefm+2lt7uGvKdZ9Bo9OK70/bY4
nU8ssKzOTLCySD3PcmHpL1QdWl9weVXexXa4g/qizcm9CsbM/1kbGHFXfNvS2tm9Ush7lWpRyo1l
hSUzb+ZpMAFI74ZhQgix80WBCiaMDhQA2ZC5SfLnzmMuFvh9OvQQg288tbW1WYAW4X8P9O/Ufu6q
ehUnR3CdOEpvSMosJKcBfO/6JYnHf15lwzFERX3jzd58rAOcYvQr9Hgrn62gahxo8wrTWoDPcHI0
HWguVvz2nM/h4I+EZun8OE+bTGqT7S0MflNL5QDtouDnBpIigAuqtZiAtHwhpWInDKOwX+mgpzoz
1Qx04VdOJlhzeVCN0lPlZC9vT9J3b0RoO5m1uTZRLWxkwgbC+8eyfwFj/Y3jwZREc0NFXSv3Dpna
pt8MDo5x6sFDsGuoEN2MnS5DzbcVi6RYMV5VLr+7wS1FZWMIcejRRTxLO9xotXmh6bsSeeeY7sa8
/Cz202wqex4a8mSBB1FflrwGmpp6LszBGOaLlopugJLdMaoeJWVbjR1QlvXAZ2lVjMn1biON7EFr
jzZHJY5MaT1CTheRTMgu84tsL1ASUN/Xe4WcMZcF30M6te8F+tnJ/mXUzNTWJBZNUQI6QqpLUfap
ReRsoKXsceUZ5erh6FRJQmt4jGrEMptvy4RLN20yJi4nUGG7jqE1cHzYTogzOiMxY4aYMLFf3PwV
F7x+2SyqN7hi4TsXOoTRIqfDcQ7ETaELLPKGTBbccAThrNZW95rHVUw7GpMs1/ukX4rywcs9jY2q
qPAZ1dTTlilBdNmhy6qUCLbYvQyo2l6OvXFyGFzRFWcMW6YfM9CVLQG0/KKm7ae+E4ToE/cp7txI
qPNJDxirkUhqOEc8TKL8sU78NcRohrJgpmZdhTL29wsanxlmB4Z+c7bNdVqHKtcZ51NuwujN1FdP
2U+oIafxaRq+7lWwqog/pyGKxhY5r6EpSG4E4zaY2XCs3pX6O+vz+Z5/WU6wWIJA197xjI9ZbpCU
Es6FHSF0HclC+SblggnaLFqtocaXJVdoetdTtqZrkFh4QjbGCRT/bx2CU+7thurS1gif9CAcu4+M
PgS4ggMLP0Ihl7Bm5P8noyJdAlu4Fazpuexdhi/v1anK3Td/7DNQRKw/S04Th8+skXdeLgH+shl6
Wn36ZityOwVXGp6ZNy+YgseBYdcwlvcd69F/16NNzHOITbi4b93r27DujfJ4HGVK8dcUd6EWergT
WpeSJ95I+lOfzMl2P0zd+O4dYjqysXW4NH25YCNeFTsKvejzCGXWNny+/hnf3fB6U4ZU69BgWr3j
yuN+UpbcKXxnNe73OXwSUF6VBPNZZJS+i/NN2ZLrTKkSElXwUsz5d1hQG/4VIR84rW2ASL81osEq
vFjGNZClplUtPn0EKu2B5Vi3fMxkqOa7dzb11OfRQJ5FFoISo69B1NVIy0QnUOTteDBTvxge3GGr
ihaYiE9GN23TyxpEStWsSP2JFa6miMtdaKg7rO/f6guUUGqnN2HQal8fjX2IvYO+8nf6bkdATgWb
f773vDBKiK1XFnc1Lc/2LvCPzDihTEUtrzGIWfd4DeBvDt0UJK7lbxeg2JWuK2iqYYO4QRgTaR7U
jizGampt4gMYM+w0X/iW4Jok+Ea+VNjh07uIqkkBNKfIQW97sL/6AWdUdxW1ugiqX4LY9MsYLbh6
cqNb8KK/DJgGV549SS+4vusiHGC7Lts4+NeNC0DJZVtG1iC1Zs17kXucW+Y62D+yLdmVcGOPT+N8
jA1HfWGRcIozpm46Jebk8CsOKEUTtRgI0JxfRZ4SthH9m2irMeBRiZFONAAiDTZRKpRzVxgwgji1
z6MizXlpotwfDQPyJ+0BVqBLHNa9n2GEC6XQ+TgRJVCGEKB20/g0E589QFLaxZzTqcJa757JlqkF
iFNvCNNoLeTb+SVxQZNnX6YWzo4GNQaWEERPSbcdN8cszZlVhoC2CeRC2rX+YUGKaJK9KTDiWty8
VvHY76bQHaooW3DPnzPoyubIrJNDSKiJIUXIZFL0z3xemlJLg0RYciwoAqNsOqhFlGkyurHRj/5O
yog3p0tdDS0aPH6J7azeWjGAy1dQsSOyYHHhu+n71G/Tgiwunsd3fmO4i/PYuL51NwJgb3gS7o3N
KtsSzTWKrGjtP53LHwipjrHP1JD2B7Vpg3vt38QEF0EsHo2PwQG8gH/iIeQq3Gg2plD8hrEbRbM+
47WF6YITSkCJ+jTyfhEu+FN/xYtCnFfgHjcPk+v1QTyq43SfyPD8u9PYOe1JejuQ+h+m3NJ1KPz3
dsx5HNtPsWP9ww9CLU/ljwCDhUgbMGAxvFEwYAWI9nvVcnpRo3pGr5BhoTlohZEnPA3dybI0DAaH
2txf10pinTG6ZRgsYf51xB95t2Vd8sVTrpMBGWjn2DAqdg/JtnMA/iBGvkiop48sGq0kdd7rQftY
9yh0TKYrIvox5ZaDjdy+8MgbpXx2GFcqwy/pLRr3EWfBLAoSsWdg76M6Qq3kQ7Je38TbMpw4x7Wk
63bDKdkQXRtOGRN2ofWTx53YqHPb2Q5OHXdEwSKztM4HltN9N5YDHGJTR9DvRnC6KOT2idAHX1Oj
M0xywwqVB8kTD73vDOGPcVAz0oxXJRRJ7X30nfA6F4PiBinNfOa1KojxzN1fg0f5DBPzsm+WwZKQ
j2U2VFSorRYCgCJy7q3rVV7j4hVf8bDe7lv597n283jGDNOZ4cLtpYKkVPqwEhhI2cU3Z7R06+Dm
FMr2PG2l9SYyCXXG7YPvr5IjXTLdyC3taD9jXyoFKKgE6/SKc01gjlIL1v9HoBr5//TykWvH/vFg
NsTnzQMDtd2l7DNDJyJI9bZ4oq5XzXR+umBjVK9fc9dIQX5VV+sxqLK0jxsfL3kehXoHvjrdA2DH
Ims2l6bEJFuHZdjO/93xKN7eEUMzHhqrGPhy2vg4/py+I2gNMpK3NXhOEEpND7UbydUqhggqwaCj
ULGc+q38hf6t5hj4dHT9Plp5D8L784Y/KU2XZ8B7fG3gFdVAs6GmLuTnW91028dbG6xYxyKTOefs
KDJXL8R2eRA4xX0uoFZNPpOeOEL3zip0R32Hvust/rnS9YGLL2iy4hY2qUB3VtiBX+2df31bUH0S
M5DijRhfY54zPD4/nCLBLGLnDp65UW0DkI1Dfv5iyq9y6CxmdYhFdgJ12BycCAxle2RKDQvTiEJ7
QBY1Vp0QXBt5s5rj59es7z8vkjPXj+ChtD+bLkwnmwA3i+Yv+IfQJSfGlABa1Kw/fscJnNan07QY
6EZutg6BSn689FXW5ZWzAjKlWlWfjIMxDTV6Izojs3yfRxOZaUwdgVoSh/NpwZ2lh6tEjgFwUiSi
S/DItPVa2hcUb8DWHuOtG513ZYPvn0QT41n+uzsvwQ65AlHcJOrNWwqyAynktbjow6lbOrBqyYSp
WKile5eGnTWZaFUN24SOGwWugJZVPT0aEnPEQFlXoo5vZOIGg/mmI1OL5zgvxWuZ8lpaKz+G3R6O
ejHMp8A88/gMJXAUIFvTK0kMKGEdHzILxxaH774jC6ZsUgVx62BSM4DiXhRoxC37wdMf/6RSYCPr
UpW8iYmsX4lCo9Lv/hebUwaroLOYnZK/IOiNr6WilLK1KG4OooZ1W6BIozZ7jZnbDz2P0qnbZxk7
GBE/eeXpzB17+IaFv3N3cXV96Q2hV4cBVs4WuPLZN+pwQ+r1/mstzcdHpGzAYA9i2YHidK64q9iS
a2cgk+ijNblwA+pAiZl4MV+zYgEdhSvXmpCaQ8dWMytr4mgKelg7j3Za0HpcHhTcuaYf/Dq8DbjR
iUXApXBngxBLKSD2bs0oRa3XqBzSW2hzDijTl3vi3krMI8M88ltkbLPxJdeRioBRj7A31qk/yb7U
NDIGj9Yxu4TODTqGPAFYtyWUsJdrklBzVlRsU0rb34J99miXn4Fbt2Dv6lTod2/H/FEDOmPKD01M
JqVHvv61FYc/WD1d587WG6LHD/4nmDLeEHiguXEy7lyH2IbOKOdzrVKwoB7jBwEtukdBYqq/BFB5
1RqJmjK73vjk1ZJI2FLbsIrnR1hOc02Tq0fdolGK/rDXMSzTgkQvt3sHXSz16dgWtGysKi0yK/DK
U9SrZNGREVT8b7KyeolvB8/bTJfmO+ogpOE02FtZS0Zlhvev/4EldKYHNwzT2O6PJRMxiy9U6nom
8JRX+Mkf5fuW9xZEvjlv/ZxsLEsPU1zMbq2RU5V+HjgiElhwvBB6QyNlFNyaVzx2K7r25WDdMOP0
vtLuLiG/4L6sCsVC3eHgfHB3t3jn90FsUYDwq3RYPRlYXcpp6UUoCEmAt0Xl5wxHu5sqVqNXJQfg
GetiYzTY+r61wi/ISdAnOKNWKoNb4oNb7tpg9681lLlFhUJcdoimKw+P538PsEO2m0JZOfLf73tg
oMS4OereDckoqOgvav8t8JcVwiOYHNpYDo9C/AhtkXH4rAUdfTlm8zlEO2y7dyCr9ot7QS9cQEIK
TH/VHHH2jiqPSdVFbvCLwpHrpV/v06E88iT2ZxCtCUV2TjTtx32IqWTQcmgQRtEY/7QXfrBnMoxp
ObOL0P5XheKtTgfXQ4aTp5/ObaNlglUWJr/UrlTueM/MIORb43Z6RfQKonx8FBBxfvW3vHtl8UGq
TkNQWNXZXk6ccj9GkNPv7r9hfQPgQ/imr0r9NSLCIwF+mckG/mZn/VMUM0eLh8+hbjEiQVw1mF4h
3d/i07uhzehybUwC9qL7Ks5PBFMO72Jk8d1ZBU1sFNR4nc/XaWFXZlVLg0z0DTeII72eJpACsP6R
WTKEEl+BB2zBqSg8QVaqpvxix7XVaZ+36FVJquLuf3hB5qpxAxrRbm1hv3uXPJ8gc+d/fChgDEIC
ZtFF/DU0KfSa3aJm3Dcc2pcQSJE9ygTAPFvlwZkXgTx0RIZmJvW4fifFdx2WJjhE+7qwNTtoN1q9
XOxUktccMgostDN8x8XA/OqAHt06DWg/kJpA5qlEyXeMjAu0rUFHjhQaK1V/u7ImPS5dyueHpgKt
nPRDRq7cpjVtfndvKWT+KY0gLyRAYYZXpt7oZCqotJ2u84vL5U4lsSkOEGxgkWUipziaWKQwfJV3
D0ljND1Ghx/OPagur0EAuwN9M5yqE0GWFO8tWnoH7WjE6CiwOmD0uU9Km1ufK/pp24Lw7ovyH1eN
icnfcXNHGpyI1wydwxWKD1JErAjOKvg6xaMtKIEehwmPy4YYOERokOtJUpAbHovI5RLFGgV2g+Ad
VxBJJzo8qT2vvurvUiyMQFoAkVw89J9Ps5NbGd0zpnQyWM4FVx6v3b2c8xvhd4Q3i2IsBS4V8Op2
M3VPe4EC8Qr5y9F+gjOjVpbv2CQBy2I+jJXoMpZOPb8rR3kzaZ9Z1ZPX760QxiMwrTFhCMoNs/2s
lFb4B7U/h18hWei4p+srb9nhtioCa47apccEwUIdtcq8yqRmLfLGbzBb901BVBWrnEo6XeAbyK7Y
Dxrh/8NX57mL/AoUyAKeTcoQvvDLDWR+phI5xbKf9eX4VKLXZlpAhkSe2wYmn/cJWg3MtYTrjM0u
IPWYKJLbCPJzwjqsEDc4HaPFJrrB27A/UKX42LVUsZGzD/9lZ4+wo9NnBOdUHuMwr/9JyUhNNYwl
MzMtbB/icsDt8KAxdQPYspEjdDfWmZdA+NxSq4nb/xfs4eJsbaJow8bVICFXtC55ebyl2Dz0DgWs
s+W9opcH6Jg2v9w1EAtZLgrinuEwzqdFelwJXBzjPkk5Mlc0rBOxOk6/lWmlwrCoMjPJdwkRZUJ8
qSZctIY740N1MrGCVKU5SX8ADvfte7fYcdk/jCRV1/P9gxu7hsGJmIYktAfkF/UcXjS7IqJwk71Y
zDQR11bV9CwZOPKTQROSKMQqXXLiwy/4fSo0po+tqt3dZO+0Ol60JK8ETK9kYChOMFVDWonfBlWR
ifL12+ZTuSPUERpOi+L/hO0BuPLxvHafimcDA4MkVK0uOe+jAuzxBYXc7wnSY/jmjx4CSO+Up0zW
fZchBUM9TYDCsxZvODvyJAgPR/plf8bQ4pThz0u/sBrN/ceDGkNXbawCw6LQV/zcjExhPnDHdT3G
G3dROdGsQGvo4ic+cdi1VRHz9iaWgOTVVmytm82XVH6nCAZnsTucyd+U4A/3rp0qZHmAbkE9qNIF
YR5S5MFpllBz2Gn/6lclDqPGommQnClRaePadULKJ5zmtqb84QJzZj0qlJM2357HXDSj6kD29Q4y
qT5Dg7Fp7/kdRks3hdtjmu1TpZK6kvEIjSpqlbr27iJ5O+7Iil3sku4HYuFN1IDh0fjSCCgLVz/N
zJ1TQY5shXc3R/uUpJFIAsZdspps8OONsPcl2m8Q7pIjuvp3jj06RKWHTZpfiZkGsKUnNBm5ocwa
Ivioww2z+nXnedyJbWGUFh8JCs1aGroztkxNgMV8xAPokHCbHAGx9ZJRMMH2nKpUhKnP6gSXzr0i
pUvy/i3h/Hx4PwnxEJTKFY+VkOJo3EIESI7VAKYNVRmqm7R6zDjas6FX18u0ZFYfVhRxodeK2cFb
4qQLHqDbB6rqqbEXVbUNOfO/f/pF4Tk2EzspCGfdDXJi5z/yGK8Z8ICt4xtWL95PlMB6vNSdDLhX
SZeJv+TsGNnbfKQ+nydjs0TBGDivgswzFXKythCv2TbrzQNt/O3/yEUnqcrbmR18MkJp+iXlR3iP
P9+h3jxObJ7aamsDZnAuO1aDfx7v8gjrSc+bDQyG/lRZGR8KDzUdtQfU3IQeGeE5NWedJdGm/SL8
rSW64OEJ+IY4WHTJ1XmiDRw2hKe3IaAP4vJDWITD1+MWoX4BGG9+CYr0NULqWlyyTyMVpndYNVin
bqtiABdk6b1jX0a3i1bLdQWslSKRx6C5CO4RD8sswlINpZxaf6IYf5ME9AeeWMZjJaSgFHjLH9vz
o9yFoy/n54Z1PiHdpSVt45JDYXuZKXDX9UgXmQfPdIuUAEkN2M9nJSeLXYiuaoLFqjN4Z8sevpxl
p1WJe0qadNSkygSPcoWylNVO+wO088z+EBDOFg2bf1C4F9SumR+f5zB0UWQqqmuOCgUeOs8nwEFa
4mG4a07CxWdBJIQu49tX5474bB/EFfHjuHf6DvqqoyE/LedzOf6OwMxRbgdf5gaqo01LJ3N/sZ+T
ToI7TxzLp2cFDPnSovVa3QVHHJxgfkvElHw74EUzvPyoxUoEJrIb0IhNGbu8ial9+qOOOKrDAUTt
GW2rbY/JTRV1RIre5MgxvA4WT+/JcFNdga1lxTu48iv3vQihUYpCy7lF3YkT0ytuuFjHiEbCZ212
10ZoMVpW8k0igPJUPvnUcbRAXqNziW4JcylcsO72HT5lTeZ3jmLOy/anqDF5/YdiztAY10Kfiu7n
+VQppjMq0NlZujW3nVSWiWRNnMyohRsDPYT1yku26LK0ElQGenZLoctmfOk4muC4+QXBQofWImzO
G0akhJCai/cxXdtMgwY9/+tQyQ4Qf001IfyUy/2ZmAU1sNgd8safh2ONlqSXvisl9BNgdCtk7UIt
dejH7XzcBFWg8uGS4o6kqQWkosmXhJSciXSniq2hSqjPb382amR5XSsTI9mPKFwjQ0ps014GQKTi
M1N/bTAWgheVAm/3xd0ZDJsgWM37HIz56cAQ8lPGx80Zz0+XEzKKBDe4/oORvAgxzMt0kOntghjY
Kur8ZyLrXYqKRZC07fT7nq5A8EHIiHIIWRE2aasVUZ5OqwcDcKdDgR9WT7W+R2/p2I4qPlD4cxDU
GCOGozbWIP9pHUlxUprcdZDDhUxwO6Ee5iwpfowvwea5e+QjuMHpKmULZm4JnPyDtCDhdBXWw9t0
iVex4DtfzU0SBRm8tcFl3I5ljDJMb9b5hH5q9VOt2844AP4Lf57NcY6TqQLNFRQ1kbEwEjVkiFBN
AqUnUax5/MKmtJOMrer5kWW4O/NeRS4UcMLDxb2u7vFBWV/z1MZBu481i5Cf4V1lR5qr1WQdh23t
8wfTgNM6iXtvXZMqqrTUJfI+0P1rW2yz3ubuDrVWNpIizsILoVVZe7qZLUceJ1S4U87hgugrgUFO
Ko74mTBhxM0fTXh8bFa72OGKc4Q6YkmAv5x3z0XV/xQCQV1yqe8FYAqHGnQ3d/Y4NOvR5rGca+Tc
KsJgchVG6mCHrAiZYmGhUGmsw01Wn+A3Ch5Wm0OAELOponH8AqdfNUgCANuZotGsFfH/LzA908j9
mXssxEZuBUHglOBU3kURYogD03xBthTz2P/9QgvM/fi/zhX7KwDJyqj0mktf43NKgQq5TCQm3DSm
87hW+S+OQBDZFz3zlt/lO1JrkIc9GqssH0VC+ag9jT1eGSRb4NOCZJliVlL6rRB4U5oRRcqFsY/D
tPTFGgdWzNmIW2tjRJgB6MNXuTb2DUKpAuSmk8b54McIZS5Bp7q9Ti4Peo036+0ei+J9V3Zk+lbr
DjMEQF0/xcrYcKv17TmoNfSpyaH5xT+tYRFMcKQe12VqFdwpgeNz3U9gjZmfrhnKQfGuVsr+tGYE
1QBeeG321cTu5mA5CPYfe1RXWeAGuMNc06pCQH2UYnBDk9aiQ+BjCXVlOmsFHTAiay3wqoDjx1f2
QjtburWFCp8mG5+kwKVbHV/s7pC8OcTy6WsoB1zeeh/P8IXa+jaDldkHUPkVV5wnTGdLs/X1oRk1
a2gx+SfBJ7hW1JZPx937ZN5DjMC/bIF4DoEFANP+8B/ITRDMIWYTdq3u8biZ+TZTUKqboCBNy9HT
X2JyKHvocxytH1NTvDvYxGZx11OEJxGqfuSNeL8EF4k1HVNaBv52F6zfU6AZ8WHEnF+SRrcYheRR
Z8AXR/xd+xFayFtyexJS+Iu+NktdLRMDmQ/OWVFVbYqD4eZ4+ie/JcDJhqCC8O8+5zOqghHNV6K4
MfIcoPLlMsiX95O18aF8n7RkhO72IF9+gm9bLxFHZc764N5iEKYIoPUE9tafWaonyctPDaQTnEAe
LS4gYQSwsaiWPz4HxfPYPSw1M4YIQTerj2EooTYbcPHGmcJ3/e/uTGy4NgdafDb7x+syH8YYKuvi
Osnda+FdT0iPn6zU4gvc2Ft5O4SMYF8bNsx82w5QXbSWcZvDp/R7AChPIZEzqJpt1DL/zplplXiU
rPo0KpwEqp5JWzeAo/P0LcM2oM4CAYU43RUdaYT4mH48/NM1+IHwO1gW9tZ8Y+wX+WGJVczWL5YF
Q183BHBRT3NBUfIP8uYSzujeWVBJ9aqiU5UoP2wL8jFX10ufHJTpzgM6hKGt6oJffhzZvqWxrQ1x
WE+dKTmRY/oS+lpSqL//r4Lm5Wnj4YFwF2ZvWeqlPIwgQgDHpNqxvd0DINLFrSfP5IRDguc68R2r
6mzxf293DAGrWESCKi2g8dKkQ94i5svsxty6CFqmCeJ7BBjsVwitG/dZ/XoacKXUym+7+huldalQ
wCnh3wJZtzuCdbw/wNEOwu9MHvWrDP2slo6i1EkkUOI0Mh4dthtGDax2KKxRx/Sk53GcVXiH/VFY
q0On2DBjAd5iCFcQT6zhfmDIcRyT1O6h/uNycSV4IpUbuB/Cfrk5mS+3kn6W78Pl9UwJW8bM8Rwl
/+rLeuwbrRncno5Gm1knoD1ZiSnheQxZu/hcW4UwbiYw8yG1ffW9iIt0Ej+JSmDVNxZkJ+HZyzJV
GrBe4ovHLbcE5vu/1SoYNvDMxCJeWWgOkef2dwuvRs55hTClNeG4k5Jl7iHLSIx+R8LRwnpGf8fJ
ZDFe58c4JyFSCh9cg3GtbtH5Jr2aCxMK0dcQSygm4CbBucbL7aMJ/F+Oxfz6eLi+vt1uSbksFjHA
wdv7LfCYXFmJuhSIm7mKWEyZBZ1ZOa0jfH1hH4pja55l02leEpN7Bfm0V7AeYgKYZUTWV9/o8Vh5
/maaHLPsMRubzl/V9pBcz/4Iqjy+3sb/VOSF4IlydgNxwh0gECKuIxFUHWJKkSY67fvLhddmeUPK
b6Ifjh51IWKB36ZA/8O4FLZx28XjXU4M4CvzejL0vuVx2UxyGw5CdI6+s36MA4f9aG3ou/Rzwl1e
B9WaFKzKchC1Nv6f9OsggPcLrr0G7QoxiVlD86eGAmZa4IgHZ4M64HYxp9tEyTU/+MJh5HhtO3dw
fHOFiNfXlaiXzd0W5oVqI1VZvWacKC89+rrvBrYBYpdM36exvote2l/HBlWuGmGuw0jKahFDeS/p
47PhFQS3yc+6DUhIffyplrnmBsbdcuCCwZb5db5noNWG7QZi3xbWKpDH8L18CKj7xQR4OkTHGa74
Tng/H7d3w88oV797POh+C5uCs4eumFrV52p1sxV410uI/JXvqQZBYO66Z5Gb8i6UIUBok/6St97m
K3kwOvogOj8zW1yIdCJOJs3sEX3y1KVdnlQxkc/USVhdfnyLP++R5OQdfEdxKZes8Pj/VAdSvuMv
rNLOmLAbGAjEoVSvfAM9M4UHVGx8E5TnjR/WsRDK/Jt4MeXYKdXb/EYLRJqYMXNWXzrDrr1OY0hB
YZpD8di1OELwcbr/ktQxo1B9j+FmCVQqU1L/+Z2tbLVsCKtAYoosAkP8WzGIQRvVPq6YH+0lwZBp
7a3J/ECWIFXCM5OoXw5aXaaCKiReHmUi5ebvYLRqjmdD0MztgBDTR8T1QcHnlco16kG3XVAbWQ17
cm1fraacssZhjjLuACLiRaldHSSr0OoG+iS/966UWUQI/RWYJqh9exHYjxnBTxF+nO3tBPKeFpz3
WfYCJN7ltP1/hR5QCxV7O3HZZX4elMSjWk2V6MF/96wWUMiYn29EB+zN1PWxQ/OpbMC8t+z0bGrm
0HcwT6OKXwv7/PTlzvZkZvAGp+v+pK1YTQD2U11aYIStAV6MAyqDeKhqT6bP31kQRBrSh1mInBho
5OwlPGamqHEuKGrKAq1j9pAcf6PzQhSMM9pR5WhH9nmxT7SkKtGrhNMEkIdrzOlXPXgkeQ5v/hyk
0vAKDLyVoXDFmlB3UaNB35Alm7UpvAHy4iVKgX8TbaVOaw8ykq0amn5034IvBZV4xQyC1e5qpq+J
qonmjLggnsEBGbdR5C8G61S1SjVEnPcLu8tTYILiBEu/C7Uu7EaXJvaYCCCYX63w0at5lbOo3En+
CA7oQGkWuPlUqGHPZEV4DoftTuxlVVlkVdA+bhKoBaOVoEHQU5+G0klj8PjeykqWlUFLNE1VnI2i
GOq5DC0UjMDbS80V95JE/WOeaZSgQfERobwwsH+7sw90dcY00BYP0LtEARkSV0RK4iVEKquIOJ0q
zPC4yw83zjZL6omgAqVnO7JM+8RFPhJOB0mBDxX/wK5BVbHmZza8S+vxKDZitd9n2/7WRAHe/sqm
i9Q3jZvQbMqWYHi2Azz1I0i/3hvIwGDEFMMz/ob5W61YDzy8I7prRSUC5Q0i3CcFllM0mjz0CgHp
NXy5oAf55KXt0AVDwQ4HNuiBtqQ8fxzz6g+C/c9+XOmFMJnDaxMVs5Co7iiMcQ3L7vIYqIiVQC8/
knyPENNZ/s2pxAI4W6nx9dJFx4oNQp0yyUCliLtrjptNsuIcJbozqC8+ehbwCG3zdBXUw+vT9J1Z
4b4865j7lfoagAM+zbnlIOQFqvDDSDrQ0A9/wl/cPbDiKsr2n2Icqi+kMk6I//TJ41vc+GQFKYUS
L0yp+PytTqj6xY1k5Prne17yP9/oj0gYE3uSrOO3BHibvEI52DBYOZFaoQjJc9QShFJxBNG5kTQ/
pdkxjJwl57PHpmBdUQ8MufogVh6/GsxAKnT6uD4pltD/1qqTPjUWySUf+0gKFQ308y0etw0bkn24
U7lcb44TZUJZrJae47EE5oeTk4KAMsOFK1e6pSocJCKEKSYcDQ8iPkMlioInoPXTV8xe0WQ1EPE5
GkgIOZTTPLA3FiUtSWyo4defIHbUpcEL3ApzP1PKQyt5TNjZmYnFVGohmnA6ka7ndzGIKScPNt3z
Ztd5wPZ0O7FVRQamY9GOt/Enp8koyv9jvScDeHcrr8Y/Hmjo9cB7gPkuGH4feWr29d7AOuyboXjI
VEGUUfCPz6jyhOcetuOtsqMVfyr46CbPVka3n1FWu42ZaYleh4lzQbXUEIAcnPGFhuOETeUxMnfM
g0pwklBeP5TXIx/IibkqLLxfR4zUoLU0/eSaxeSQu11dH6yheB6pLLHO05//qfQOI3iMPrL6o+e1
kcftfpC0pJofXArsBkggWmmIVhoZxfPZ4/cYxNn3AMQvfZarr0KhbRFfNgZT1Aa7WKFGODFZbb6s
t+r+8rQgzxwW2+s0lufSIO5sixRrTVjqSN0VRizN/2ZQ7+sNwqCMgmVCspCYFc+r8/fORWiY+fDK
3p33UbQ3N0KcjW6wltCDx2T4iD1tVVYQ+teZhF/DlSXHEEiqnOc+9gaLfDyZPBpiZbNe2p71XvAk
/+EhJQeUOvwHxVC872V/j+nZ+/bgVl/6DXab6hCCa1v1OmFPkYJNmEr7m7pSP9Emy/9ib2HPlCXg
oM9sMgkPAlgT+wzgaBQySd70N+ju+wmF0GbOB+MLJooiSdQLsd3jgjXmXm8VQGiIokoCJ9ghq9Ia
8miKY1KHhBUhAB/Y2ORTgRlZqaEA0vSrASRK7SDTUNqOW6ZAYADSa6gUYugqZTrr/ZY0shIv388Y
WR2SKbBzuqxdPBnxC4rUv6jmcY/a8bPQcEv6rtRRNDR9YNEoa+Z5a/I20mzUddWkGBl+golEIzyu
Wd5uoXEDOwYN/B4OgwFrEPYWmZWb+jpVdAWATJPPOvKWFrzEoA/xwDLmABFKysjHb73IoY2txUml
1pZVOYyULVk5JaKpOmA7O03keM6JRtdajs+dd3aEnUWIGFJZQeboLcU3frcZab+UUhMEYZ5a0GQx
WYetK4txP1v/MDmQu51H29aB7RmH7GHy0dQI2MGbRvrpAJ2kxMSYcAif6UM07r5mPA1h+mr6yQNz
gwmKBl2H/lyin73mlxPMn1tkb7fMon+GxtJO3XVBRrTJQcVjXe/Tc05DtmzLJoBeq2LMcdQQOMAp
i5+B2QCw3oNJzjnNkFsELgk4W3VSHcNbPsi1mf5T3y7psFY+inHgk2aoB4OZUdkIXM/CUaIbqt5p
chLBGzNAVzsBX5sGxtbnocVeaHc3Mf6fELDYTjz6JfzRNNx1ZgfPvJPjUyBR6XjkWKuu9bmoeOlx
Ozw0Y2qc00qofp26eDrrMTWXNw1rVVkpx5Frhz71huUQiWIDcps5kNNH9pS6QDRrk5bJZLL7P4n2
XFH3UyJQMMH0Og+QkbEo0GogBAlbm0KWEBhCdpujDqEloXLr5oJAOKuo7OsqAbg7BsVuY6WmD2pC
eR7wjYLqjeznhM24ibvGqoMDYM+WaU2lF/j0d8sICUFzOAl/o1RqF3FkaJTHBlQNooQKJNK1uQ/g
ajTDkIAFaqX6LgKwbjUXcyIXnvnr1Jovcq/sRizl2tKGrcM5jEVwaHi2ZtCow21TrtVsPYL/xF54
qOs1oV0TxKYYoisVmL0URkyfjb47Q7gPMU8X1jPW0cAc2KnzzVUdWE35dUZe7KsIU4EwmXyFVJFN
Ob1l+zwsQ5iX0f8IdF9Hg8ZQ0fdgciZ7eRLBvbys4HT9uk2bNegapz66jJX/TZMVCP+vcf+ju/tr
+RJGtFQedUdQE07CuqG9wL6VebLbd7Ncjrb/q6DXg9pM7t49kF93wa3WTY9AbXIAr01BLPRQi8em
Qx0Y/tHhNTTpERqipbWGshLyRaUp5JamyS4C2o2AGIG/BKJmOhCjw+V60LzGee0Jhb2e01LT9NHj
PnCaGOmE3QRkCaCwawn3ZnGPcGLIipi92B36AEmP3P9VLApNk59HxmRurBwVWU3g89u6/h8cSBgS
ipGwdphQGZdu4a4v5wtliAaRqKCGmQF/fs3wQumovxba6XFwfvTVQ4ISKyB6aZ0cnv6kUETz7jFd
Kk5Z1wQ1xlu8m8RudoEiqMLQenamzvW+Nhmo+ttvFzINoghqs0nUaRSmbJwuliIHH5tjjWiKxA7K
bVjfhMlTSI9CtAKLA56g5CH/ehAkGccYHZA7D6E2FWNEVR2Ue665WDelGrBa/CqSGlXuLvJQr2c4
5oEXGMk/860c9+EAfJpqdk/DEY68IlPnPcoLTbHkN8FGE0CjOpp7RR/sB4ecWvY15OFWXwRC4YcX
6PX3zOwpTaUcqk0hTUsxbLQrXu1H9Qo5rorSiYngioes7NPfCanU5YUjiNz8SzoNb5k4saVGAKlv
9jmGkr2ERBKs4MdhnquLg3Cl0aH5wX88rGl4YkzMgPEqRFwcA0b0d2+pdulWCbUZ/vhzLhkU54BV
udyuYVUZN8gmyUXVaSam38RIqhpfLA274lLwk2XMW+PTFhDrPzXoa7rBcOmq77iiQcRqQfCQGuU1
Nvvsu51mcMpQRbMnwuGFeNQiOVId7Qjmow+KDIZQg79fjI625kLcwQtAh71pLKyByjd+TSv7ZW6+
rs5mLdzFXerwaHCJd2b0oyvsKQMIK2Vf8Q/sXRmFD6nRaoBXBfGq1IJ8WS1/92PVX8V1ozgdJCmF
KJkD357zmNGkvUkHSPrbr2RmfCvW2YUIhxo75olvzu+hB98wdFUp/V0+XzYx1OJDCsKoHxntyLx/
2YHOYz1ZMi8BY8eRexlQ+HzM4Smk/nU7jr5TIbOFRGpILekGKdDCDA3oF97j7PxB2SRbjAquO4h+
PLrw3m4IvHzbRHznmwZAWETYZCfolOIEbofNHp6Fm8o8ZQ9eYtURDxz593cZMbR1Tf5sJSfZFLOk
sAl6tAQ7btmsTNnavdgcuY5MFNTIg+jkhW0RbnPLYxqTqLJf8XaZpEyb+y3FMxEUX9INuE9IrnxG
0AwdsVWzXk7dSioX3s8qt+Fu4aVXYiiQsuic0Udr2P9LvtjwD0Hk/jEVgisNmFfqNiPsZRUGZYWr
piVr3IcVhWgCspJM/5SJiB8pFH6i57oahOC3mr6daC32dvxJ8FM1wio38i/abDwDoD3ThONC43qG
BbrNg1rIcMOeB4NufllsxlfsjsMZVPExSxProll4kr103V3BeTPBio7YU2rcdYFChavMi0JqGbUP
Le20aEXnp/5SndPW+A/NAD6L+6uvH5drMEGTzpwjaniUJeDSjgQOjkhHq2xjHeM2hrjSRwSutRRp
yN2AIDji7mPF5K1JrIc7hj1CippDxQWZeVqMTBFRb7PEI/bKaEt9fqI/PP4mHLkvnnKwS2Ic+TvE
SMhj1zJeEftoeJeK1xPNcWiPMScDLyedu2KydzszHGHm+jZOySvHABROesosxHepwSdTzEoYmktl
tTWVjZrCmoo4eH3gNpadNfZpL854mS+9T8ip8Od99NBvEads4kXNkWNLiDO540iAUDnYpYBCxMc4
d3Q7EllWhbNd6FvrD8EYwZwUkEwFmxg7vNqs93yJgy87/flbFrA/dwbTv2IkplYnl1o7cyHy4H8Q
hR18u05ixTWEpKOslAcePUSXYrcHI+byIm/t74HT3uwTlJAM7tZ85LSYiGbr2UVzJcHkK/MPwdxw
VHLjbdOax4DEJz8nXm9yWrGfsigkc8mTVNze1IKTPWlp7Eh3oY269fYBLEq8aInCbz0kvtkoFEsq
Fw+HXOn3cXClSITKcdq6p+X6Iwp7KlpSq8plTVEBtU8hCfL1mlB4gyVpBsYTA9Rt45sJpLOiRMU5
Vc3ygi+upPWU8q3OhvPB2yV1WRMjB4u1Y8/OfXTcYyJl4o/YlYHzbxDH4n0Ot1+bDLvst4qg57Ak
4vbEN+x3CKU6S2SZdcrDSNekYCRF+7/4F2gBT+hsXXYGkG4qc6+/RgzRhPWu5XIXLRtIflP7UDcj
QCbZTcDfCd87ezATnbYd9idZFcG4N6y2QWYeDa0fygApcjEwbQpu+/HwckWfgiaNpIIw8cPwXmCw
G5vNTAn8kvD55l9STWwxFooUN3HdNQJgbv02VY+rYMHTwHMBeX086SifngxUJWJpuZCvicySqiY0
Eu7p6A6J/kbVN5EXu/pzQfUcAK1j3VZVMTQ+9LWf4isTN4ypQladGdYVrSaR8vQeagk+Z8UPPWpD
2TLQTTW6RCN5wSkT9Pez5ZG7U4T8vHhhUn2GFRE3CjN2dwwttpeEGfojp3xS1gsK+ljcIMNHysEB
Kn1Es3D1ABwbiJfP8ws8VkeQl0bkqmi1Kfq6hSiXVUfQXXPA8Q2ExxE2iTH+gCa2oAfKlsuOwU0F
IQiIghOfsyGKzVQdyJhnu0V3anQhJ/BqzzWmzDLcR81GkKLADUnmuwrP81tkakhbrNaauj6BDHEQ
xkyxreLeLju/mDPws8kle61LDfvVAbpbL4a6RxheUsLfcGTwhq82b6fONYfJE6UN48TbJyUtkbLL
tRz9kBEZeF1vzoYKOge64hPIiyRpspb9UAqpRaP/GOkq49kWgZpU25V82g3VMCxXr7xHOB2j29+3
i8pTdDmt2wK80/sOE9VccYZ1Su2x10f5wb/bLA0S1F3Va6L6CwiFLze01TDHbRE+Mw09/2/kKxP9
y324aofQqxhUbleJRufrguIKcE1AB+WuGFXYP2sM90xzdznOHmwyXEzmGFbr3/JvveWBQQF/bjtL
I/34BTn8CtkM0+JzaZrY7W6XhKxgqHVgQDFd2p4Vd9ZG0z0/KBG0w+JvCHhgnQYKnlXafrYTQwgh
N4YgDcVgLgewa74jF58ThFizvgQfPIJv0atB8wq3tnkm/LkQAl7vyCF11ENZX77zglaiLoWetXOH
o3eNltC+GNmmuPUEDGhi8BcRvi7NnO6flmgj6pA0U0h4xD3HAzEe6B3/lQC4cD9IIzR/xygF0Bcw
mOvuijPxE+XhOWgh2wsLEpj9HlvkIBVr/d2xznY7n4BIH3/EJH/ZKwWXKmauQdrqLVDjlRQM5fD9
C9zQemScOkQ5gOYPcrw+HcLhlLLH1dQ+wehdoNtDMzG+DYZy8abj1LPfkuxFzZxdwMP0R3Eua6GP
JZRh+yw6+QQ+3mfYbxR2STmyIwbALOGckSOB8VxeQIVQAZ4pwdCS5kNEcHj6KDTOuXKY3Kc5pHCz
8YcVicDqGsh0B/+5GX70lMaw07n0F2cZOGfTEHIPlOoCg10te59dlEjlPQRxaIKkDlfFjMe3g2AZ
osmkVHSMnRTIS8nxCyP9/8PAp6HhK2mahaGFxbbRL2K8A0lBPek05syX0RBgE6FMv1EgyWEB9Ztm
tg6Jv8pOBcTFFSqzFkCl8jlfJRtSazQzPwdDVk9kQEQYDkWIuQSaZ2ID0xcVKvUus+FSTaQ83C/x
TngETjkXnppQ0TDU5zh+L+w/M/r4ByxSAgRvt1jEtqcLPDG1cX254Izt0Hjofy8mbkEOXyZB4yU2
r4EJOXIO58Xd/uyyXpf/FEdyKWltCTwpF0fl+2Olyjf7KD9vCeJAeW0scL4AOwSQIahNrQswvzWh
3mH171PsbJup62DEm6DlPR+2njuaw7EYEXKqoffS7eDH8LAUKINog/DDJno7PmrnDFiDWr7kPevD
93RpYlUrOk2oaFojLDL2oD41tKNC3tRyvw3+W3tFX73XqQ97g4CvaZ+XPkr28/JC0TSG7xySAb6s
DwzKd81VCqBFEXZxdBcTd4DjOX2go0MTxp/hL8FgJlW8qAQHcIj+lKhPcfUnSp+jZ+3uzmfMXGCw
rTdWv87A09FBhYdPuEjBo9h5NzpL/X90E4FQsgDnhO9O7xkk9/27OIxInO5b49izQsmHdPSGFQYu
Lcb26/NXxWMj446KKFierbfhfTWbifs77XQDPBuE72ud8XgBMvR/1R6/edavgV8CdxUsPgSMAZXf
CvB0vDfTFfW9QIw1saeJhpKp/Bi3Oux8PXOLgzRYJlCEC53oq2cmqODS21dSefGSAyKhq2DeCcok
cFHNct8wH64/kmbPv9x/WMLJL8OHPSTAvw9DJBJdRFCp9HbRl5bplo1QQdazbujDSq5xjUsnB/mo
C93Gc4lIGHdGtnjZd8MD017wusnYLVyEytfNSNucBu6lW2atM583FqIhoo3MIr+OCGPjTr2/H6ok
sU9UT331p/TQge/KamGMb8Uu8sDBgVgHDZU/sPRMw1LiZ/w9O1feknX3lFCYK669CbQ8jS0X+V+g
Z4JLGPjYJak2oPCEM87nRuiztN+KV20BvZOgkPo76dHL8r6cN7cIULST1oZ9+3NEXsLgWLINbEyP
wtSTci73yxpO/qggOua8MJYfTBsE5rrYZ/4KN3UQ0WE7NAhInV165IWeZvZrOfzioC/zlh8EUBHq
1HMPHwHI3WltkxnxIV/4/M1gVSlk4awKGWw+VjAdFpqGTsuFd904hGqxbg8iP/VdfVK/1lvJkjSO
TnafrFJp5j7Hud88b/N+JbA2/voc0i7IXSzFQOQWSBOAetalnAZ+CbuuDRgs/dthmSjYHIAjy0nZ
Oyrt9IqpCk8Sadri4Ea5QEcrpu0xEItZBNY1Uuh8U/XoTdFmKYcZp3JOCrSnab8Oyj8Dc2BLRSu/
/PUkf8fVgoTbm1DoXlXNc9JmuhgTqprVP+ccaLiM2vFRccnpJNOAYYGCk7xH/nHjRM0qCbn86w8j
i8UA2N8zmmeAUCJQan1vKan3YMJ5/zSoqmoG3PnKR+hfoNDzO31QX0hev5ZCxHGRZqqF5GVBL83/
Rqpc/c/l3UZ5GpC7/QtYAbx/2b8aLkP8hgbHZm11ktCSHZitD/v3zLPB2shNUZdVDOp6RKwSarmL
4ohpb32ayyeaC9Lma+a/6wfnbiXPFNJ1W3E2BbhRxOBd37P4yR3IuckN5LGXHQIZcAr4xfbae7PX
atfjNXuCi9/rxNfqvFLoa9yJjy2dZgnln4k12XDJeChn4qsms9MJ8/OQo4emCwtxNGc9EU2FH925
PVqsGpHRszOUb+WqG0I/b/LpKu8ycIF37aQpKvmx994xIxTMcNVqviU4sfEa4I+M5r+wZWiMBIxL
4FERhk1J/LgfYajD8GVc82qmuw2P3LwD0eMPX0PdraDZfW8h8brTIL/p46GhnmiHR/HoFwv4Xj3V
fbnUez/LuXtk5yKa0NgH2T1GPVh4HOTFqOa7++PvCRwP6DaDBWBF41ceSXL5HZW2RACFj22OvNcE
fva0SlrHMoTIqolYXNuOkjxSTb3T/1oD17x2ZJ3VQDhikOasQ6Lb/uOJ9CpemWBMyA7rQfYO0/gy
Q/dpTtDgnEtDXUBdUA9SETSN/3ao7KO+3OA1PB4lAlLLzNtwtbHYGk1JGua6e9X+hlxC7Rnij+1m
bkfykS1Rhr2/lY1gId0VFszzOJon72Yi/9jgXKHM10JERzl1kwhGCF1N9/Ywlo4QWwRXaLzJhR53
773fsB03prdip9yJtkJrkVXMN+x8cnrWtABOBusVGn/eDkeNpXY+yh/ci8ZV2+Fo7fGWdH/gQ6za
Cra0Oxx8CDYw1H6YSPNEoNVXet2l6gTXJjGQcZZZjWnXgh87JCtLCNFblaR1l2d5pTQLK0wcnBb1
GVV2Fn8+RpdVL9MGRsMVMwULacq5QHcaV8Ys2vXLKiTGWEQc8FNtD1dnAS9D4RDFyjuS/NMoPcjg
xj/Yi9D63Y1v4j7MxAQzjET+lzcBVfn5WnLtoDh447Uybfgg5SrK905IE/fTHQKYAMPdf8mWWwZc
+1Y2TiMknwUZSd5uNUYWRoyrHPCpP5aPT2/SFOTQQ5hybNMPJsfvohvdsuM8wRBduOpzCwRYt4C4
ATC58TrGRiu2RIF34U5higLiLLQe0j7cPJ+he62Fg9g+PKBeoSfeZhljo0h3PLtUQbwVW28/SpZa
Ns1JHNUB0qWJlzJk3RoaQ1CxTX7JHx9dVIw2ZHaGY8whQUVRYE2g1nT1vA94UDD6R7LxSIw1W4nv
sxAlq7tukL/BfyE0jWcDC784WoCp6JdQx5SisKEhkRE0OPVICaiD/U0wyGc6e2J/ziUNnIjV8TzR
u0lTTrqo6i6tOC11Xn6bUveWnBh2IHAjJeuueLhQRO/nNd1yGSXfRYMJkhXJheTVMHgg0EmQ9GF2
RtSh1V6QE7dQRB6g7zH80r3K0wlropCZJLXZBaJV4haxDBgAKyTPIGd6OKEVYw+9s6dUhI93dZcB
rc1f2+lHDegcCc4ax73Y4A92SaNHPl5/OxYQ8DCGxQunhLKryqaOZiFkbQx7T+e4JWjhg394neYX
I247l5c9+HNohvvL97aSe2Vs1ZEYaF/S0onWTOPQmZfhDKscVsn/+uKpQds6PHBVJZgTVneVJmag
gZK/PPLNv6+pO8XevhJOFFuoRCoRyXy8Z4q8FgFBNwARdnjMu+1Whg8RaqVVun5FwyqmwDWSkWqI
KOr87pHRL0LZZ/DK9GvXqg086xe8VgzmXblpONMHYlV0+/97SqDb+AbQJAQhKORt2N3BhYedeqIA
bDuWEbsswmVeUcIUbh6d+FopncQTYAISh7BV7tv/h9LW61GqOEMj32essPYpT67f7Ne5wc4r/dlB
3CF+HUiBsVco5QsRDJrMb5KUAhLzy8fWBIIc7ocvY2VGmhVNgR0t7K78zDs14N0+BKQHmWzHOra7
06ouL3pnJw2ur1+aC1PI71cmtdwscWDmKroi3TlwWGyVvYB9DDka69ZbFLXF8G9SqBll3lW6izfs
Iugl3+xKawaQUEDRPLxI98a98VujtxV3hzJwfmvvP71URk9E8I1QZ4wT7Q5EiIA9FFvKUIWQWiNQ
lzIulC985Lqz4Ne1CADkBEWt1r5QIf3Iy/hos/GMMpekbRRXYPuJlqNRDrKD5E95oiaWOVinDXb6
1o7nse8k4NuueniiGhKv5wdmTtpK3IDgp6LzeszN2hcKkA+XK1RkJ9FqjNrxq1Ru/bSuFXVZ2aWr
UDZ5wpPadyRSlrdfmzST45XPjLVN937I8yjN+ch5+ZSUAhCukK607BHRrsLvK9LyJNZ0i8qk51mW
04zYz3iIHyOSxsLn3XU0tkP/FnQYaxukGLu0ub7Se50nhkMpFmRo3iQAirlAiyWYbQt5L2T6A9YY
u5eC5CTeiYgkn1IHJSGPsY3C0UAsEaaDHlPPRzEekdZiMcds0TMzYtlhibYyY001p3I2gNtGKLUy
Zi/UVEbaKnTTo41lTGKHdA1MK/Fm2ayl3uO+UGSikyRvQ0uOAk/nRPXsYzSmn7HStgi6DiFqTLhw
mX9SaNf19o7WuSn3AkU+B1Zy1djwIIv9DCKVdOG1h30OiVfbK7XLQFaU8igO9hYtUCgI9YepM1uu
O41YiKM8w1dY7LcD0NlUNr3SbbczqFoBuHBm29WLN8HTISbh1RvG37UQNlp+2Fo3/Jqc+9ZsMKTD
yyf56mp3xUJz5fNVHHpqqv84My3l6B8l39y9oNJDxCJRywzfJl/8T5CwabTblWks3hY2fERBFgSh
NlVEHoFNaP6lWpGIHiEtqM74qRtUZwUSSyjlStJn2M0xc0w0Xlpzb1qQbq/NhOL8JigqtzV2pD7k
po00LURYELTO3qL4/JJ0YHmSM8aw+YHXg+gsxSfTSdNav5ul+2D+IaTl/0ZPbtoV7yOIwvKPZun4
XPLzfGcBya5nStrRymdpwJjR9lRjqXotlm7Koa3XJvteQAtd95EAGJVa1HYMUJFn39KpLecvblUb
HMrttP/qK2Ugrc1c/Elkvu4XtCmSoP1R/uOpubREV0kQjJuF/fFMV5ZpJT3q109IpT5py5ksRCzp
jcOn/e5NJj8YAWANVp2KruwsWAi9xWWg/Qi20c9tyZRETmg+L7Av50PIQG/xGxayFygqBBQ9+HiG
LQOtVy+sT36WzJv5LS9KT66bgXO46bC0DtLan/pOSB+9w2OfabsLiMPPXNCoKRcFua0tfPrqSjlh
a/hNq93S2/ukyLvz+hB9pEqyi5Oj8IUM29wHHUUIZfGwpegT7m1rPGVJwzNVHqWDWw8xfb0KWhHs
AntJK5DQPfsiUFt9LSxfyT018t+lHhSx+v3kViSLwiJIE1Kj67UT+7j9yaUl9RqkG0yFhwnyJSLk
rKMeOlUBnsg7FFGGShCW/dM9l4OGRc2DzzDwDKU2x5methsvyG66PmpW/JE6QUenyc3o5mTL+nzV
w1RGrLIj+KvJLyjKkGWKZySgdJgdACqi7VKQEzDcQJZ+8YSY/PBBRajTM7E9X+QPPDPxPPTgFIoV
tNDF0p4qUGN1D35kPxzd/1qhIgwoFqVLakZMU+L5lsvfSU2KTClXtnlZhZ4nh/gId4oMLEmahZQe
DAZPl0nxs3Ifslu5RWrZJy9MtasTbcWvjYiWCpFUq6feud61yRWL9vccCvbyVyYf3RG5TSDH5bb4
deGnx9JRZ0jSnr7LoPMPOwQFkxzauebY8aG8D+PZI1lO45UwhuzhXdZ82uvr3LTJQtevR8s40pgY
BZNBZAETz+kVQHKhA0+J+KlwG8IG0e2vlhkvdh10kmGBg6qs7SNTQiD104LayfxD9laKVbxfJFHh
lUIF04dXwKBWEm6EvmK6+Qh4YUMxDEV79Gyu1AdZ2PS14wci+kFTrSCk+x6QzVCaGJ/W9D+7PUnG
gl920VOzW5paoeEqQnSnJkMwqMijXq70cTKqjhU/5MmDc6FIwZm6aGT1vytbM4t2EKGrAdFa7Oy1
PCqoqqCSP59s1ximea56vgs4VJA0anUnReawrVudM8PWSTESW+IgbMtw8QL51TrJYpCICl2Uygbs
ZUZiEhQnuPSm2LxPfdfw+zeKHV7BYswDde/Bqu9uxu/qlsaj/CqXoCsA/M4UcdJMYPvVZVqy/kcH
iGqTmoYF7KqB0AUbVkFP5sQHpkai+rB3JtFlJlUQM/cnc21MHkdMYqITHk8Tg+wW046hOMk7G1MH
7W3ZfWqV81skqExLVBZm5ETF/U1G/P5sWshEdJYoMWvIvcSd42HLl2YB8SjdE1/OU/nqiUEY/QC9
Ox46sPG9eLMGNqmAgizxLbwDPbJYMcKsE/lzfnR4IPlvp2i6V1fshHSpVF3gwiDop9ah2GrrqFsz
hWADPzvitjrSTimcvVRIynMKNOADJjPeCiqzUcRSrxLI4d42VaGqFvZSN4UEqWVqoZl55+WmvU/F
5nGTjbXCuFKeedMEdR1IQWcAwDa9jymc01mRgneJ/gHGaLT96g7aZx5HJLUoCCyBlVcFPgSLNynK
SI7hEAFcdM4fsidUJ7qyWYRmKkWZcwz5JKra/UTbSOopd41IQZSGCPQoNGq6lXgr7UgfWGyTOviH
MZyL7HNCr2yIQxGjmLGuSv97i476Qg7p53MEGnduc535roeUfOV+meX47UdV6a2uVSmjim+DXOJ4
uZ7/lNPFEmmZzSOIJSmNMD/0cydIXF7DpIW1u4MqHEwn5SIyP2tGt2RhctPIHi64BjdwR2ZwxqkW
bgPW19N1C/CZivxuWQbzGpTOgn6F2zwBLLgmhF9mHLckxtaEtzYQx+njqvFYwi459HwA3tE7vqDJ
MyDzAYzPEzQVsiu0uHKmk3tZxgYqVq9DzmnBki9pKimnQOKzHKe/KA65Ct7P7KKYriIb/HA/v4X2
Kx6vUg7xQbMvVQ3NLmtclg3X+G9QxMJhjA8l685h9cdpYH/6qSuYybUDQCXhCPENN1vD579VdHyY
R777cN4jhBDml1mu+szq5cbpvlpB5QUc6vobeC3i2V8DBIpJloshhJ0GuwvZpp50P1tDLSSuqskl
XGM73UBnrWczOhlc5iwkIcQVsllZz1XG4/aHvpp6vLqwepat2C7Gx5kTmxVgY/KM0pkeHt2M73yX
9SM4UGdbME6sjv/6oeKKU93Iqugb/YPuMKfguTYN85s8huN1n4hB6IU0E7DdR+aKQ5RXyNshXGU1
lZHNo2UcIoEqoJx3LgOmchBLFAOcp1KwJbOI78DaD99H2UBZeRLe3PdvpU5oO6K5hXnidYNovgpj
DA6H38Fafyy6O/oTM9oBG/GYVHQa7A/ZdLsVbcpodExd8yg0QTCzWfoCpvXPT3Peyl7KHoe5s64X
TZA6jIrwY9t4y656CCXsb9d6JOEydTryf4s5ZHEF5KVRKqxIW+zL7lGVlGxLpiQse3yQTkAfeqR4
LZTDgxD/OdiVOXsPPiwYxi5HBnvoOoIogeenN0Oytv4wmHY0BwSvmU9RX0v98YWqixretYPDmCEa
Sio5B7HEa2vfVp1/3qe1NOS46eTWdNA/3YKu9f4UZiAC8QjdFuEAuOXLEbvV0L4EbDRuM8YtkdPr
E0lbL5nSPYkUuLK1uZbdO46HRn7qbhbXLmI/U7e7F398Ok/QsvG3lp3xQyfoFYyKFXOf253f82zG
IO4j35ls8P85TZ0yWpPEhOXE1CJFvKDkUr/z9MnoQcPI21Sf5VbckDC8Mfy9e0nu3DIxwwuv8iGy
iNvkq9u8C078Aoh0SdqoKpkvaiBZfZCaSeMa10FBrxVRBaV+peUtKMQ2e39BYLzOW64KTmfeTARD
9ou00jAOPe2pNCMlsCSkyAJTTuHwUgHEvb3zRljXXUaYhd3l8OXoRpmVJpQXR1JUUVlcwvhbt9iK
9W1wkN84lXSSA5XCNfUOHaEl82z4qBabJtR9i01Ws/088ST/2gA4imorXoFblIGf3OnFc5DboDpS
ik0CYazCwcjslt9E+kLWOXy9nVwO4l+OF7bE0s0glp+DyVu09PZTDYWWpYMk2C9L9Ebt/LBfaOf8
JSvIlcJQwWZcNngKymcSazv8nJL3vSLfZyoRREjnzN24ARATrZ0CZ6GQGQXthvnJBlfO3q6Jeih7
GWfsP6nizqON7RqekcHuUY98FkDr8Iuprj7Gx1lcoJQZC4D5kxaTEiCEnt/hQ72pKMyzpDhWIdQs
irN4w87G5b6X4BVxWxfu6j6YoY2tNGgmNnawXvbeQVQZeHAABcJrTWmpYd+EQu0PB/flg+niU96a
gzWF+maQ/a77OUIxNekVJ6iaJG0v6LsuLYBIj0ro2SKwx4nhJ5Phl9McB4PQ6cnMAugat7esqWOe
9um3wta3pL33EFkwHJG/NdwmLLCR8GZMY7Z7IMr+oQV02WjoIhzdWwyg7iUY+PmIc702hAATDl/b
2cmM+uO3u0pSVMT6b/F3ywSITcYxhbGHo7JewuvQv2S3hzdOjAn9iuJUnbgUg+fE/2ODOrE0dY8T
MDXtfDG001oSzaLCihlWhB+yCqGENDBJkvctYAfsI5p7BJaH89oh7SccQlmi3D0hkL3QN9+wmlLQ
z5UI3GpYDPb2pj4Gn8YceNyfn9KPaaSHP2ddM5Ir5ENqt+z0f4IibCV7dRXmxD3fm6EByJ7jdopg
k90ghjmOK7tRLPnpaIY0HW02KNbwDtnjPDr6t6f9kYXvYJgdgVrXOTqvcy7OOI7kvtwXuzzE1amX
25Sy15SJmTa5h/5HKNVohX3AFXjNOl3hUFdc6oNb+Wrn4499IiukhdJK1tJdqT4s+s04bSfqPhMk
ZHExCAyC0CwKCWoMKObkagAD4b4GFCPDJP6qk3c0UiXAinOvYNBvhTqqqU0ngvkOo69GwVr7uA3u
Vi0APHjpT+moei7Pr9zS0NJjj1kE/xsIGvMDOfymwU8MAjWujl3F7lhgivM1sU6K1JH9vgkJNw9K
h/91htIzxztKWyQmZqxFOcB6w36klicOjAUIvQz0raXQjBKmsAFwj1oBa5ShitzESH5CEGX13uQU
Hbm6DiV5mb7EWhkE4+CFg9wAGGOCLfBNAIehlNlKDt2coIcPRYHWPnefwW4hy89/VvXnP4A4w1R/
OMXx6E/zXfEl+TFQxpzrY7lgWxKq1akd1mXjL6tUcyD4BeF5VIvuOfcUD/6iCdmu+9dzTyLhgPrS
MLSxs8C3dZKJJJe88brttW/3WqaBRXGdWhtxOZVocFOQpOh+G0BKBEm3qMo6G3qqRfkX+epXlZkw
pN1A8fCZjMeS7QHiJuqvV4tU5yePb1V9nucuFe5t7dwPSZKL8ArS1un+vOg9R3mT5fxr6zuWWRml
0XJwOJwQKomKjayoVVuR0YX6YNYzGcrzq7LHJVlA23Ag9raJ8qcGFV6SJ8d6gvZL1U5Nmfvbhnev
WEjBVgStYxpm2FLx1S+8jpQZxzvn8tmtajZIx50mfoVtWD9BANwb2t+pVddHJXcQpcQqJLInhgbO
c+94cCcytUhn+AnpxfQCFodEmRcGELxFZg1ICiP1jd8QJgzY9M4TdGb2xANTOLTjxVJznfxZ1HIn
AYuRq7OICEK6lt7B5RxKXwK24bSDTjjY5sI7SIA/s8spD5Vpz6jn4YTnIQDxFWouAz99uKGCpmaX
+InUdpgtVQVn2DuCkdfnF9IN7x0B1c3X4xzZiKyDWTUZM+7AaYBgXIJQQYlu9zewlIg1q7dyM2AR
fqP1Fg18bJI1MvOFLcSpDeQrrLplaYvK6RHS82FmUsmE/PQwyCqsPSNz2+2l4dmC+cZzR//bkXfT
WMecPnaki/L/XKDQvT5ys4Oums6Givhsf6r7h3yzgWrunCUqSuEd1IePEF8q4NCvy08zlaOXQtim
AXnhd39r70jJGDacDScBMqn70HDd8JMl4xgP3hX9XFRMDjfyu4lISR+o0d7Y7Cs3KlHgWptJqlKN
tpAgT+3bcdsbns08Sfl58lvTiddtgr4sbjARGJ2JqBM0G22yZD8K0lEb1SgwgOaczgykf+QxsCze
+4cvwTFaIg90u+zX+zpvcr5g7UNXK5UFSrqFzEKT3DlVYy1ONeIirZn0Kzjk0wSZlLoqhM97Ulpv
+jckM2JfrZcCqcyJFqkioG/RvL/MDQRXE10p0ncpO1CfLL7lxzQqSe3VrcE6/7xvh4aU37QLRbRL
iNi5WmZFNy7FgDjzdnkFiweAPERFsrAWwJssqv9bOBDomwLMURXdqx6/+GZdZbYy2ogHk22X3FMP
GKEDiboDwywgNfskAZNS2aKRZXS0GpLv2pZRW2/UiW3sTckMpTuQ6zQD7Tn1v7K1upQkTz4/Py/I
che7ojG56/t8xOuxMswNnE9ZtUVXFoUwaUfuVRJwYHD/xh7utGeC9Bk5vE6QaQBQegJj0o+A+zzm
Xc+wOiQ2mTbxBtnwiP7BDFcgOoHO/zQtKqSL1y7/1b1RTX+N5a9+JOI4ZblFnKxIq79sqMA5OXCd
YJNU3lmyf2OgbzvswNwfmMdiPMPPAvUuNA7dslZSAPT7axZknvgyly/YXNRkBXd2wNaY4U935to9
/gTrzSZwpvRIfD50hsnme7Kz12vw+1OzbQze5SicHGtOCesVrj2ZVaNa0CXAXfl/WSPUGbEZjHSK
GcbiQtI5GK/tm1fNsXHOjE+rJ7ugfHhoOZUCx95uHVHw8iYmUmr6s9sTEkmC7DhBWQhI+vYTb/ZW
rEd2gf26THFylo7Fciyrqc2ztNESlyZnEX98Cjfiswspuimp87TcgxJXycuJ8joj7nGwVb6CynP+
vZHKzcus629VYItiD5glydRujpCpUA8c8U6uGBt4bbKvY7t38eRYQ6qn43YjWHFe2TAqKnI4Bvai
9qJ0hBqYySfomejGXiEHKmF/HDE2p7HqmLIM3dCy4Kmjye6nRbehQe3WO7HdG/En31smtdRwLvd8
LFAPgcQz2PK59/OCnN6lJui/JVbwe8MdCAs/gVUMoqGKUu8o2Y2QQjEYu4tLiDrL0Egbae/rrh/s
yYOhZSH/DhfCiNHJlcQU24ZvtW3RwNUF4ZRM2y8u6rPhbmw7fqOV8R4EQVu2gshX4k9JiCIzK/iP
LnPOt56kUbhePe2Ggbjb2EArWApaWn9IZcHg1c9PzP18QuH+Xc+feiot8po9x01FSZGcTfhOqiTE
C6UxbelgZHVcS9Bcoy2mrfH945IWiCUyuZfICMsRxyGyQp3cidfx9feOXXZPTzrjx/BCGHZaG+Yp
HUZAxgYfM3UIwyFzIHHvEXwKkNYEw/Maj0knxVWl2uaMNH9Je3r+s3GFEe7Heb7SPyf6uq5G03Q4
MjB80RTM1XOmqcrXHoqMVWrBuuhOBWj4yld7E6pMTR2bdp2SFMUxOU8O0NCUWrI4BhM2UCuzv5H8
zHAcfWl12Rud6jwDo9q7So2jvmrWffQAfLjVAUd68xpK7ab2fzZjlQ18PZbXOhxZi8eop0Vy/ZMD
OznhorXjcTIZrlNuE4Z9GOv/r+O/vpRZQ6HJdQMlSRiTFRqhs0pmodwMnHciKLWPY+AtC5CXF166
Sn2pzg+TJXAVbmktKNmZa6WmmjFeearklvRBpu27yj1x3USS5Mi81ta4iOynsOh4PqRm+ZGDnp5a
5TFovE3fRm+Sb7YU0OCAMf84wCRnMjG3OxFyj364IfNCcYJNcTp019vMtd3go94H8c8G4uM/Rzu4
0aHUMYt51JPIK/l17rRZrylgtGpGeHjdHlMpLQi098NOn9vpKWDigFmpO41iG3xPdnVLVfJALhiU
Vs6udq67CwRoNjdfJvmgRiuxVET198Q26YWWN2AAmUU7nQ5Qhap7RAldT8rXyq8QiZLS6zgsd7ZD
qc+raf0TuEFDAeYHxy0KaQEJ1ryUzbbG/jmMapI0zzSlqXIEdExXtxdoGR7++uHH0M6+30if2taZ
28vTXPR7DHTNBsWFAE8f4nKWCVT3w0p4xUtA6aXEnGChXQbT3k/uPonmad5EZvEjsD4B7ieDhqf7
zDbQkOyYyVqF2iG3dUEEOf/Xn0MX6GXwsDPL6BpQrX42yWkbrAcufeQplK1HVkzQbAnZrmDOQxNw
y26GI6ciRuC/K/NIQ5FF4NwWP1gwtROiG2SWr01AFfqRiqxz6ANFsZmbqK1q3K0sp8XOyhGfp7WJ
YPG4fIXaythimDMpxRdfUhNEVbHzSff7GWo09OebBcBfN1xRoQEi7i8M/vjOjQLLU9b7UIqY9bya
Mr6nnfjw138dB16JN/vxVXfa/JOVP5odd8aGEUUKb3NmyYn8nupuk9aNSougRLXm3EeZeIUpU09x
xHilFkJiSGjtII77lx8O3w1bjFzsv6Bj3ViSQkDmMcmzOpLTpdYZ3bDlSFn/UOK67JG6ZMAkWq90
SfxM1C6Gsy1LoEcl4R11ovz8WAEm7v7MlBxAs/4fb7Whp+BnZ6u0r32uX5A2HVnqDCwxAhCizXw7
nDubcSttDuFCMSX1P7mBFapJdeW14H3PDe3Q+dfUUSFmVHeqsrsBTUngrFv4AENIJ2uwtywGQYIx
CPO9L/dCHEBNfM/ykTIjFYLMtF1iRY4CruoTfihKO6eaOc87dJ6JM8I+BwxqBRg0k/b6ipEO3IIV
XrZg7r/HYMCoeDQyQxCDxRI9HhSpdiCyhbxCu7LRbnVr9up89ZPAs5LtQ9WFf9C6RA/F0Ei0c34Q
coE+t5OstR3HeQsUloXyt3BQSWD43DZETkPjcJLvMNgr+bwU0/OqT32K6FOVnryT83jgHJ9JVo7N
uMd6q/hseKNHAmaqrQwtJNnSwOck/Wrl/rycGfv7JI4WAYA5wT+YtzEGZer0vPj9PwzEpbn0mbnD
eteZXWQnZti0wjvjGm654I14nY/6CCpAynM7TbUjIg9jCAGtbh3ZI3vHk+SHI9ETX+klfz7Kzuh6
uFtA2VblOumRxxgtetyBDmB3tVzO1Up13i2P7oaqpB0B/0juJR2Am/tKoAyuNLxnzx1DlGSAYm90
3WkTc9YKFP9kq5AjO6SMFW8fGXfNI+bqCeruav2vfvp4I8+tQRSoEaYsIcJvc3svQ6KudL0fNkw0
OaUqWtODpw2FW8+VJOiRclYsuVne8lPTbAq9rSsNuq4n5gWv2As45LShBIZ5bM48bFBaL+85/naS
8PnCtqWgaz1BQaKCXMwRbbVjScQKFysLR8RTRbUd3CUOAYcJoslNgct/EEOeUyDSl1EQSzS+n41t
pCSlqXjUrVpWxqHmRVleu+rSfymnIt1SpojbIXU59AACIYu1fDu+Vb5hqpdpco3i/jOkp5rWVhS6
f+svzNk/kqqpb25LGKwENP89hxbIA2kUjA88eyD07rjK7wEvC+zN8GpXf60mWOF8mptf87Srl/OD
Y216f6YFjCFKWIEccgM8furacEqyVomasadMjQLIa7EyiLQMKkd8UhiODJQpGo/ab+RdvuK0S/Yk
mt7KEt1oaF7cVWGYIcgfrOHuxoyqq9Y/Y4Rb9u573yCAi1U3SENhaNL/inPa9H1twNII/+6Qb6Yb
t3PRXC0xrfpgxhgpuhvoYC3jvFBqoV19LnZzYXlg+zDDdz2+4gEK9nr8pVCUdIHXccd6xt5j70Hf
3/0MniChiSugDUb0t38umFIzdhpAJtFbSJVSj7DHB2ZxhqwKvUvLCSl3DCI4ytSyJLNB/2uPBukL
731ZnSnO0Q1VOvUSKzesv+0FUm/YGZ5QexgU2QYPQ/3agOIscqdyxzbYiWr6pS9aynQ+BZ4U4bug
mtuDwVpvrkraGKa7wTzEnJ1pZxGJ54KsleIfdmDp7EhyIaAw/ZImoEiJjs/8iDTbKhNoF9divNp1
weJCB6ajeqrwiMQ6/NHdR61XD5hjFfYXXv2VWG5Uql8U0CAjLDYfaH9JCwT7kaEfiXo4JL16lvVq
TEbbyyCmXrq1+cUQlI3GZCZnWMs3T4i2Be40kiDQjxZbKLfo2J/RvmX1vrdANc8C8N2eKnMQ8Enn
tpFs2f564JkjugXOalvAF4NebUm/IpjDU6YWEAp1+o31viiRwcoLAIgFyJ62B153pmkqsarzE6Xd
xplGZxpRNg9AV0UNV9FtipOp/u0ABuGqADcxTJ4I6uiVQBTbHtsdHPNMy3gzO6Kl03e8uY8w4qva
Oca8JgzNPMI4660c7jZnSvfIp5V2riYb+oYKDEReZc1n6ZnJbK3kTvgJp7KRPeA60Qwk7UA9mT1N
fQJv6J4Epl4kEoC2a032f5HHjVQy8tj6NH/UWhVrnnfc/a6BHqalFvKS4kN5MCA5mpZrJo1Z285n
v5ghs1yXwpF+RCgWUJn3GsYqJy7ES8C7GoMRXVgEyOadMDPkqp1AnHNwzrzPV/ikoJgLQeRp5cwb
Q7pj2bYKCIIXlnvehfl3AS1bx/lSbz2iL8lSdkgGYmeruzEGg9jUHhzTbBj1qdvw/w0XGRq7upJ/
hWYDFVtt2M9vFD2R2WZhC35qFoKR8yA5pkcvdEDIVV5Z0d5DGzPzdPPxF494j5+BnKr5NKeV6Qk7
aDquuHcfs8xVUJTMaK6i3TBrv6BqAufvyoFsp+EzPFudtuadybuCAjMhAc4b8qv5zqsjh7NOgUQ4
4Yl92xROZD50O5OXtk2QldUjJ2s3YbnIdXtnbErYL8RSgx3JG3ISN3BzWu9hEGRCdE2Prg0CKihB
JXZbjtbmNO88sQZBx82Y4laYLEmlXVqW8U+3m5+IvoIdFjsGHUTO/fz67tgxgrXf6IQfuOHr5lQ8
wXwOlMMfO8U0IHDXOFc7SpGmrvq4ShsS53l62aspxYifPcljDVLHythC6Nhm/Ffh6gypeeP6r6l1
ZE/6SMoZKEZo9TOIz6Ue+ywcfwD7H1WTAQ/dO42o/G6CMhG/4ERaNmg+ninAtY1baz6X+mmh8iAo
CHZwpt2CkbHKwvrwT1Vh4zx6ZfJlv88WNbmpmlOAR5r9jsVYhk59XPNUMlR4YrDkMAZsMr5KpNUI
1hlGW37HitvWmyhFb89ZOu7smt9P6gb9unr81uKsnHIbbAvuJ5j2YOI3jJ8h2X8C7HqiGE0e2Pj3
jEFyZsI6OU2f6g8sRqKq6VfBvbkspherfSPdxCjNlFaaPgKeJq7dCK+EirNTNiqDlTnK2fPjJ77H
qJhqxbE5ntu7GKWjlBAwN/Bh9hKIhz7Yj6TbvengYU8LB/jpjOR63H6kPtwhmOrVLgoWWoq7KHak
xLOM4BgZUCi/gwNBDdUi1FFwI8ggprI9BOecmsPGJKTuCCAwwkdUhQw+Zf8RI2FOYqEZgDB2XE1K
0BwWe0uv9wHYhpsBDGK8c7Qjc6JT69pDVHnnQ1ucL5uQRq5MCqcFkaZl4nuIw/T1xJKCCdEAVzNY
JXhzTosXVVKLOkohVxy6Pf1nw65kE62w8UJZdVfltX+Ir6qeiH3ixV6U3WUAfYW0+JAO0mh2mpQ+
V92w3eGeXjjT8TxwAFHkLOAaUet2+HORl51hLhe4MoVY0cfEHSf7pwAPS0ayOMLzMT6ZVRHv3zTt
AyCl1aEMh0fQyhIjANRar8S8023nmiykiJuZNcEJPABPIJ0b4EwcpDRtShvQ+5EIkfSuh+/t7oPM
x96jfbfzeJ9nPWB0k9tlS24h9jyMPDkzSf9aMiIEpOuUBtnymNXR+FZzonZpifdwpG9T7Avqu+VX
Pcusy/iHaXGv59QhW4vQtfMc/t7Hz6v8Xt7CEym3nj4eZcPl0uWz1sW2B9vVN3hWHHr89ZMWglAG
l9zovJd7t7aW+XPNGzhA5CiKD9zabVLbV6VFqPDV5QiETulK4eGaa84SnuGbp/Ubo9pcoxrZr11B
/ptCNvbHD8sHxc4F3ocWOp1YUztdMdjHWE0bxTRnJa4Py1m/y4Q9AqZhGRWxYoJRbvcpWZo2QJTT
ci0mPaBAb0BVrkrcluyC3dY/7zrnH86UPtocWBN/bUvlYdgaNwU/aSRl7spDWInbadcMcTILpx98
/vehSioJKE092oO6tStIDk4YCSckZ8n/3ohDGaVSp73y20KSNEUfG48tmwmhEabW3l0eqDjQEVuo
uFYRl7dQDt8F9JkPZX3rrO/B4oSnUlIZRwbYbI+nXVA1zul5X9GqOJ+7I2z1X8vn3ZmBft1IpWh8
gGbpKYuHP1wYh2PKkgRo+YixdWz03KX1gCNCKJjKuXpUeQX+uWu6J2RlVsIb/rg+2lZsehOtHiwD
TILkhsvLfZXzTxbBjwlXlCrEvuWH78AfqP+BjfoPPiUCDryqsfeCOn4V+E9TaHFlmpRMjV89bm+a
NSEiXcfjUc3Y0jAhCBDpyb0k2ktGC/lerUODhEtMMH9W7BXbguykst6pBgtIahxOfx0TXBzEXHz4
Fxln+5Nj4Osa/JUwnCsHPlXt70Lh6UlkzTWP98V7KzrwamizUVpXMvkFyrBujhOAY3yBnJC2jrSQ
kYq6OYflJ7SA6JFgc49PnWYUF8n0URb5HdMSSMosCla4xYT8UJkkbBVEBJgaLhSayVrnwGx9h7jD
EQmc6NFelEDSNnVSXXqF5TczFYZYvtV02fAHXBVBseGSSd8HMNpO/qrOjGjo2xdpl1HGbFEPG6zc
vaiv+nl+lg/k5jIO5/QaQ4x24QgqjFIdC+haYxRYUvWCQy1ScH8nMdALVrPR1VfH6bcERbSJ7e9b
N2zcl+I6Xi0pxFBHVhULZbkg+phP+k7c1pYBVcu1kgQrLuPgPkeWXL3peJ3firebAu8cwfrgMA+U
8P16GwOa/y0MDIiEeQr9urO5Zq4K1TKkG6DEMBz9PPK++di8YNCcn5N1XjE0G5jE0mx7zqMeW03p
yS0Z51qsFGDKg3suMaBDk5tlh7HudFFApbA6IHQy0a6Kqz39yCgAXK0huzHG5/SCnGC3rL8io6V3
r/aSp3244JunF1Upspw8R9S9Mx+3+jN6ToTezPd+ulWKxRDmhs1ILFqWUo3o5pd2NMjMWXsJ7nMa
cZGMuXul3nhNUnsMxesC3xy13lrD5ouERPjxgo6q1n7KA0as5x2Ktiow26KUY28u6tritcDO2bN6
T08R4x2nZgOGgowTBFrGXCpSfSFSQWhfWeH2QBmW9xb7FIWgof6cELoNCfAzsXEV+xjBb+LyqAcH
rftBdwlsd+QijMoicOsBAuGnRXZ6XQtyqSIimb86Iudhw8qdu+u95qF3iA/D8UCqMOjk+DMH5Qo5
OH8VaF2zq3q8igx/HkbRZnJIDY5Pwmfb4ZTjLXpcr29nRKeb97wQkt87Jf2atvsKjYYQKRMiShMw
iDVF2F8v3VhzDQwEo5eWxKH5hB0Rzo8bWzwSr0QMzxb8KPs1h52CpE/91ogoMAMfg6rndPI045lR
WihKSFzyjeNpirGXBhDLxOFznNaOxtsMHqlWIUqkZdp+wlPW/LN9BGf4fBJkEqisMvBOVPbegZlP
ZfoRWdyNKodONX4qy5yW2mbGgNGZL9TywPiFM8887Zg/qmnFAMokKBWNSs5jQMquQgZSNxPPLJvi
Pr5Yqt/ScV9Hph5OCMJvx/K9Z9htBwt/FVtA1d1pxIJ2E3nWCrblxN27uF/ZpqBzI4SGXO3iXZu/
srLW8peh/el8mw+gQ6SfpYJxR8PKQEj/l4h85iLPuj/V7mL0d+pOFOrKVvSlcmHCQaqFN+NRSvCd
eB6dO5110y5REv/gcpRYwyF8DFLskzjQGXeZJJBeUCWyiE0VV/Odz3R/nHbk4bNlCcOjfv8Hndz2
BU5U9AwTqkVLysiQ28tY43HmFan7RUqnJ+7jYRQDp+rUQOCzZiivoAiFXD2GJJSRpXGSwyShm7/b
Lh1sG1V7YALMZtas0HNR9vfT7j2Adp8AqM1kkBMn9VBxkuzJUc43y38gPmZBbq+X8gTeDQNLcdWQ
/hcakj/thuneA/1H7gfuBc7mfzUc2TEAZU4hO0PlM+b5qhN4wnHNSgOusMktUAZJixVa6fGf2r3W
SLRmkf2jcwxSD1COR7HWx0jHN1EQ5TgfbX/d+8KYlk0oErHxfOYo6wjJEcDBlysBamQAXv8x7MGS
qvHntcOjE07q+zMYFh5o3CqYbuJiGngDlDyJdb7XuwYSXDl7GXevcgDH8+Q3nBEO4QqGUKS0KGaz
wXP7qK9ZpHZEc0Kc5dRAGOyIC4hqm9ThKWFSdMfZiOMmdUs74NIlGZ34FgGI+5j7HBMAKs86NiPA
4CjZG6AsPpTPwk55hIljDsUO6c7VIpykN2VgTBa2tK7zS55TPZR0Gq/j514+LdMelrHU3AKMNNKV
Ug1EVD57/I8HXqnUfPD3qBviTsbdXlAFFYhHK+EGBGVsn5qOBH8XtmNMoJhRVjlzV0jvw+tF2MKW
z6rb0rH5u2Iceq37QuWWrLttLY0LQ1QGgX5GS4x/i7cIgmCDS00O7SW8VXI/M0QXCEAJByqbLw46
Se8Nzps3HGiKFQQe6mvP9sNq5zIMhgYIPecXcZASFoj5H0wPYZf4jUIGQspDgEEHnDNie2rYuT0L
i+hnfeEH8KW2XBRqDPRZOElC0M/5lqOQ4kIHrmoBNZ3k5f2+Hg5SbKFvi/+LPOwvSoRt5q+FXBRS
em76tLy7H0r5rLfyyr2I0vBL6LQWp1XHcFOaxqHjKe7LndkBqZ9fwD35zFVkcd+Gg3yDK+vCgF7j
xRWQxFhGEb3rW2eIFLRMQFtaGYml0sEgkG+IuyF+yf5mDmDUbVbSxt32XRgPCLMN+JNfh9Lv/XpW
AhGMCiyZQlFaDjVOxiocizsif57yUT7pP0vjANJkcSLMAwpX1+GYdmdSxuK3XgHOlK6FeP05c043
PajXkBx7VllQABsFSRXGgmjKlwSVHNsZkIKOuOKdK+HdkPqmgarihYRVnQMhiiR+iX1o3CJLxxql
Pf49nc65En6sADOR6hS+qCl/SmIXDu5ZYBxl+JWev3sg3kMfJwSe/AA5/ytVvtEYXUzp2wtvSBau
rQ5czOGx867UtzhtQ1yXunVQC8x/TEXguuP+nxaJxmq9Sb5OQGq1DxzjTwxX1VSba2IRC4Q8tAGQ
W23pqepUh9Spvgteu4ef8jaQu3XYQiiLCBRc692j2osBiEYm2iyfUPL1svYRooYAHDPMoJ1yb9Jt
WN3BLKN1qE2n/YARyhlg05FXHgpmU7S80JpzT68XLJLvYLYALTktXfijskEionbn9LHbYi42bvKj
Xw6v4EOolRQwqyql75/IthRXaHFITqWSk3udXNKb9YB+Pe3SYgjwCR10t2//3W8TsUSS9Yrj32Sb
K6t0UZAD8UK9IfqljGYzwXISiMkIpR0Lh9Vj2wopOA65NMPIAgVekaigIDI+DHNA38W/LEhMGUT0
By2hPV7LBaOIdcThuCm1z4ZKjLl36oqbDzmvVIrqQh8ebCuMJFSwdWtSaPVt52CcaeXFe/qCe/s8
qBVEAHCV4wtdYqM8gghLHkYC5MUf8foINknjKGkBZ14mbqYhB32orJ0OVekNboUK08OJ6VZfdfxJ
vltH4B13Nkj4Vw8E2xkZMcjWtiz2Ke1bmx74iP6Gh+iyObzFebJREn9OUWo7SubANsYAHFgP+pWF
IQ7BMNG/lBgRO8s4n+WKBtVb+RUMbsqo++Bh4bOnA1bSDVypBR+srLA1d05CQFqO0ORuZ4UIE4I1
aTdyyP+7gIMr0prw8yjwd4Fcpxgp17JPwSZX3+ka7yucljyTGa8ICLT7woGQtfJXMQIvkKTfx63O
sU88kHMlL7txo3j/owyzVbcL4aTE2i/A+G2Q9Ba03kQ6MwgMHb7s15NJICmzKbUOVEDPKIFzPMiT
ln61kFuq+Xnz/FRs4SGerMdYb8IbayQolN5lJchBXpf9WLoeMBxkNnR91cKxgHakpsxchGrjm9jH
OP84IMFBatizwDqBziqN5kR+pFM20wyZ9LGnLynZxMz0AYVRZG5nUrMc3AFYbumlMgKZYH1klE2Z
pTZlHHO621AyZf2isKzQ7KJ0f2Y6e5MatElfPhTlyHfT3YgbMRfVYfQ529EGvQRMvUINrElanQDL
GzMyWuj5nEwdmFq/vKyVOBvEBUw8FVu+scCSDmdCennf/wCqV3YVIwnZJKDOgOlsJXsCpn4yu/ub
F+fS+MhLBYVgbDSHXZLhbTUJse+8Cvv6JrqvAkhejSPW179YPiFH9W/b2NvupkW/Nw8X04xWB3jA
p/fLlQrU/PfbIvXjBOMZ36pZJglNgdL2A0i2efm6UhLVc8A6APvwNp1Yo0Hzq5O7o8Csl5/2lrgd
GOxY9pYFqkyN6yatdR09YkWsESWjZ9/xgZw3cQ2EskOKvNkCKn2lZfJo2hW96qYR4ZAZciUpVwcG
/9xW2OB6RlvGEZRriHbZkH6eTgs+jkzBZe2ckk4YFHTzyXB+LUMcqbOABIcWO5tOwaqW8PcPcwDv
dXNT22P6VpSTXPJxE1ERgD+ZL73xMMuDbvff1+/lmUWo4bDnMd4rBSa5RhhNTCzk9DvTM+u9oVyI
7aTyYBv+EAmrB70tEZooTrd5d8ydcRD2OAP0eK5Mm42OQl1EPAyzMwbltT9rtHPcYJHqNDPqTWaT
nwDX20nkn5M2uSZqwLsXZubaz3v4r0GJgcaUqtxKmWtbAqyhSk6+AFsI+qBPOaKVN7RAOrYk10w8
0nD1nZ1Z3KYsjk08rmrjwkRpPwwWM0ijbz3W57lqLjSMsAcU7tEVzoMx+GLufSHw4c/pUmmKEbvM
dzmTa0AZhZWp71aRFCE/aELH7M3xHm0+tBKKRZHok2bbc5Nn1sYafujv+7g/s/aycSCjQfFXS0d2
iIQdLaSNVsihjvFUMhbXiWELLoIYtDrnaNQSq4j0pWKn7+27iMlYWdoXzdxnuG9XULT5/lbNAXF9
9ab0KVxAEWpF91ygZp1soKjcsGWhKaJ/abQxmDIF6Ie8n/G5iNZT8uRt+vq5unf9+W9ALra3M6ME
aIp5BwKMGBapRuwfnz+tDoitBcE7kDwQvOSlKPp2UbIHzcMA+B0ilAlVmClXK3TdMFCB2oMNKaYy
LTxYfzi90+puu15/Wnhvn7zpX0Gzc5Po7MaAVhTcVcYLmN1VwSuziBX3UdI+chFs8680TUqgdpC/
pfNdBP+QZ/3YXrFDlh4nqw9NwvMWTMaRy8QxN5l3kRQX83xqTrowp3Mi6GgC3Hl2Vd0kPfs9wcCP
lpo/jDdn228BGdaYvhOvSpyI5jZap9mw4uQEoT6kGaiEqHudxxWKIhj+cHUGQbBO0ZcE0eIL/COQ
I01h8MfQzfTASbMTi7ydKGiyAt1sg5EuXAqWKlg0YnmzQmvmysZ4Dhz9gh9ndL8C63cl7MqfoHMl
KNoY/aQ9/qxvOislLzW3BS/XonsWQ/rJuWXgpnictOTseel+Np2qifBWmyxLOuRVLwuH6S87qvLD
UJN7JLmX76Jj7SwTD5xfwrHelQXMW11TN/m4NcevahhMrxdnHmnPZka2uw9AN+gKc2SBjk1+BG/1
tk76YnpcOt+6nX7jHLRCyWJeYSYW2latdK2R5Qv9AwpTaJEgb7fQ31nz2XwH/e6o40jMDI+BNKBs
0cJgBhqtNDQubP/VkwBwmoQyRHR+PXkicU4X/9Iv7g7IyubGcVMyLCCnVB73xqBjtbNHWNQ46PgJ
qfnSE1WQWkOOHvQdL6t7yib2WJYs6xpbuytc3w2QMV9QM7UNwqROb4LKudq/JwyAESW4LcX/eMa+
sZRVaAF2EeIT7QslptDxLZBabcg0suTXRhOuSa9nNVERY4YheOl4GYDmAxtxdzo675/7jfY3UAMY
kjKDy6zNZnufN4McGsxnBRyrvKnXQlW7Ucx1T2BwtEplj204Pi8uzrki+JXwv8G6ZuRa2LeVA/u5
sxUYqXL4u5C4IRkG6b5//fjF0UnN5YDqPqfkAJUHoGIrS3Pxgr54B9Bgm/JcQ+su0RNSffAg1WP1
9VLK0zhdbeM82CRVED60TVDDujYz3/8YMujdN/Zyd9HjM0O8bz/57wHzE2StMSP3MDAnGdnz9d/J
PBh4lUcyv2UebzkKU/Hxmc/U502JgClmrpGbHgRSYS5lt1xOlb+JgNtkMo4Mi/qe6FnldPuzc8gK
aYZ4a4RGrKTGO/4X6s7hgbXty1axhiIMMJIXF3UPCbERDoHH3TLSA3Tfq5mtYTML+g8Yw8F2fFdW
khzmpHLGhtc3fAQlYDqoqbEA8DeLnoM5XDeaBK2OjLpX3+m83z9nt41qPdADm0xnT8Tj4iwEUZN5
0gsPssvPQcnfWZ0sciCnloYIjjOUgBO+IzOzmE6UVdker0vMwRkWtQQFTcvQ72NKpLPWZMu3bia8
FkYD7XWcO3Uklt8uExf/g1SBBNnjy0Mntdnb+pY88PK/siJNJi4GcWMDyKhTgyOplOv4qo0XGYBh
9UIuwkiKihZNYk/qbJuOsbSRg7eA/s0s98dPn1rm0Uphhy7eNK/TrHxIjo6xMRkzkU7ekIrx0oxC
dyQKqQ4YnGazWu5tvsE3jutZw2hKLasQpTLGDdAk8Xe/UF4A+e6HCIfsnMJpLM0Oo7JQqGZJBtKU
nDBrK3ky6LAp78/AIIL4jTxtjM1Z1o/66phtE25/rlggjBYYNd9aIVKDLsIfPVlfAbzBBb4JYQ6K
jVz6JkVDOHksiFs3zDbTD+1AImTGKEcfbVR0MhtAsefjYbGgfl4MUIeWvWqIbRZUG5cuZlp0NU+M
AU4KHo7U9xscJd5HkI3Lx+dtaJaP/RJdMzxbGBJwg6Bn/bztWcBdNZu+NY5e3tJVmM0C5p2SDWH0
Ogl73Fojum5STkikBQTnrN+QsGICF77iJ9n0fJEhSWfOPeAWd/8o8JixGaNdKaDch13AQlkiTCeM
VCgFwhEhXyRstSUY06SM1h2z0957NEAGSTsD0LRdQMdj0h91LiB740Erp4iN2apvDhnmwhQZTHa0
1FbAV6geDo57vEBo2O5MihsevpLNKpiK3hYSZMOkQJQmE/kkvrlTLU6sfGCIG1KzZuE9Ope0js3k
eYG1lkmffqysZxbWd9QEO54e8XboDjvh6Bwcc0PiT1gKzGrbUpuINKPq3DkS/UFKJzVvksDfWpdm
XaYGiMbJ/fieOsiSAXYYnftZo9c01vUlaYjK7SjYjILHgtQxo5MPqy2aIZTtdxR33HI2zPLpc5mj
OrAwbauJ8W0E5AKG3WyW+Mq9OiYg13as71kJe5xMSPHNQ0q/MZ/K0Iyr0j9PC4vE93igKmKQhkS9
luC/gCzouxCPlrXRThKVmu2q34KLi0ynxU3dmbOSZvPE6msz/dXu9+44lZslz1WpxmqtsMFxVPsL
5srlFQwDK5RxAwlv6hzCmBM/GiuTMnbxayZ+3+fc+ljBmysKqSr/S0BwHVPYow/FzpguMGPnCfX9
ue2IJBmrvkFH/dtvBAgK+oe8d5gdkTFIKkdBDmGEv1eA3IacKKjZVHVeIO4kwPcOalqWMZ3ZrQK2
9g+rMN1U4GKMeOzsNgKjrNkeH6DNVUtMDRZhJmyOD75f3H0GJFlR6ED91wDeA5GFDZouX049PXub
u7v1aOGQ7w3tC6cFmuUbmeliQkIMy4GbNB2yjQ38bwZLgM1TVeufws4pAHDkDXX8Xvwk56QEL+tO
8VkSCmG963cV3qvlq5uQneXYaF+BQq9G2U5DUWYXKArm5XsVfGQjCKBaf+MWU5EUDD2R68G1cL3r
Do863vIWzIREDUDI/a2JMFAaiQPCZ0YohGz1U/2lDCuXBN+KAn6QmgqUBTi/w+hO2qKPnJmHS/mq
iWK14d8gcYE1RfP20RiJTKlGTB+cEWc+LBmq4txacFE1OmvtO+39sh5vg76Od9dZ+LklfbUWTIOr
unk+6lX4Lr7rC3f/gEglmIzsNQoDJFjFnxENuhLdmr/JGYdoWwKdENSSlADOojyOy6gGszFOtFhc
HcUExI0VUst4oD/0SIrSl5K8gXQakmw+3SGxqhuZyma67GpgX3TR1hxP4agPRz3OV5rUTNOk1S+X
EUDEIwcarsuI5q9nj0fDV0Dk5jklGk7ErhzdIWCKH2yL5wJ3QwEcJaZywSbrt2aB/9veD1gYfV0Q
8kIVrrILIEUmJ0r27hhMoml6QE7D+mxW2cOh8M3jEpQcT3p2IR5nMPEm5PNgBAdvVugTI0om/eg+
YWhjjl1NVDlzG5Q5BW4x6YwnSl5r4MkPRbnZ20gL0Fw/NzflN+kJugfb9O5x/Xayti1Ctg3tCWvc
fIBoe/glpTqFgquliIMCVI8+/rai+5eZ9+PmvOyCIFw9LgF2n8QyHd7XQ1H15DokawjBJEKjdXJu
hpcifeF9QvmlEYLOsjvsJIZez6Qu+DEMqDe1Evh2zvwlLkHfljIAu4kQaB2Eb62tkxfFCsAgpbpS
omk2fZBKeppzerNzxYv7P42r0CuTbpDNG/lZlf7R9H9udmtrxAde02r1euH4Paih8UCLlvqm3ZU2
Fqjqbg+YkETZogJ2o9pK2i7yPOiJb0xcbAmId3zRgNmxnGK4N381yhzWQoMBXUb39Q3c7F1c4qAU
gMgzkAMiuqGx1e2qCHed1z8ErfX8E2C5NGeo3CkzSIuqfrwM23vnIwaqckdWkdEQNY5GZVh+5oEI
lYsOKKyJUoRuYbe4eXOeGI8K23Ks8aTAZqoaTrh9E+8y1hQdoejQ51o+HdSJXKLoe2LpNzNiD+Ks
3A7Ga5Zt/lKjSnrurTN+gvkh14ms1sqOP9IAkzDNzWNP57dCPpGMU/xDRACHGoYgmKzNptMJWbe9
yyspdfPRuiciJj1uPPZPrFcdbCANDPHNklE/tT59KwMkLJevexT5ADGF+AQPT3pbjafXkNo4xIem
CFJpOsiJZOzLgcPiIsj4z/GvhiNM7cUCsb0mpzyQsaKm0UVbVThwv7UxeNvaOCX1fhXKjRolON1J
kfzV1OeyvXmIoEYTe93ilPujnbnighnX/AjCQFyCcMHL4EQXm5g96tlXxlu1UeojMWdkHNfpe6X7
tOy+sG3GgIjdzDJ+SzY9SvVKcHRt4cI0weyZPV6o2Ven9XcYQkG2nei29JJQTNMgFIETiQlO/M4T
IoYdtxaRxHDyg5V0MPGD32DKOtJ8ljwFaDVsOCHEHAIZGEYlqSnBMePD06r6ZfKu5VS8WBl9laL0
9OGg7fXoAq8h54FrKBDIHZSdfWtHA1Hax7pu5TDxI6AASo9CEUmclKlbcl79OorKBscCSehMfXSg
Wej15m/Ct1GoYIBM4X8FtI0wVReXOluDdkbTeyX9aaXhVDXDQnzGD3fgHl2ZOcQJI3TwikD2fsDy
MhCPa6sDwHKPrQEzSetoKDDuYl6yLpb8avJLwCCdeJ9Oy8fNSuDzKyBjvTyjHmSNIFG6jDkGv383
UweyMgSNC0ll34b9CLMdvIXcfm6bzPundOXkTrj2PfFtaPT/rHTj52c61mjFyWyVwRH8iCXtTnJc
Ww0+Fz2zIi52l4eIVyR9BE3tu4GNjHIdnG2Wa19w/yC/vre8lLAPuDw2LzJuw6bzGUeXIlSEFq4b
t2Kec9OKZMdLBiFLHiHuaslSF2Mx3c7unxlzFjqLubPGWo88WXhl+ZRFEXiR/C0b/3BMqehxUrZ/
rl2/h0XLZqwmMjn8d3RGo3ZAFaEfRJPgd8QufHGpVe4cdf4FfonlmRQkFGIZxW6TFt+thzMB3/Ol
tnOV7UaNMdO83zdoeEPf96klRV9OTTdLARW2C0AMbrKH/WMjpHiDa3zWDvXKARwEoWu+27fK2P1r
heEBgAdpaORLlNum9n2+H90vw8uFAmMUZMuG6QGRQRXRBYWyeacBMx2OJxvvnPrnwZVB+aJpZS7D
j7xpPX27fbX7vx1FuJD3J55UcEOMgcKYM+QUW+HKpz9x4Qpufznm1yS78wnbyjg1Yt/fiyYR5uHK
WlI9dx22K2TSbmwy286x9BlrMDK0LZvZ/rgAMnY3gICpeimkwjD+MaDcnl/r+H9FyFtdNaeBsIR3
nqTvksQSLzpmpALfgxeASaY99n05F9mfbpUX4Yo1+fVFbMqxXZSgxSX/WpEHfUtzewbrBjW89f7I
PNNtdRirxNPuEXYmIWTI1KWMcLd6p59Dni4zvpfrBlNTeBvDHjaQgAi9dEf2Chs5UqhQDVF7F2zw
oeOCx6NEFo0Kkt1L7OxU9miYQuorOUUr7loAZk97sNi38+LHvzIzCeaxItmO9iy/rfdwThpKItm4
cPdPg+CM5o+1S592J37GHcWd/18Os2T44luWvFEyVnRwCG3UdVO+eni43e1Rj96ljtMMklUhpe4g
AtWgEAUUvNGDpaVDkX+mW6e0B//yWc/AoEOBxbZmJBpjXMDvzpuzo2F2Q/+bWlG/vOhWRPuZMp4l
SHq5NCB2zRaq0HWDH9Hz7KSsFGjMR0KT5HWbKEf99we7ezkFAyywVGTJluPg68JWYruZMlv42cnS
vnqDW9X7s0RGHANLZzyHdIJ2YBthGFwfOc20yyBUPqItuOFVx5OUdBFmVc+A0p7ayPdXc+grkKac
Ke4KU4m67d/V3ueQRB5GPut/0ntxaawKNSVYp2rFKPE2vei0ucH5qg938or4hsa29EJczrrEZpVx
J3KrFULDQN+gEq1+ohk6m3Xio6gzmDX17CKJgvL2LXnoHTHpX7MlX75KKVH8usl05FQmb1XO1Whp
/IL4UA1elGIGxcxGDvxsgRVgdeimbfFG1Qx5hSmuQaEgxF+6y2oucEAVdrg4B2LOpUslFIel0BP+
Z1fp2/4JCcu2oY6mIVHKk2zmIVaCCD1XLgEhxjNzxRDESRqwKAha3LQlw+6CJkyuvDJtumYhdSsO
VEJHCJhcb1+7sPtk1ohS5pcKKwMA+F6NwiXMM12hsXacfoqKr266U0tElvxvQYljcn0mwdq5s1i2
oqYgDTCP8bfc/u2POWZm4IJcGYh788F2XfqqGB63mYGqJjjYrzghSgFDFJDjYDF52qYVW/9Y5utV
hu5nONp3GvEPq+IsC0FQakjexy9Sljyw/ENxe6u61YbSQZWLyJwaRQ3ZunolnF4etyvI88PQ183Z
hpTdvKAktuHtaSdbVO5CFZsg/GUvatW0glYU3mTbk6AUyzfVSlggesTGH5EZLx3zYDCAzYCjQ3QA
59x/bEA7Bk4kf6VbDtxxi3RK9of42rxVADnARVeaHhnr84mpkltiNLxJF2huK2GeXtZy2D+hD6E9
EGHFhA6BaylBxMYpso1/DvjCWVm4BFW16WE4go579Gn5owptZnZO+q1PVLsMiUB9tVN/Y7lCLBtc
08zOy4vZA30rJRk5eeVJbxhTuRSyYXQB3+38oZV0szUyzWBizRC6BEpdlMx5/ugA0J4LPtF+p4Iy
jJzG3ZQRUP3SOwriTUMrCO/VtqbC2ZWo8dW7CAxa1e1yHP3PhE0E7DS4rPhBKeMpTDweWAvj4qu8
UYU5tpKWAVMFLNprIIyhoWOAgOPa/f47G4HKN5Kfuvr8hzwabqrcM+MFGc3Fy7clwvZh6dgX1rkP
/rlTQKadgHk5G61iNap6YweJD9UbZHkGHbFfhoXZr27g8k9xW4wlEFNQzHrQOmdoKOK1U5yrBDm3
GX4SaOqTWD7gKErL4WH42mwlBbDYXUV9j515eSEmYeemHJKVIhmzuo/1smDLkVZCRbhZjIpBhd2B
aXe92R0EOFPuPEnLNVTdS0hiGt0BwhPTzCQoC0SAhfnliGs/qJT8IlJKwOBpSB4JPbXofTk0qpWP
4N3ZMC8zWk8DSiOC38m0DN4+lgZ4ILDeCYCcs3C85jHEAeYlqDEn6NrSgrRJT1nPNj8DiUuS9S2E
/MZM7k6Op3YrkvaLOonD8yHFZ9N0c6M+la83jqGtsBRS//0fhtWfi1d4EVI49ERxQUa2aWoc+RoW
n/OCKof7cC9na4UttjCAsJBEcXeYIsojQ18lZryvZc6buWlNSQejCcxYYVrGB+SV5Bop+q9jMXKc
5Ot/TjViyrt3Nqcfnh6zJvqsBP3QLTKK0Ocl/jzcp6mc69wfVM159550bfr0CA3dbaU8GsVCyyvu
8qcGQyqdTR6Npo4gJujbcgup8Ee80QIB6Jrfe1DK3xGohnYUvVPWDAqGEjQxguGLDSdjkLvrtVv0
qfxCoVpRc5lt0/dmn+JX+H4iZW4328L4y8kXiDZC71LuRFtFEr8sB3Xknm2worg6UeMjtyCyaeLb
vg5PRBk96km9WdaOP5qYZEum07cqNLLtOnkbVbU3j4/VSfbyCqJMeA52kQnzvhRipgyldYgTh4mj
ekIALllvFNaSZPQo74EIIMm514otulo+eqgmmOtzkWI0hI/BU1sClRU1reNuiWypkylPdVMKotV6
p9BUmr6VcYXxFBnCC4qfpHU1DxJrn21uRxOyh921dfva8TTo+8KvCmYZ+4AqD6X7WnF+c419q05h
saYKCKEwUqnm57HDRWpPzzIfc66KSCHuUjXuiby5zgsxgbhtvll0AMU4EPUP2Iaxuj042TGNJSk/
QDzZu1fTKj5gznj0PGZ6XJ6FhGkgX2H3+3MEYlC9nZxl2r10W8EdQfoGKOAv54p4uCXgqrXj3rpw
kIuQVkCwnXtxuxqUwyEjeZj1jsxj0Yje7dogxmAh3AEQcn5iOGpif4Umh874KGXl+JwNZeLhXoMy
F72MnMtQX4MSgHN+1L8r2sQs1D3R1TKAlxVqN1oVbyvK0uHsFZdsKGDfiSEwOEx+2a/Hy/FcxUsi
TiW3lHwHhm72Mh3yOexvmDS7x0XBkSiVar4oOTRvDWkFyWpeT+62H3p3IaXgNLo66fLCUB1L7e/G
ghoqWjydbRw/dTsdPz41Nhkvk0jZx8iwzrVBhq2gjJTP1TEbsCCcH6T0w2zqOD75fayg9d3kkA3f
KphldWjHzwvJvxrKGZBNBQ4I1kDChRyBZkkI7xzTa+JOokfAfoqUM/vp5OnUbJvmILA7Kp7JWpwz
HokCHxBXD+YUawFLfXfeeb/RvPVMZkTNMEcvmb0cB6xEvP7i1CaWCTD1pVWXkQPmk0c/OyWXgnH2
VKzCL+2Uo2tLdXfXyYSvnieXGCrUDAJaBLCa4x9VHL4OeUIs4L/fG302UKqXEXdStgxVTDmkKBDB
roej0C219YuipF2xcjn9t7geOuztKTWKJvvvdvWq+d0FtJKGXGtnFvxtassg7NhNQRb/i/pORTMm
y4k4D4w8+jZXi2wCTaOPtFJs/mhj/W8qFdsO9J833X3WwAFVFkoMmhs1MoYL2/i+Vb7k2LU9hyXJ
4dTnP4jaxIZnIlgU0yodjwaiFsEujrnedl/PxH5Px5QYeHkuOVTHsFwTxp/hs3z0me3o18NsGEmi
mPaFlS7K92H/5g+3scOioGWOpbhvuaNAnQYl7hzl2X5DZlIi7YbK23vDSNy0jRLXx7EmLp1KrDw2
3WsOnF6uLc8mQtHuRuRgI8AHX73cONd/IH6/XwHJpe+3bRdn7gTt9SA1GLM1jHFhs7nkdNefdPPt
qc/4hbfCnBgVD8FofZUP1vAtwIYEMhAzS4fwMmstWY/VkRmNR4SGFCoMhu+IEGPbOdsOFY57y7v5
uu35kMeTr4MpDnann/AHFR6ZVINFp2VbdkjX/ZPQAprcWaOvxcHWcUsvOB/QuQApC1GTUpHdpgGP
7TQynRHxVpiXbCLJnaPgoxbrojAn5l4p63G53i89OEp2enPzVymnNOGh0ACaep+3U3a+azHbcc0S
qrrtcrzjFYJroeH9H7Mvk/IycclVGQ+1A3UuDdgPnnSLzZJa4PfTBD4ZDizdGJLkLF3LI+rtEApE
+9/fVkTXKnBHHeCjB5gp4Qw+Dr1JM9zZjM7X71X+eL9FxHynhtCTtavnmHiTvis99I4NlXvX1AWm
Bt0LRvld5XRMFJmYx8UfgrtYZSJSAzAf+GZDdL7yaLtzzmP4W2eRnY/O0kuqRvmrAJmPWbaNmg0C
yUAO+vcgsSDZfvQEZBLGMeplo/EtcHtHX9WqRv/oM0Q2AL2iJ1g3fEZ69WjTAUT5n564tZBYgGyw
IFnM91t0mMqUbHdrB/SINgDkZ4vcBK2W0iysDJ7knQVQLonNpatu6yb4DJmjbiUSid892nZHvXRU
ByVBQw5LKmr4mQ5t6VB7N3WjD5/FwLQDo+OZo3DYO9N4ZCFkbel1P7EVhCeIRIE3/SuAknvQvuyf
L0tEZ3bwqPXwFjFGhscrKfxy37mAkTrQltcWEsdGwIQWzF+tq/b+JSIR+X2qtq3jiGfHfz+R5nSC
iGR/ZmJYuJXgwxUkGZBJ0hQAnoaNhYL0SNCp01u7+UJjKNfh8B+ZDVG4IwdLUQbPE5GjsCFPJixk
XgC5ztjeRNWXs/Dbb2oSnTwtNeLZbJALpAGoP5dvqyJnVL60y3GMVgf6/Z5u9VwsonkZCA1uf/Xe
FB5na+BexkQQkQq+B7DdSOq1cykeZq2lV/ezwtbvbQ9tez7gQ3oFALt6Zmmc6QxTLkPlespD1nif
G8wVnnsBx0fL/LLTbC9k/6SIxEk9bu0T2qqo6UovdahxEsrZFAyMiGB9zzhq3tDoINEytykKUO/y
WlM76v7FLhDCNPKj5A+KP3ZtGzOmcSssNsLGTAExhZqHyponVOpO/6VHQtKs0QKcLsTE8pIBQP19
TEFVjtzIiItsCNZhMdHAj0h6ttXH0NRFQ39Afymt/XG0dsP/assMHf16ort/9SWp54BVI3NJdtXl
gRHRiyQSBmKhNQmVcuCBJjMKhDUDhirX4K6t+njQkgSNwLxqeOkOUgvtne0qXeRmO+EBE02e8vuI
0iZtLw+XLxShmFrruQ45X6H4wUDueKpycM+CdXsuoCbJd20qNkhp8VaRCuPQUPU/PB6/WBPwS+/a
WJYp0qo7WbaZ2SdWWb8Fgz0wQECeO8IJWXLmxASzON9/gt/PBONCXBevo/4oZIMEYW4TpF+rjw5h
v4pxAOjdgJGSAhSoz1875JZzUQKkliA32R7INeOVJHNEwgEnKRYah9EOGtsOPjiGqn3nbrX7K96u
znaF7k7cKWrf+kv4L2wVSrUDNUkNo5QkNHR1H4nW3Qs+rQ/Y9CEKo3BzcR5fufzJ7XDZvRQ4JRUn
AS/aVRjUxjpGec4+cCyl4PwyHenteUjZUYbB8hIfXSzgQW0ji5pVpKVf8gl05yY5MsXS6Z8p0N4K
RT8kChIbe0UO2gsO+kDJ1Xc/+Kcb4pnpA8GVmptSwuL5F5oKIFHyNMDuhBA8Txh0RszNrNqM+QZE
1iHQ4AgVHPtIUbOyZ/mZJow8UJrN3BoLhfkxv0jpryfa4GDDOAS3psBQeJyH1dxk2Z1BDVDJxLeA
wKKyQ3EZ9OMeMzvKi8qtZkWs9FaVv8L6elGPEHl9W5/un8kHWuT6akNPsLxeGGbTxNAWf7rhP3ME
a0PmpEiOElOlKt8eJozLnHQVeF0vDG4iS54OfHN2e74QTChk7qkSBKXHFSAWrbuI8aCIWyBA7ye3
YyK9wlHfWQFON/JolqqxJsAZWPj4+rt1u1LLbOzSJGt0ZC2XKlK102zvgyPzlH2k31gFFF8A/u45
rqGT7j6a4llzNJ2lGDWY08ELSelsvsoN1kH/P0bAVA+L1QFxcvgTL/byYsuo3dgODGvLtwJr+zTN
4xvNwtTDXLoydT1Z3CfAJJzYl6U/GuInh11GOIa2MyA/pwu8yYL90rgjoL3M3Yag452fxBLJlxxM
CdEumiMDLDOrsqdQG+4bHnV9Lj+M2pmBzwYe0TW49zYj/VsTg9Okl0ZqlhAMkyDlfxGXIkzKIZZv
rLVh4gqoiNfnE5xull4BQ4fJOkW+FbjcjKXZKo5l1Pc0WyF6OHnPptQhxtCLwrw/1EHBl1Az/KEM
ULDRVonjZAy5xYJQSOmjAuy/BBUYbYilNcYWlwbornZhbY6GGnKeqSVQGLsyCNGfnlKCE/sqiZt7
jY0McOf3XnXWLnI0g23RqhAs8w7gJyQa0uysRSy7uWcYw2Wj7hTlfFnDsyPwrNJMKQEnOe5mmn+D
wsN1YdCCIXHQC2p40f3KTXvyhP8EnPro6HkL/WBhRVEGfjDC+XwKv4S5mZL6taIzWsWqPmnR4JJx
674vIGshbKBGzwRXOJyglWoJdsjXcLgD/ZnjhvH6IeFtzijFR0wZeA+Q3lqbagjnsCIZYDJ6za4S
qJTWrUW1BnnBfm4KEgVEna11C9c2eMqI1PKadlbgvYlprbItA5lz+qtAORPcODIO0N/NB+Hlu+A1
aXcgZMegkGvoElzdeiPN9qIZaHSfhahx4kouuE6pfNl1kb1VQw04A5OPgpHIePNIeT1mlA4fbMIJ
XBXyK6bs6V6LAhoHmSvjH/98zRBxJb2fFl6t/UZ7tC8G2bIRdMtQzFcC7ocv9yMMp5M9bExyjJZW
bIbe2r8u+2MQdt4RI5cCQ3gxomUiiW3qzGFf5aQC6UBwEFjEj+WCdw4iuOhXyNcMjUhnpwcTf+lI
vjon0dWoXFwS4kDDYzPfQkTN7yg9sKaisEUuW+1uw7H157P5Tf2oTgwFYTeUIGBIZ4Bury9UX8Ww
cJxnN9tqqYiQkAfqhp7DQnYywfxAs25C7rV9LYOn9OXgp0F8skmTXbEOKlx7hEP2On1ZqYqtYziU
XcBfUYBaPEf8eHHLhzroZE2AdBkSJ2/ALcuFDjmOigrpjZgdAZM0aJRXVGpT16WobtPjDfmh3F7p
4gJEhZ8bdz/CIcJjBwEizkVUmkTDXYe9MLMor1Jq98uGB/PiWom5Km/VO/rq5Q+5mCDXNgJNlfhQ
KM62miVGfKtQX0QyeIZhsi5e5B/X/i1k7RTucKLmFuJhuRSCZKEAXPJQkQU2MmC9+Dc8MM7ycu7Y
daLwAiKKnwVDtG+vhBRpdrXg4mP+ZVqog5vmuJ4DTPuypbXO/lqQx8HhE/d4dwOWJOecz0U8Q+X1
oa7syCXFthrto+SXWVFpBcLMP+N0dFb3rU5cowzSkoT2bpo+CJBWCkCtOISsEqqrNpH3t+uPTzf9
JHomaHDfkhrqrPFH8Hzm6dRyeI9Nao1cHMoWnDsm79d+tVjGNx73JgHD74lH9NT5Q5u+0IQwZTu3
+n6jNuCpIKuoO+PkF9QLEEhH/A+7Qfx1Y4E252qKCU0HXT9CtXmU8rb3235IiOl5gUIBV7okZ23C
N7Xr9YsXYHpb4clKJnkXwBSiz7fwkqYKSgzFN/DWcoeUpeqwYHXIjvyF5Jly+MziXpZ+kyGSLRVX
a+6wwDAsR0RHSAWYz/rW3z1jJKWAsFyiiM5ZmxIPKCnODbSw2+7Nz12LaQbw65Py8efS7hj0Rh5O
FGWpM97ukF6iW3tEWogRMA10eq4BYma+1qrC3lZL2SSxwS7yp40whNxjqMhcmJpR/1Fnut2REFxe
6XawRzkcKMIn4aecErfa0YyWiBWGLzS3rAo9X4Wnkzh4t7wiHiy649CdRwVVhbR+QEakIS1NLo4z
1/x5xX5AWsPiQrplIMRQABYPTX5RalJdYBJdZ03JSgGNRFT8Lm68UNs3of64n2uU9M6+jyqHRDyi
pj7w5lwTUkAhYT0VsKYRf4vtFCsiDyZwdEqg1nl+xPUvoicx2BFF/Cj4fXocw3LxmIULj1a5/TqS
WFNim3z1aMn3KvVr5c3Sa57YdnNn0lFIn8HfUZSb5Si5O5jv/uOEJId5CLlMKv/zLrv58ApSQBIn
yaYxcrEdkqcGkgASk8Rt2svGgK+lnA0xFF7QM4CYYeQVwB4p8dK0zj8Bd1Cg4zFKtkQFJweNo7Z2
eV5E7jb8Y5WnsE0kQmPMEPgv2dEcEkPqO55BD/k3ijXdvLgbq0pjAU6RWIeoeiIgNAgUC66MPlk1
WiC+zBX0eSnipmgGNpPKTO8xSvTqlmcSNo2oIXPMcMZEhDmCyW+4+Cv2NvjWNLbDKtTVVaHzuCdY
jhZLT7MoYWumydgA5Sm7I9/PG9ZY+GbEeG9h/aAsWYZNTGzv1zzQsDoRG1l8lrWz5tIBv6d3NUwz
3OoTNldsYOqsWLb5bCs9SRwz3wjHzDW9cRaBCtj3ceEFJ0+RQbMBnnVKgUV2GZ5Xk50sj1JNPJWL
8r3vP6bZamdudFenYZyTuliBIMSHYVRzNMKOTvK94z0oQ8lhbbk9cnEedmEwBtbkcuVHPzN3ED68
je+U5tLFFb5IzctLO4CdpZTGztD9JJadpDxcbJyGzK0NTEUDz023rixqWtZCNf+nSRo7xLWYCz0i
0Lc4l4zHHPpl8INA/LcQ4tJGN1rzO+cBxi2MduKtSKj5MvVNshc1DRS0m5QNrT8FePD46IVuhNNb
frHarHKnOPIvI0BlHBR+SolDpwHSY6kWz+PRGFnmsYDI6SSYwYbzn+UigA/tzOGYMa96cVmW9CB3
5m8HiJkXAQ+jFzc73xylR0LV7ceYq9xftb4r0v0lbzvU3AbN5Ooyt2uNZcFK+DgTTFH9D+KgzheM
V0botO3mV0GZrPheGjS3PUOB0G2qWJjlDuNUJis2FeDzc54kKQQpb1Id4AN1fxy8vXE3SUQ1ULBh
PPDS9K6dTtTjKRjAolB2oxTHdZAPnX55zT6yJ92AdjUXYPa5nK9CAoiXXWRWmO+T374+xUQCZH4T
6dBX7bxKH9JcQ9dcR8XHa1rpdUqbuDShlKzFELFXCKDDmri5HzUv/FsEpYficpOBMQPV+S3v+SlG
6aKkBLC02TWqMvKTNMpt/URYdk0wl3+321/W+pAxDcsBsomVSxzMKYpfb9V8lj5pwYODwKZ96Gqa
mnFkpWvbyPeLzjbfPIlCMax0OO9GPTAmXvlQldQkjCeLdTJ3FU01UJC9/64ACExPN7dcq5b6ijk2
dix1jDndboLTheZqBfj4jnolv78Z7M2Mz0Mq8IkQq7w7W4/ZVnADlZBhevYJdAMkfnDYh0ZFD0uk
FZJqnG3A2imqqBxhKehi/1XjlaeTun5OfN3a7DA+7VTFot4IrmIQdGPZo/9Yz2Op4N5ywzp+KScR
3hZyD4H+gxw2Mqk7LptllF1bm3040Pdnv5kLrHLprMUk2ovaKUgrmrXpWkKyjwNP/yOGpBTTaK96
O8vBFZOX4ZusM3elYhsOygCj520ShdlGMPINnqpMpbMWdEZ5Os2MK6LyvLt3eMuf0ZSAJFaVM27o
CDrNTM2UnQ/U1uF9hv7SsxJdZtHopTZMRiyHw3B593F8WD/NR+mg1BwBQ6DfwxXyJaj8kIY0Sqzx
pzC1SUh7H2ja3SROXqZ3xmUwOB1myF8dvkmdGcDY1OhBHWA2/kvsG1G+RbggrOEKRu7Wvn8+wNI+
6XNO9ztYPNj+4+7Vg2iaDLqddgf2j6gqV2zap36RSf8dm5ltDmjkXG6nCzI+xDaHI5sa9wv0A7nJ
CS6eeQVXpAyIgBTaUawmMO+EZEcW8gCm7bUEY50T//4f3TNeFhXEXfJon431326wxSidqemZymbL
emdsL1EVrZe4VIuSSAFO4fFrUV6DK+zO2Tyvy945jQ7qirMoP9lZOHAJ3PNysSOl3Qcb2buV9Nw2
yyBPATACagdmuVYf6LYtf6vmgIRjhCguZp3umOiW6iGGorRsX5A6yt52ZSSFo20bQbW8YHqmR5zm
rtELjtTLqI7U8025vrbhhzcWgx5t62QjsKzZLHGbcXYr111ymtcdIE4J0IW8y8/2OacdwrBck0d1
Z0uEqbQjr9tImcttnvSfZ246atpzX8kfH5/iJULC9Vdg+YYxt0nNJ7aDC0g0xeo3EWgGaGq8eIVV
iz7831/B4gF8VIINd7wzRbA0bCoeBt6YtmG8gQvZLqyeWGOjSZsw0miu3QOdDylkPHmuFJyL5m8q
hztoOPEk01dYzpr/WL0zIf2rBqrJLH4NVHvifa4HV824j8Y/SH/pxnG/1UjATVdrpNhmg61SzXb+
AzxrbzVbUUYZ1ru4fhjrsUalUd0kZRwmX/rpMFdlOS3eZQ/SYHoZ85/z+kHIsPSZlzFlEnlKxQF+
1nEKQknGjNL3TNoYL7H5HF+7lMIS3q2S/6XstyJEeDyg+92T45IrGMl4B+ZOToaK4vmM/DGNYZiY
zC2knSS2Vd1m0tIZfENzr2IQwZM09vdram7Ci4ZuWrE6CnlKfJQzfmipnMWJirbslv7WCfkANcDi
B07YVqN7ElOr8mUqZ9CCwMs4/8GWn9TpEn6wzERq5tkA/AiAZGjohVLX2MJQDw56d4IvFOEcQUpN
YCFrkaVn0U1QN3eCs9eSe0dnDo0mI6I/MW/XBD3Q/SaUguc4U92LfKJp+rBv8Zbtw9/yJTrrhopH
yZ4j/V0CloEkOXIdgKfeOFPtVfNarMqYaI/R/omHh9X/79jEfVVe1NiGNh0GK6q7cMVY0yLMIg5B
Evd2DshQkhTQAsV/y5M68qGXC764SHUqeBINEvZl7rqOHFOn5PJAC5lkr63XLyaJs1DXFwrmdiaf
nGxu6OaO3L5dzwY5QRVn0KXSRr/C33KbA3fD+ZfOO8GyQsowMZ0N4UAJGA4KeHMqnFlKOtQ+ZRgV
wgpQDpIoc/dSMQvmzQW8yJlQuhrwrpPOUpB7WaPGbhSITbzGVPpLlk46cqibl2GRC7OiiFDIRUYT
7Xf/AN1b+qKvgepdJFDgM6ujTv4yvEMY6KmTaQ1wxwuiGW/5OqBlO2XM2qOGxSayxw8BONa08dkg
SeL20GM2g+H1o35TDgnKxe5qVeorMe86cRSJIEMOG+Bi9k+ef3n7bmlInSPSWUzblzlvP0xD0edF
On+LRFjHSz5oGoBEP/vuVbMPz4/1Sw37h8MBk1z5bWodB06uyv1XQn1WQNqfgVP5RnVglhO7zw7l
eh8PYvm/tuoh8DVJMkyc04BeBxyEpjCs7l3to2kkqu6OWAJoBV31JSH26br9NzyznOrivp5plUwx
bU7KEJL6X3d22hhIPALF1vPTjxcegkEq5cgTEuX8mO/WMA/2QZ1otBF+KSMMiJLzZVaaUiad5NTN
KMqnlUysBvMEg7X9fxzm3372jA6mvkxU7hsGV10T995uAuWXJXJ8np8QXQ0eIETHN6D9MAbCgWFh
MTyHEtj0/Ef2B4F/M+5zSZ/Q4VQ4LghkElc0dXtjW0KA5VKRIDV5goZrBESQVWuZpBrgOCQrDLc/
GeZbQTZnL0FC4AhTZbYhAe7wG0x0G591xPF3eJ1L+IYf2AY0MCVgkb5CkcxD7F1FsNZtwCNGBgm6
3kp+HQqd7ksdOozSCJfpK/zAfdt8Wfyu5n9vZbXDlD0FHglxvCDsIH4YxSNF+mC3pfm+IsblM4aE
PmyfIVPqNe4C0skgIHka51ps6WvMwe2iEO1+mA9BP2y42zVe1NshutwQ4VoTT7JPwJJLU72DLG+W
p8LS02+M3qU6C/qBNwZljWIYVXMUlxhD8iqiizuOM2tdJkppdb5ilgyFVqKPdtHW1DYG3UjEeJMC
arxOjgxij76YP0PxCbnkyaD4ECS9cXKPJBgXB3pmiTgcQaoTjrq6GIJZlCklTgHs6Wh8KMct/nNE
0LGMBg/ybdaMit0deTniecRO8jBjNE9LoLoOEblaZYh9x9bt6MvMO7BL5lplz+2lUgaGOmI+VsRy
Oe47JAaR0IMY6K3+Q/uw8PzFd4orkYSJa7pHlAjgiWSyLomu6DbIvZoA82zgi2k/6Fza6itTKeL/
afdEXnSg7csuR7LkMzFkR07nJdWebdXVvhYv3tAV8d/WVZRrA+/kvCdSe7DIXxr4JNOU/tYO2NrQ
zEuYob2wutoiWQX3I2tNFvSOBknW/59uHtsM3GiNuyeJSPrOb4P+yc6qrFWo8O3sFC/DjWPkKlAR
gemBC8Mru53C13ZzxCnz5+sA2rPSt9xQr9sRRKN34mJgTTLXHjhF8rqRsmK3fM5UXC11QOfEHSWC
MnC5gm1caYztQRNFLyF4AXT+EIOOhNalePn23P36gsDlZnpwAbdv/83dyN3eyGPTXkL97vl0t0YQ
m+Wuk9uap9kvA5CfijSOJTxP9nI1suyvH6llZj7kzk1slL9wf2OfVlhU/aMeaoY3zPhxGzFmTrlL
TOAheJqtOlyR2V8RTKyr1yKnJAEowvBkOczQhp/mppsXZ+dnbpC/ttK9F2ZZkZLpYTUd2aZwLeKQ
eiDzEzl1oHO/NjnXb+ffSe9Whx3C/u7TDZpQJNmyGRSdF5JK7ic2/hUNMnf/6RE9V4NVuaa/NVun
yUVEHM2byqVOKHsOgVNbtFxGoYkt01ik1pnyNodQF7pFcmkmS3tWzr0MCpqVOBbZnewa3aXtoG+k
JeWzSg4ofCaSskVHg1H4rLkTVaOw5v+AjT6w6QhhBdqLGOSz6WsotR3yQvB9Uc3GSCfdxix1gSZt
W7QFdcGlREVWkZU30+rTEYIWbhpUxkW1Svh15+5oIjv2u2yyLhqyPH2UEXciXo7q3b6CDGM9MyGc
wTKZ8BZ9oo04Q4rJeSSk6PPvKB5MceecEt3RjxD+XRHqZ7CxElS51BlXfS7rbLpANX5TdhOSpEWq
RuEcRmbc9vjOND9qBTTT6JltCEdo4MMwrN2wuk4HZVWgSict7Tve57LdGuYyENlrghu53VIZbwsX
h5MywGLWZTcXaxtQjXMQCq3ydHjwBBX5J6/KsA56qav25B8oMq2GfDnIcNymUhzPbFBGX9j7gWBq
GBRYRUl2WQ9Ls3vCtrwnQVS+F4IDI2E0xczH0bedlI5SHJrKQCWYXjWNXtc6BPIxv17/UBYgT8KE
Dnw3wvwSs26i0b6PtcLjWasMYFZl85fXc6BQrGbvwElJ3TtmGvojkl9v2ONpyOBL4EBUFkRgJAI8
uv1WUabh2uYbKRIKu61JB6TLztuSaKh1eZ2m2WQeLBmbkAjIpjoNj+ynyWdsYvK/8Lw1i0q8b1AP
l4IV92OtWfB8k+ugywwyPBH1FQPMebNiHVnuwp6gsiaAFow7EBPztFSSU45XBxyoiNd0YHCLQODl
sxdlpLBZ7BlhqtOF013RNTgWNy/bh8EOAXb64NkAWOKNy9N9uwZmtR7RN7ym5yqg0jzbIzx5+K8l
9xYy93BiJN0tfC4D6hs69fmZr0Rpg9vMNfZcp8vTMjCLbEHhdf5vIJPSpH4HuvBHNLqhLXHA8UQG
d6ZM7cke6nrd4n16L5c+BSbJ75PZ56P03WFONi1g0bydP6TSjRN4AN79w5St4Eza9BRduHeOHnQc
Nn4nHK7MfPN2+3X87387JsUVmvjry+Nw1jmqXRNNFj42djLeaF16w4VcI9+v7EWvi+q5k91cVTRf
QoRFMx674WZRUe65QgNqJLCwZmAj1hcPzWGiuAtzU1/1cjBGSGIFDRMeV7fbxqd/6sL1Db4agnRm
nnKlZU56lbrfqzGFux7sW1TxoWSWZqE+j5kPqRqPUEaFA9VIzcL+iP0B4wSFn2VUH7QpYqDu7QrH
yfxE4/fb+C96ydd1CTTnyVyOn7BZWRcEi0fnakzL/cmARwvedrTwPLFXTfwwjTHOnjzgMAM7oeOd
drosxk7ArTI5VVluGEFK0GSSABBVpBZZdqR5Xv9RIVvgg7t58CYTX/EaOxICBWhGbCMB3tYkd2mm
6lWctKVle8VLYVse5F5PJnHAdc4wVeN6zJaMC8dMKJmVXfp2rychRlrgvXDzS5dJqml9SPAzNKNQ
isM1v3jwZ7hLVVNSc7Nn9Qf6eBxkHlSmJwfyB97Tiiu/fWSQwyONUDuB5OVFXvnbYzIf625ZhcLO
tbRR6FnKMFQ8MwuvWV/DYETb0MEDJ1u36q+PBY6JKf2Wmq6Pr40nsb4Ur5uWHm86T/Lk7IRo4+H2
x9BynjNolPG+V07rrWNY8hTD9DNWrhb0rM0nb8Y1wYpLVb6Dx8ggR7/sOXVWjX2LWDE5fxUulvdY
r93MyP9xMbY2gfMWCbJO74eXNUFedlwEtQ0XQHCSRKBCO2mNggs3jquZDBZCzXZ7k42ycObOrcm0
XzWU5Rrmrrp+bDayOEpIe/mJzXPNmvNSo1BMTacbU+tE0cIo9unuSndsCP3KqTb27zLf2PDmG2Wn
IZZwDyhLvUEau61ufMqTvqlbyyu7Ij6D43TFpONxtHZ+gwcGRdm9hVmnDgvlyC19DjqAulWejg6O
GC3rlyuAdMkIQlvePck7ONfDZhOfQE6NhK2HSqlk37Wd1fm8h9AnIQKS/SZ0q6KftJ4DspuUihKK
H9mmWCtIC57oSlpE5cBRlw3ZClp3xSAPXC+B1CqVmv9MmmYGfG9wOTrRlVHhZ9D7kPgm0OTdIT5m
hruCq2KDydhnjvXaCXFtmdjh+a5gS+s/AP4nQv9S34IMdxGID7UWL29kaWLs9Pi5hAM9/87jMvFA
0vUCp9OX7dkqWg6OR0cbrGiPzKCH6NB3cvv7kkQDVG6wd6F+DDSlQaUUTVIOiY+e5enpb6ZRW2pk
d49g17Ew7nTU0cRx5cea2u2618Q2+MkY82/nfqYyMNucW0ku+vu8OTOvCjyxyYBeYt9BRWY7W4UY
IDtxuFrXpcyW9YRjT83ODLtmGF+yrtVTEWdezMYUByT69BHdVxPR7rf3UIYMrPnUpnxCtEUDowW1
op/ijt6pHjRQOR+5gN4Fxeh6uwzxepqFyRyFhmg4qyVNdL9S0A8mN0VnPb41XJ3lvrmLe5eLaNwR
YPJqXFtlONJty3JD+b2sntCiLnz6WemJt99tLs+ReYZtqoxkUJzIzlZ3nNuyyMsNknLXMvioKV1q
VZMd7CO7LKmEwX0qpV4prKieuhgCpz0g/0Q49wNHBmxtVTXjgHZrcVA2NCzKQsA2sBYw/n+3aFrK
Pj+FOerU3fYuYJkhNn9Q8tyFH0kk3WQ/2eXmMmW7tuk2NOiYvEzCgyI4dU5cSwuE4e+Nu+vl9rLQ
jvH5kql9VvZCTDVPCOnFupLto4Mvl2f+c/ZhYEWZVyMqimyVtgVwhpaASUcMGhWN5BvHbUoqc48z
gqxcfFydSajbB5v6eei4bbialPVPh/RsHRi5A67V60LolL1wm5izWa15dpDypcrfiXogUM9F103O
MSUcVj83YqDiUUKKZ2BzQcppEYKbhtN7qBIdsB1IP+FipvavwZeGLHDP1LBtrUvczy/n9K9ENKAg
x+ijOVVknJUqWiAv3oJMnxOrYbsrb/v0F215uJWCm3P0/pHEDGZnvi3XVljvmb/y26nuFIiVkobx
kMny/Yi4F84g+DsrnfTu67S6f26NTkPBPVnTeqLMPPRXwD2n/Wg2bCG+65XW4dQlTS1sZWQs21x2
c2FlviJEAxmPtsYWZA/AEWqzGln4gIIMiXWa6nAABW3ZpCNGu0Ly3DUE1VqNvHxg+AjUnFr/rW97
LOlpxBTRmeaqg3jDVMn5HHyHJrUJTLP+60IfE0SOVdK/wkyPgv9A5eHMyhZOPkfSkVwWPRnU/vyB
GaB9W9zr32Vh40Kc/APQp2pOGY5xO7zokSuXNa++QbbeZIxwPCyOH69pLi6JZmc41O0D67VdWPz9
RaBMjYBD+82FmPsQNru73VUYbm9B5510wes7sMGFknY2yt58mkN4zu6S7qGg5NXoNXQJONUkJpwU
6zPoWG/FWLuRAvsHkj8JVcCxbxQqRcPAxeIOyJNiwP3hAwSh6snkSaycOp4EDE+mTHBtLQB3ujoh
XltRiuShePF7kGPi/tXGooyrhhVVuqlV6oOtmqL0hvfDUOiULz0MFBxw46zxCWOeVtZkmhQJIkxJ
liX0CZFxjs7ZkVAeh8NdAAJFf3F5TlBOyt6bFiXZQ7ZCStQPG5Ns45bIIQCn1JONzda1/PX6pS54
MS5WkGgzQFFZ68ysFnxk7vEV0tptkNDWutMd7h1FD3GgRWDrIrHiynKr5PcgeIv+8FzOv0UePn8p
5w+gCLrEz3g/REbg+yLEgrLEWs4oc/zVETWhqXSnAV3hORfOZ6ZgIFmHzn70LgTHyBa0DshnVzxa
ttp3t1v10SiX/P1U+k5YqwmLlpO8hlQQNqug6n37XHDIGPKkF0SoIAIz5SQhsC24H8tETfI5gfl+
MEc4ZtPmyPh1NRILN/xVwBUw/3oS8csYkZaAk8du/K+KOfwE76U98Md8mqU5mlmWKaOkcikG2d8i
mPYKBFZMB0oWkVbxNNxSAXrPtBBLcQAtfaj05G2eSyyse7x110h2mtuFaJQESxWiD38RlYDDoEV1
cKzIJ+9RezqhRbKsOJ9VpZru2cFkmWiUj+rQIHJDIbCs2d5GkhnYFQ+HVgKxpX2NcKEROr7QdvRx
wRjpJ30xqT2NDm6cOyUe5HnR/oPHntr+6mPl5wYXDheGLyGs4kijhqXpQhpEHKDpB3kmXGNX5PuN
zlDuEA3vyCnNx3v6skSqIvSuqPA2wOAPZhdx0lVCXiJAnWbF+iBmzBLlp0I4SlCTtxWaMgY8UEb7
wKdUdCULaZMglbUi7EjuTR1OXq0bbXnSXRkQwsSqRshbr73jSDg52Arpm05MDnVYLclqCY9Qpcvr
jeYnd6MmheaPHizghnbPG0Kr9dpTy/A45vNfAWltSdX1e+I7Irk8f15HJMzFb2mjiU0vrUhMDTf+
PbQXpz0WEMTWmnAK37jhAg78nagJRV0r4xj0RiQNGwCDxCVR36exvbt82jBF5SVJoI1hDA2qc6eK
utBf6Yg+Ix8Oc7OPOoBvj2GIYK0ets8Zs6o70ORr9KrMZOHrY2mQm+i1G/rZRE2Dqlm8E62359fs
cDSeLWOx3OPCkwMmGtUN/95x3sSZ93z3/g8uvVErsOgask5xGQA0gdcYNMZ9D0rg2mRH5QuY+5SC
+gPC0Ce73/kPPoKnKMSdSjT/jDzu+rLQ8g2Y18xQnA2ztNxdIaP7UdfoTvOoxCUl4Z4EcG283vc/
NaQwufWJVDlNDbzwByEfgfU4STMFu1j80Ov2ETkKSL7EnmWqZJKERmZSUOUdwUG3dPoeic5vF6FG
gLHvaQwSTsOCk3eDWk0uHEgBHw2nILSA+rg+7hLxbG+05Q+jz50wLzg5Pn3oWIhdVhIrV7vCywO6
9BxOS/pEGvBKL0mQDSg1Ac7Q4/OpM/8a4ZZ7mPTOX/CKUNJ5JU4C7ip5ASeC5dZ8Yb6E5Qo4viDx
McTG6QFxqBw194mWUdxmA05HKBloS1bYRq6Nmmc8iwmvKDBMtyWnc4OjMbjeqxks/TuyO3Pkx3DU
9PjBDC8U4cAickUgTE4D99JCanRKmiZtjr/ECCV1TQgv7z7L/kB/8D6HQS9dn+bwoScgrSyA5B72
f/g8SiDdgiz6+mKbTRgIHgoiQ7meZe4B1D17xLCVsk4c2R9mH+ei6k+QNWxWaYJXBewgm5I1MYXb
10zHv1HFcNsmtMIPgK4l8as7xN6VC0ycXZdEdI+w0ZiU5zu/EsYeOal6wEyTAVscXXowHRsnZ3+0
j3kphqzM5RZmjk4fYieEYuS3/K8UogUu+Bn1M8etRmWMFd16hnf/wTWMjtdcA9SGlzqLrCRuaNFH
J8cbCt/7GL6zVqMRrqztO4aFGvv3/ob+NuPsxs7FD6FEN9A/arSV1K7z+ThVse0kWlADUVoc3COl
QotPlSqhxiyjef2KZA1iqXgi/1ZsaEWEOJT+xGyBI0dhuL03GDea0hKL8fihgTld+ijg2zc+spPi
ZWq3W3c8OKRYhDkrTeYVAaYMi88ex/H8Ih2WO10QFFwRMYd6LG2yoh+C80/DOQnSWolyil7Nl3dr
rd7ewVac7ceJRex+RWwFnZ1SGMoviLJmtUq92C0wPOWrjUV+2dbf2Nbz+eTsGS2HZgxrUOJ8lZe3
w6XHvr/+rRVP99ITf0c+ZEFaIu9JLMRor4d8WBCGH06pYqZgEIQkbHZ9fk++U6zSNKXpmJohry2z
F8cwHy3ciwKv/30QhZ1Gbaq5WsjNE257tzTseLsqDL761FJnlMc2L8GMjdkf4vxjT/9M8Y1lqvqK
tcjjOPJ2l7DL5LMzjkilP84St4zAGudwqJYthz338/HSxEERGE78bfqn3L5RryPzEER6XO0fuBgE
kN7IEVTK+66CwrIz9urceS6x4fabrma/hb0NXMfvgiboIm8MoXRmXJDWBxDgjCI3GBuGt9GVTKJ7
eeFCk7oh/HigZz8Z+vnt1FVxS+f+icmmvlbc3U6MwiPmK74QIkvTRqtjoIC7/6O1cjUnI0ghSYyU
fmcAmXCwt7ZneVSPUzSaEdANHZeLFSLK9USrOnCG15FHLoLF5okYBpRoIijT72jh9rEHUNQ7N12K
J64an4J+4jxGIRJdUWpMUlTmXU1E7ix8xsMF/6DPZm7+FHXR7pXm4PCxJ/g1+t6j57nWnBQEjH3P
pIdcrXrrEqS6bB5TW+YyPxiJl6JTW0A6taHbEXLHIIqsFUSO/+V4xQ5zWlstVEzVh6j6ZC5SRCkr
TLx28OCnxXossVij9WJZ7yM1Mp4Y+OSSCSLBB3ADjW0V+t02Pmw/p8Rl7gzYxeV9+FBwXhj8vgqr
jJsKw4lj7Nb4F/5+SzS0yjlT5XQPD3KZNzQMCcQOjulhLxajU2RiayXtDwpeNo3aoy4/21gGMVvi
YMTlDNX9qcF/jaXGMSpa0M+D8G6UB71vVSF5U3wUq34tNx9+kx8k7OzW1wAuAoLqXrmHP4rC6Rf/
PLiamoNvqvCdp3UrQoQhUjp8KaI0XhjY0X6B1XZrARSWCJ4ARDI6NvAIlc7E1ejYTTuJXInX2DLX
xEAfWFdazJf074nYz3OGnYyUUREWzQ7kXf1kI8l95tVUGHH7rwH+vpxRU/rxDZhKTwQw5BEmvso4
GwAIdprYRrSmbiQ3u5gduubLO5meXXJiwj1HQd+fHHb3SblRtdjnz2N5bngWwVDwrWU8Bimzo3fl
o/4Cb3QHrboQtOtRJIAZjmHmtymios4i4QH4/W1LJem+BheE/KDaQUN0dtRAjlqpD35YKgPhMhry
N6XED8kcHcC+bpH6340DxTh6TJKuKNquFzToSQyIb+7QZN0yabGm+IbDbgcTr9ZctqL9avTbsSKU
3Z4KltOD9JqCz/vd1rjObia0OhmxMbD/U+dX2RFVaK0Jq7EImJDyiglblWduTyEr+3u+tYl3AeOw
qaf/7ciCzZvPY+Irv3Tn5MKNL1AOKhY5BKyia1fgFO8nfjVgR6kTo/lQHgGlzMmDLlemVVGuw2hb
M3E+HIE/bZXZtTpaQry7r9yEK6lQkeWc0Xjrsi4Lrf2RaelEgafRQ+8LI7m2dl8NgC7S0Xko5A/k
3N33bdF6VoAJ9QjhOB+PxJkEqAfvliEsJ1b1URkDl4+K9Hyqeho1iSOVufpCKuVVYialsh3t07o6
72SgLqCPAAWDfJCo/RWFoLZ9yuh1uaZX5zUpE8x0wwit5aMMFBMo5lAswIPUs05ylGxlSLo6swjK
x7CnFxXa3g0jhme8BVLlLbml21dMt9K5sznzJ0gEFfSnKyl28oMRSzps9lAyB2sOQRgKU3mjwcSp
OPjoSjrTKhmftp8+nJFtThKZUHTfoApZ5x7pTL5HiIYS8z4CFbrQopZ+XMphSmERvDNklEt6CA8J
WDdyEotfPh+23WXp+VoT0Lo7j4v3HC3WwB6eOn4oXqitY5yPHzszkNAuZ6N3nutDRA74ayPBji4x
pmMWqOg4/1O2iti2cKfbnO6QJC2FInDb8/lS1S0BkUK7dQwmyzrkOTU5gntKzJzY0YFn1Ojjt/kQ
TaThb0BBHxKp7F0NUzgEz2ZJ98DUXFB2XD+qayviO0sx/tu44IzxZs5lxs1rdDaVQJJcDLgu4G4B
R4xEKxL2YcsJ8DPN/JZVG9kZy9IbMdWeR4ZwP8LG2M7mUFnzmUMJDlhZcraEiudxrax5UayfBFq7
VgWQpoTdYFV641p+aB3r77iSr2BPYxQgiTq7tpf3ZA6VHzicN5wHdHdZGgmujH8CiwqJZ4T+1DQ3
zNGrKRddh3xE1zxUuzNWopRvZEDeYzZ8/JtSO0SY3HiKTkXsksDsH6RGGm9xdGpBN+/dO0rjmjF0
rZK/fABkUsSgpnyoRHbrqfBch1028t8wvztGgNjq85AXqIljrCO3OsEWDUOzh4rJl7dtuLvSumPb
X3ezjE46xLShpwqxTJYB5m2gK62r5uQW+an5ESFbknWfEhysLBjk75ufi6VUbiVyOyRHkHXucnsi
QWPfKNxGu4n2T0qbk6Z2vEf6/BLu2ZQO4uyPPjgYS4MOZZeEu0W6s+9NaRiF1GpB9bIWQAzSm9/n
7EAa/9yS7CEylZsZLBkCRxYxvvWoM8CiH4Tp6nUIskeQZ7KGEbqI4B7iMlrE3JwdGpWzDk1W9yN0
B40NozTl09KEOHbRZ3kvOq/MXCodIWeNQUYulI1o34hKW1mJT1O01I3VREXl9M5Yt7GpSTVyELZh
UuDPzCEsdsrdEVRZH9ZK/sma5n9/zq84h3mTidesKlGApIgGcMs/DK63IC5TEJ1cpKe+G7ZX2Oib
1xMnjq8V8fmXEbkx0EHY7aS584/7KUNv/q0Ott41b5tRB6p+8FQpu0s/gOFei27mK977vlX+PnW6
YA6EZOSbQN8C59WRSdTTXKHy4uIpebpHban4bITzh7T+4CMOTqMYGtNJE6hB6U/w0DOZAaJLcU1K
O+tRlew3aDIm3n5OnHf+a/xqNlUG2VXLCtdh+FP1NuKlD2o+m+6URUuUZh23v1jBVemhbLgsc7ka
544pWYpLfTHlJ8/l8ckmHJc1HH/8EWuT+q/8rIPQm59Zy+lDINP+Obmng24bzitNQS8GmsX3tE8z
r5VHMHDnVwggmp7EhYjzQyzU8DUrdXIL6YZ1rXWQyKpWKgVEpZTlI/SVBtkrc9IujiODCSyhU+E8
2YNuIddZWadZHD2Ik01SXk6D4OIG9YebfrQpppdfcJnoNvZ6sZBtMtzvAJ/5+jjEutSwcXmU/E6s
tL8LODQ/Uh00iqXpn8uUto3rew0SLuydysAyIIZpVwIN/kP17Tgkft5vIrhKAOypzqB7JH0o1uFh
ZzPGt1PjsStpJPZ+YJFkNTRIhMipBjuLBI2RSyS67U/FfbnDVBkDL36gFEkhScXSg8LlnZlIJBdi
JA8yNzewUWNvKru9xOJgdDcxR1+y+NAlNjENYXF14tkJSqppl42jNpwo+fR8YCC74ODV0Z/aTYmB
N76IdPzkQs0zGYv0kN1pjNybNmnt8G9IOd8BR7BHjY+pumTpV/N0AtOa3l/zqo+t32Fy/WLXQ7sh
CamYFkjtQP1E6uk2GzdTnczzqelIlhm20eun3WU3pqh8f335tWEehOUelglF7ltFTKufVPPTrS4Y
eZ6Jb87nvWJDPOdNUenae5wvq/PmzUB7Y72tyblB36VbTEP2eQ/EdQbcpfduyiRWqfltgeyOyz3w
X0bwYtcwHfGsSGN9hM44RUmb5ZCmb87tAOQbsDal0ghjKprz5bR3BTbc31A3NFzjps9WEb+qysSk
vhpeMURDZlPhY33jzG0eqiFCjWEXq5WaHrnUkQz9TqArLLRa4EsY+bVasmTtqlqJuRuqeiZ9OGxC
6BYkmLZPsJbxwp7fRhkQYZDjDNLToZ+uQ5NG9EnO3e0EYr5ttFVfTszcjoN4SIj4kVUTh3W1a0Td
I0AzQAVt9w2dt8nP1fRaSrbqq9kHSvR1fNCzcsbjyzgb7VgQeDEfLqS+93+XRl+Ds+Dm0utEUAmT
DCT9OjBxbK9tUElGdPoSCNGsxGZW7Rlhw+rTTNKPVOZUB5vUkb1RTUgrg3pVjzGWivpEr8vVENLI
DqMiu1U/yPt8qSNcLlEW9vSKVKtckXU7yAWgIukl32FHHeSdgMabY8vjcqH6dmnlruCDcRPM36Zh
thxAe3hQs3CFVFVfww7uVsXvUplXUxjWJ+EdnhdbZ+VJdQPFpXojipF3JMe8FiSgPMISYlB6cisV
BFGYs6LkgGU3nFT7C5tRHt3ZnSq3rr0Me4eknd1vBd2A2mDkdxHq8XBRekCscKBKInqt+wodQ3Un
aNDv4Yij58XQZRaEKzcmLUJP4Eg5ySz/wbaIVozkfLY9/PAlUr0BbLKdpsPNptZMsW/pvowX5ZhA
l+w74SHxmQoNA8/+1UnU6BCh/mIBzO9nnmREb3nmU0mapENzZbH6f6L5pMf6KOlUgIzzqjKHelC/
YoVz/HIcZipO1VR15j7FMmxZET/zvDFA85QzJAbEbJWXb6ib2hatSgWfifUkL3hliqHtilZ6jOiv
6HgeSvHkS+C3h3esQVhELIuzLCaFjScpR5QRcxXGOlRapQNzlDO1NG5Y67DI99TwJi3mDh28jdDm
aHd1zJE59eVjCJSZjghq5lg8V4cyYf65k9C4nqJW2lKaE5QKviSapHrItrdPqSD7KbFkvXOL8Lu6
v45t16DQXB/nqRoRCLKMY15orQ66al/56LxtkU6hrJ4ZLqPmfAOGqd6gQvCrJvog3msIAkOKmlT/
s0ugpFK5iRWqi5/ewyeKcrV34sXcOoNic4A8Ynq8qBOE8AhwZkdogw+ibuO5sHPL3pRtsqtNU2iU
b1klsksIkxmuHcpic4U55Ins6t65aJXmq9qamPKzl1LVxcUoPTlb3VxCt2ISgQ9NIN+qTNOTQEsh
7zCYHWtop+V2BQP6+lBLTr1p/vVABmfr8bhfi6rQxq4nUNFc4yyNUOl+Bgr/o8ySZume5cJiJaZo
o5vaiR0JhjEbKuMkueR1x6nbnnaSFmJvi5iZV+nBI2rHm+K1AgWVvovHf5eLR4e7z4dvQX8K02UC
110k7g5+hybT0agVjpO2vqcy6+Of4wpXNvEF14da8TztYZhKPQvPi27Vn1teY+F2wd/q8LmJbamt
xbKtFqoWdH3x53xKqV2u1imTz8hwxdC4biTN1qY+enPSGyXeGah2JXGvfRZaCfBax8IQ/iAVJ4R9
TlU5sZlLWgzlCpxzvFPw7SgePualTu+Xqiydo2DatAUARbLCvjFdh4jjAiQPYukb5w6LnDOupxMs
CYnX7+PrHzv7QTqKRkQjjcQ8sV9M6bQgP75sxejq/j/gXrVmiMQBj2hEdc8Ify4wqBMiwg8PLMUa
92OL2SG+zsfI5xB+IGskOAF40pcYBkC/dPXbIR404jMJOfors7l1UX7F0bWC6ctclLXPBCm20FwW
Hf0J74Ou3u+HRSxd1F7ixrSwOf5anm1if9NpbRxK7GkyUQ3izq/uITPJR7KrYcdUa9T4fwLkhCpe
5KPTwGHuwxi3253jTNS1sBMs8I0S8iHt0mGq11Cy4hHUKveN9NOmCwkQH6GKWMCv152UWk+1g8cu
0vmUoZaul9j3Iat6UIuFRPHC6II3wH0TGzPqdGfkQxDSOmmbHaJy5oGKmg+fg/kE9iqI7LMW/AmL
283ukumtogMBAQ4am1TJvGoc6+OJHrHD9Gan1wc8qftEfv1gk99aQyJBSQVpGDQ3dEafKRpa4Drr
3jBaegJewWgK0pQiom2YXajcBrO53/gWf02fuOT4Gzr8T6uTpkp1ct9CcW91lDn7epYdA93yNVsM
H0qJNwKSIAO/J/ELqyfgqCRjUM+yZAHZL7YG7Ti1jzZxn3O3YgCxHz4KzEyO1nUh7VggrrHT/7q/
3af/AC33nOZj8a/k9zqRw37SVYuQTdpiFcA4TTQCEBUxamtK0UpDcjz2VLHIsmZHCCUUXFErTMdW
sdUmX428P19Vn+xDeGfpGm4ZgGD//EddXxuKcexoBEKSXPoNVDgupGa5g1D/N86O1K4Q+98o3b9O
6Kl8DFjBQhCSPwLLqHPAfsSlMSjQ5N8y4rUZllDksFT4/WwdPuHF5fhRISzTuh5m0cq+2jRqWYqZ
fne6NFeZ1NTYynXNsZe9269dsR2idsdci/bkUX4pXfR/8+rlmNdogDJpyF/faW6EkAcZI/i3cSPj
asLADhtRSSyXk4tRQ3I4XyUlUUQkJL8HGLfnuVq2njTUmnBC1UYO/lME96gcnyg6fcxzjCeXa6Q0
9XSCOftR8YHC99b3cls4dRZJeCzy6AlODwSgbHyFZHjYigEm5rU1OfWoVfxfyWDkk+goitz/6vTf
kfTsUkXvxLz2mK6jgT86vI0/bw0N42dgJ1JFzE2HqMjxAvwtcSa8c7hUITcrLQ+ZVc2sKnYR9qvL
SbmgucEG0iz75q45g3+2++qNOmcIpBBC65bxYnwmzOjTvthCJLb4Idsjfa7QSj4QDrmBTwoTxglz
g5SN0FfjRHbioUV+VmlOHdBwCPiTDkt/xl0I/59dBCgT/syEsWQI6FNickcOeqMruaGrxy3u4u7c
JBeL2ugEeXOzzCsTFu6Vkut/kt9yt0A0aNynbHk3bfIVIpZkT7MISs8rycZDRhZ3bCmNKgkv0rec
2k9gFuwlmpURlO0ANDAl1OolUNM8BnfX1dRrt6Pp4CZc5V2iHa6t672bUja4eizIsG1FT9C5PjfA
iC8tNJyVEvT486Y1WYQiJyasYB67TCAlMJdXz9IuCumzbM9giJclspggChDrJeYvvYvtU0hGL3Io
qAiGQjFhqPJHqJnD0oxOIXI7rV9oLZ201yJaohG3jsjSoebfwet+2oK5YyKYhgswUQPw6TBGt2gU
3ls7p5vqKm6NLfxJQGDqYRdNGMdeyND+pNOxH4lasxLDlgtZgppREYCYRBthciJD8sdTKSgPSc9N
3SXQmQa7dHyR1rqlef0nx1o/jbKlllTTNwSNdRJT2msh06aM+Xo9cLs2mR+rPH6QYC3uZDMRZJxe
VdedxcrBrPjFiYtSRh5SItbKBShvyjFX0fBbEKdQRkFPmnpHKayCCAX1Jz8ccuwHfTCyXrTUv00+
CZhQmvvpsR1ZKaOF82VnN49zQdL+doraEHhKB3cuf0rDQCT2optso2bv3MmbIsDNY0d8AQgE4oSQ
K8lkk6aNxlKKjie64D5pZGAKf1KoGX4R9+e+2MN+buD4Sz/USNhk0S6VBAJCYEHd2KH1KZ2625rZ
+ZloGdKeRGj8hUUpFO6GgjcZnFF996i9y5GcMQMgWX19TszfBkRVkZ+rZypz0xcSkDnA313Syg6m
IruW0ofEEIswzpFHTI8mqFuaUhocv3DqwPmXAXlB2Exf7iCT/w9gdKfvhlKZMbDi63fezu1hmDxV
nh/8vrsuIYfHofdIWdO7fYe9PyKpP/LABSxZDS/LAvh310C9giWvjqj3f+ifhrqt0oL0o2+E2VLt
xXmn9kO4r4Duhd5rD1MkJZrgMVxIWusd7Tn0YETAx+NhPKAG/FeUph7vDgNSvKZV5hdGuuXDliaW
vvOgv7j3YspY2gw9L/ujCHf9RxfX7LbmRH8gusGz1ghjl4X0EXTkGzqECNeHRceEBSyPvMPsN1AY
MAracl93FUqb881Z1BLi6kBp7A9SvBL5yvv2TDuO0hygF/92zMM1M2H9xxOoDGMJ8QzzSja2kyWJ
RMQGp14pPyuAYF4zB0bdxy+E4IrKlWYzxFE2dn5LybBr3bx8pNcoMt2/AE5GsyqYfvsl24JNQxms
1Wqn98WMvoWkce5Y10YeBqDmDBuXwbmii2SJhzgH3IXGp9mKSg7NWkp8l3Nvj+DIQoiG7oiyZ7Rg
7eoo4aCgAhlBWQmUIM4+jEAWH7R2V6OgJY3+OrZCd3kOCHVZwxtt7EsnZoV+iUQHGGy5djIkM8QU
vdqRr/Z4Xk/TK5xOjMgD2urGTKQ0lr3y1xaJ8oqdvm803vICu32seo/I2VGiohYonpcIYkY9SGos
UtPYvWqqP0jpTjnkOYS5Lq95Ik6SszDSDjxz6wAihjd5MeV608u+L7mEJ8EdrDBJKveMNcqJTz6m
cbGL+wxd27vasjHGKTb3JppsWMGvvdemwXBLGFGSyFgNIEfdTMmI4/FgjIRk7ZoxLF2VNyaGEORA
zhw9V1SyaeGzSNss33vYFVdPYx6mfqQuC/qmFR6s4QJfEM+M7HZBuJkuoKL7bb/5gGuIKeAPpS/z
SDUQGZmbWoGHe1hEE5j0CC3FfdjvS9xk8JgBH4+uYuLdMH4Z1qwBGbIdlxTtHQ/LNMQJEKemn2+j
Ht+ZFwwIf8nX2eysMJ6VqczqT5CjCJOM0PV0n2n/gpBMQZz6yOxLrDGgwcN9ImskkUkx6A4oGReW
D8Qb5cHK/a0UiSuQcP5WF5SA68Dsw5YcDaw5wb+sBwsc5g9Fn/64/f0F1Q3PSjkD3+TGUNCfPyhh
tXZomr/2raZQfYq9M4jgoGax04tuEG4eJQwo9XtSJuV/QUCeokeQfr4k0nBBVC2DZjy29nIks+Q2
ebn7UOrTXeYYQVqBI4+1ma+Cah95yIb51LhG+YUn+DKCh8VHgD0m/CTruonzJXvghNAxPIEFndUj
SrTrb9yZ2NrmHC4ALXhKk1K9LyM1pDKBzfwnuLw3m+ai6/Bc9gcJinckrpDIzpAsVQV3lBG+1fTb
5d11ZOct18TAfhE9SKdj/dSRt75NdtCyfjYbabwPqZtABxBYM9CAjUVjpZEAMvkwHT3m8BHVN5GK
/bV2uDObD6JZTf8y+VoPWhFKkUSaEuvrnAHuZFYyGkgIE3fK5w6Nh/uVMKyjPyUTZw9X+9B8P7tx
hPRJBLv3ApiIdbpTezEcRYiKusSdjgVxhrBLn7CH1UJMJ2IJetVqOtDCFQtfE2yuuwFqMPNF29F9
2aTqMeJNSeBJcaG662kpnRQpQNJOoU3jkDzQzZQzsGcBzjJdq4ONwRdbExj8QmmTe2rpk0pCYK8g
1joOhYSjE4dS2O6fTHhPhQktNgKdjFtzCZcP58eWmw8VVlffY6qGgwrjCdCDwjef1Fk1XAiResL3
gr0bp6/nlP14rYIkEK0Dk7yjOBJmlSQmaTiIsqSiR4MKSO+fBiyVydTmJh0IH0wT/R/JT/PmW9sJ
pdRa3LTvtfMUaDwEHw5s2/5BccpN/s88+YnklUlf6+4Zj7j3mLvSiTmYsYZyellgvm/NE5Weqc/T
17vtIdj73StxIVOecLLKw+AJy6GDlip7n9lWpoWpxJ4YDLkbPrl+ukpjP2iCIcYlPlJH1nvWtEPF
2aT2xb71YdSsjKkBbfNUDcIRB4JlwCR52hiEr11SXEIiSviQOMzpxIfIKGDWUz/V0NshMBisknbR
WQLJ+FB1ZYC8N1O8M4/WBcU+QQi2eYb68g0DGWqwcE29Hzubn9TNLtXNqb7nsbeLhTav9fRctzF4
+EZvUjwO7u83IKhAut32TIZWl2Xylfk2NeSELC7Osyr0bDvxrQkRvHrIImF/AY8xEQjjPHomDi2+
eoAYpJCImbR0Hdv4WW0vb7v2Q1PXTHpS9ny5srNLRgmkYnDt8KqNCXWPVhDfT2RZfEPyFxOoaWhO
cga8zmqGGQXdBHfjg7Y2ZTJUU8yGeHTpCdYeyoFgOuIummo3D0CaH12iKTzrbjk+fS5RvRhtyZ4M
LSiSz0+5leO8Jslod0q12LKbloz0FXNcFYYZms9tZfy+mkNofb6hKIhs991wCW1DdPc6fwa5akHL
EozCSBev1mVZmBfSK0Sx3tzALxsPaRI7Nsw8kssRDNOy4RF+K1vPhMf7zeFT3iZs3UQZpaKB7dQh
m5WEc9VCr7GbUGLNlepNk6t0+8/g7POcaybuPPGp/CL8++Vo59glGiyxcYyaJXuPlePtSVmiOR4V
uEB6YN3SGwOXYWE2dRjBl4v+jIStfeKVo+vJXrAFDDKO2L07V3F6NakVQ+pW2k1XX4mz9fvQmmSz
cyeqZQGRYqxrUvmkZQjz9ZVsv/bAUhQGyqxA9gto6QO/2IKct9GN4gkcEe1HSkWZENZKP1kFqBNN
b4TDjz0xUr0RwtPu/kHF1TQW2ACj0jhLzEsrIsGTkkg+0ESlQ/oHEIlPhnn4nNGyyMQvYkpQKpF4
y56YJUth/TcRfqIT3WcA18/8eM0w06l2tqiv0etyYZUQxAuC9iNrd3D/JYCi9Gr+RPueWpn7kAW6
OSLUwGSw3gklrf+2+Z+3R+q6G0XGgcCKAe8/csYki+Stjbu3JpRSaPtUn/M3gbR8WER6ojCM5Ley
gUG3ibNEtcw3GdnvKtI+I5AXzJWm7AEajbRKZnixG9JRgubRGH7HkGMZ8bWL9+F8YpOyGqE2TzO2
UrOSp4QB/zZsc/jLtvBuZIu1Bk3zbLT7kuWj53aLlbMknRN8aB2cPylS/DQG6FslgejPUPMjpqwH
UmDB80hyjV2fJXS0t205DPUOXifBL/mH5Po+N2QvNgkRYcWBVG4QfNpO9+z8ItxS8PFldrEv1cwr
Imfuli+7dkb//S8XfMKG9gzt0hJJJAChxoW4ifNmdT0+oAaG6Y8gWj+9UNotRr/cuVTkLYkQbtvV
qhWsgMYWBOHT2vn1NMM5J3eCJV3Rvq/ecq6YLANTBA5JKbFqCdhWKZXJk1ZvMna1WLEm5b7MIhiS
3C/C7A1lG6YMULgypJMcZZIzNS1Pw9Fess9rjtSs9X651YAOZKbnCCJWWMFjsSZKb5qK72vWVhp1
tO/w6MBZFQZzRxrgllS1AFcPcFcx+5X/8boIAdVO8XarQAULLqC48zLc2hRysJ2v9CNG8Agqmw5t
7Y3rhM4evjjCZHEvXX0KYedIEQ9Nh0I0928eymSjG8L31maFTIKiTqTaAGMi4k3nV2vUkj5R+YsS
zCKefH+orkYxjnNeoZrIRqN2bVeP6SUU3hrO8RWA/miczpWRv2ZxNcUgmwecCiDQjXx4vHJMszqG
39TY617s7pno80qYDw8iaV75Cp4cU5xwghP6WQsnjOA1pA3XIljYidpXlHsBxzFYZ6Y1JosLeYc2
COn83IWI85eKJUyuoLcr6rLlWGZFyOy2SW7oIkYOlwUtnxoKydMb+DQbpxiX1QjV4ImGPKcteLlR
bnzNys48WuEKhbGNEymT/NWWb6LlrLLe4ptx83GzN0IIDDxwisqIlJvQbv45A5rJfJ4Bg8CPEQax
F4Kfgrxw/Bq2B63EuxeSAwbNcEASKhLI5MoT0cyKM3iCSr6HLqw73F7vxJ1ZiOxQ07h4GNiZ4na6
aEZpKLMYclrTeRq8gSg9yODZRcFv219LQFbdKI4NtANgNtNYaYjyAy2fcZx1KGRa69aAJeSE8KIp
T2H58q3lPplpYWMWdkXJagwl0fj2a7kIPqPBrsCNL4F8RCZ/+oGhUzMoqZU5XslT11gHSEulMLZl
ZAbIZ8s5bw7UMtT7SgZViDIz7p5hinUr0AWx2ogYA2SZDlmuGi/qtCA+kbr4HAITRN7AX88hxlEs
RxZl1Ig3R8cJ99GLLbI6xXq4T/rhWUdXztcU9JOzUxwSb/dqa/cqxCBRVzJ8XtTFal2c4ZFA5+94
0ZmCd9SiAcpQ3aoidYMoX6DbbesXJqKP4QrGvEWgWBK/c0L5jE4ZUA/SolacoDt/7tkb5KWhkUVd
KKym+aQaaGc1mfwgV0O0zFFb2JoFLWGt9V11pHzjMimmVxa5FpeW7EZBeB9obgIep3eHr2lO0DWU
eHrHutQPRavwPPvbGkQjJn7ARq6CKtwqq1wVqiqrv0j6RLxn4Q0tZONzQ7dryM1ApSGCT/TJjqI1
D1OF9qVxBrtvyiT7DbcslIrCdqMSD54pZ6TkjB+NPo1Np7bR+/hSLQ229N9MoGT1tBULtExlBiWL
EBn11am0wxN4oZ5/CL7seHwGEGSGSFvDcCD2nweirAWPPWxAHFyRJDgpQ03mDxSRQgt1M0zkD89p
uTwNeWRtcfXDMBIzar8DbtZQ21LDFmUcZBJQdNexBXMoxW3yLPiSSi2eYWH4Cmh4H2e+iISpKd9U
0vt1g2rFLa1JjfPbYF10vEMAspdkWfHnY+XZONm/riE7l9phiNgRM3kR9MCTe5JtFTdxr/xpuEPm
hRsJl3fzKP3Ejf3ThFKmA5h0wcggUJGVKzuIqRWbDYR/G4+dAd2IkHOCTpzUBxHwQtK4I0moQRmN
VDg74RNYqNxNA+cg++lMD9ozLU4uX3l8osBTTx4GFGvdGaH7ufWJ1Y716OkAKMwnpv66PKWCgxrB
zpBkEBSKCLvKP52B2qrhsPaDM1FfAhbIEPD83+3Mz9VIJrPJHwc4b9umo9AAce5CNireB2ZgPL/f
lMlAMrKgrG/XXvJUunrlmJs5K5imZRSlP58qn1nEup4gpn5vykSIIy7BOoishC4a4szsFQCb/Qo3
sXO5342wxezA8AIDvEijCiSRmeAaxco3KVhaZfGXIrpApHrssYq8PMCGrleW6dfDFLGtNlm54tA4
LfIxyba0Io1uf/53tHT5FXVZrODTk55fy0IW6VUvv17Ik9lfkvvdC93Yh69zEnJhjZ2cpZj/THcq
o9FJ/7OyeqV57cqPA3PqahDX4TDs3s1ZnaBAKM5cwZ5vrINkzEtsOWqcisS2zBLBCHRbylvRgBgs
+exV7OGuqNIGiGtzWZNvihXRF+waEKR8YAubwqrYciZtP+1KjPoECXDn1rw5YZ4MjoVLBkT+gzZn
BEv/BB82P7nZOkuxYMfQaOWzADgSU6pVpDwyPIEcsrvR+i1mAosWLoI3/UHH4XorIqn3hvAJDPVb
aVU9cD8L9ztBrDIe8hGu3pwscrvMtp/ZGuJ3OCVXwuHWhDDCKKgEZ4a2tSh5hi4wgYU17iRxsoPB
qAwWVnwvvJkpguxmkGuQLAqgYaBWMqcxqgM25pMZRm53AID392PFTVwVHkiGyvf5KXniB6I=
`protect end_protected
