`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EsXeRsPajYX/YxoQaWaSSiCwfBR719VMFy+WbPGh2UU7Kp1+dfK2zv2NuQUxEGnYh2IsgOHOYx/7
4D14E6T+Iw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fwNmTuDBeFQhprdSkaRvfqp+4JN2uTi2veIKP9lTdMi6V3vFfJL2e26ZwNopnqXVxORqcIxB7j4G
1obXJPT2WSCL/0R7vCUMg/xfDg6ZfHRQ4HvE6Q1qt2f3x2eHE9gwy6LqEJ8d1O5yddIUz0vAxT3E
MCeNfnm0nCRZRRRR1XE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kL9kQOh4E6UtbQ/npzD9A5qvkaHmW4Q5TOqEPVqfbEiuDvKyIkPxWrP2j08vuQIG/7EyOqE/kj5s
ywoJMmW22K+cqgqvRYX4CWXFmZSBkvNI1XANVHol7+tm1Q6zcn4x8jo3f8GnUuBouEp969uv5TVb
C6W8kRmH5VAQXDtD7qgbVeYKswRn/GOr03sH8N9Ixf3ujy/rBmCmzDHZAfpgrSzHpSBDLuEk/POo
Xr9RNXhKMiY0o/UKBWTOczhocmLcg0NMSjuIOOn231vhyhTbXXcQqDAcqV0PuqZO7OgMM9AUBcta
f5wQBZ3NAv31WeWX668oqKgjV5YgAh+FAy4XhA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RtCEHK8hoBVXzxMIwgNIEMWUxUkR5Pqab6pK2iAMH+eKzf39R1Vn3oDa1Ljhrvx1X7iUngAsgX/3
LcmaDU9gqDte6ddNPkmbNLHvLhT9m5FvOkIIYEvIwBd4IBifYnydM1owSggUGKGtS8XQry6CERrW
2IwC+w9nzwdB76vItXdw1s4IymWgY5uwNq4//tpnCTkR/OMjCa2f6M9qEfWJYNlBJ+GXDAJmYmUS
wk9As7MfL7ue/D71kahi5ZCHlR1I+tDM5txkG5hGeVCdvwQTXth7HwqgDY5sYW26p5uvO2ZqvlfD
UgWjG10wynX2xKhSh6d+19vsIic1nRD2zh5zJw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R3wbUw2LtZKD3E3fbP2KygA45tQjKS5V6VfkBIYGo7BlcceQkKo0rH9dIS4uarIFJdlyweFapK4J
ePxAwMW5ynwhut3dqSMsEu3D/QC2USMsVE09S32y+GwiJIOKc4yR4T3A+F+DpWiAENZtryn6RnBV
jZ6etPI/ggwkkZm9cLyFuFK1/x6BNvCtmDYBz+NvlP64/yJ4zISqL2xL7EkNUjtPoWrn0H6hwsMN
LWmwS1HAvRjP69CtcKcn/ZrOsenLSCoE2qMOpIL4p9JrIN+PO8HJDrOUWtQU8AFS+CmCXdRF4XvA
aw3d/kbIocHUShnTob8znWjsVn39/MpEWEx/5Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NPgqApUBvoFW73rFSKf04YnhBIrA8CIHSiW0X2nssipI98eewlp5fI3AW8Y627oAGytBSN0EzSw6
6mWHpipQLQVJA6VeUIO+8/hOLRzTb+XgsgFpVaE2fLeCPOj0g3idUo0VTbgU5/uqesDE0Vbbrta7
T5odN3Lm9NJkl26/v5c=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ejAJ2cG07D83mzglv1+hg2mXZeeRNlGMZpMWRYKoOLgMgbw7dHfDf5ZV1yQve7ZbrKv4ydzeaMEx
8KfLuTCue4KY6+jlpd+KL0RPlmYfM6m/B1rwwR5ILj4xN3GdnDEXXsiMW/kLFu6ZLoD4Gg0fG+Vt
XWxnZfKM0dgbJWSRVoxq2KanJ2PlZ7qdlRIn3DOrtTjcJYuKzzGfxtNYdsTieTfk3SVn5bI2qSkC
3ck6p3do36oxO4wtfit92yihFVrV0gxzgLHMK4c2SX5FGVkm5jB2zgUjTl0KTI72iktv+yeDkEkh
cO+wtpTtK7QSUkTWzCgR8DX8WFsIX5CNO6bleg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
77TJFIvpXiL6a4RrmhfhZm/72rCPM62ubXi0Rd1zlwbibkA0O1BadaHpLDUUe/TgWk30/Hg5B0gt
0JXBDCRKGSYFfr3Q9+rqwqoGI9zK2klcmF2oOv2grRhzt6b1xAAAkzrhrpA5ds80bkd/ZYBzfWfJ
M7yHdBD8EbU8+dXNXz+9C/9HUg3LdNDr1FzJZ0Cz/zpeaVDWcSttT3gWJqJH0lnVQeEVtMLCiOtR
xVRI2UrllH4xzj+v3hXmh9Bu9S7LDXXFJk9ORTpj9mr1FNFhZfppAocEt6FZA78fKMiroYWzS9PP
ouCURfQ9SVVZGiMwM/lfGOK4ysySBuj5k1MtMCsKaRIDsjd/hiL7kJWMPZAtc5Lc7m/MGe/MriwJ
V97WZrmqJ5yrhonMZGFf+BJOu9xdzRGJs4pIISQA4FHuoNKNwiEolQQHlehX1OZKm6+2mK1A1B+y
s4lWL6s0LU+36BgS4YbYI1ueF8dJ8shjT4VbpLhO8Jg0twdUGgOQQ8YII9ywIrif13mpJrM27tK4
yf1uCbZ5EqiQR2VBNlLt0zC9zMUzlgXnAACvgnl3Nizg3/B41iQmSWbqoacE4v/u6Te7vo5cY4VE
cUkkeE6HEfuoFeCUShgrUzIL6O087f+Zr5VaigcRNdEJIPittBmSyHxLdZjxURkdlu8bDi0qMrr+
EFy35oFMzGPf5uucqrtEkfYGoGMZvsXPzUoxJTzx7w/j/WBhm17Hv0i0Dzd7wIJ79npLjseaqDTL
+pQIgQtmrNtZ0r6MQHEy71fHRlMtzMekL1aWDh8rJvu4XvpSnHo0upaygJrKu/9Ek8lhaXn0jXNb
5zFIOJ+0UFAfnYBrrmO7LDyz3kpptBdEE13Y33SVvRsD9DmX0mKjn3Km6Eguirq8FoAZuiH+Eejp
tS0H7WM9wCb0fP7fhkY9Kon3g1cXQsVBXvzaFujtXTK8ToKJewW7FC9gKFHdXMQyZbkjI3f1k7+P
BZlJsYs37AeDtzFeLSoovNqe+SXBNnBdFkt2YWIjjfltwvJ4GQYeoFp7j0VCWOQTCgM2e7hL04/f
3vEqVamCuTbRwNZHfr3IW46+9CqIxid06hebf0WsVK8tcIlGs7RkgsMO8qLbvjkozW7ojGcb3UeT
lGcwIF8C/gldNYCqo38DEq8AHKA4QPwLhKa5MOpOzfRmJirAOOcma0gOiF2f8h8FvDKSvJB6ESnD
VgoZkia+DX9EdOhd3Lupmp6r4m/cSZ+jp1TQYQC+s3r5zV3ogfYuj2oRxgmV8zQU3wpwWNFFIKt3
5xURxe7xkeW3kwdNGmU0tdIwx+62efEFNkztesSezv72ndmZjMamWBbWwA0ySPcWZKIqMtyTGopQ
2A0kMYGBBqkadC5kOKksLSSUmweovfXZ6Wk+H97wnIgB7w8HucEjz5kwyHnt62tFV9VaMC3qiMp5
FykY6mPf0VfYOOC5fgx4NwW7+H1adGWXvCybVg36GfrQVD1BKL8DSVymurrOaN9LrFrkGmPPN0zc
MU4RrZ6GOUHIyIfI1uUU9L/IvWFz1SqJFpkdkSRwJYVwKPIio5nwNydcB0uHGNvNpTfvCbQJR8SB
MeFQAHuW2JOivPXgU7wGJFiQikjl9oM5CbzJ6/vWmAUNjK32/00Angm2ELpVxHge9+Xcg1xj9njC
tTyXl8EaE17xuSX9OlTQpM8sF8Jgn+jxZONJRfpD3BcwderRCLbjSxcG5GAsRHHMZTtp1muMb9ND
oqZJCHapye2xbsNyjbRUS/V/ZOXOgTuXpEi06g+znwXy7XKnUV9yivu/5lbSNGKLMCN/F4xhtfNM
iTTeDWmSaYAIkgFEH90YUPc7tvPvB9MBl+jjz/44DcC+w9TZ0nitxgZk4k+0xOOm9aocjyN0qjte
0qRkjxawBX/E3q2mWJMtAq0qr6bXqZBVR5GoXJ75iW9KbgqCO0AX71uyJCJU30/qwlGpGliFRy9r
U4XUzdxKfKFDjppx0uDD3V3trmSQ85qCUKc2vkaBzS/UF+IGC6WiSDqm7iRjYA13x2iv4ljKGCQc
xkifAhI2qNJ2tGm8EfeLWco6SLM0yRFrZmqiYFK8cBluTrnWF3GBwbOMNm6gr9I32wWGdPnYD2dQ
DLkic/rmjyjFtD+x7aufFEjKxvqHGFfub0OhJMFDGIea16IeTjuSyog6VQctKV/G97d9H1am4EMY
MlU3xZytL1leHn09GuQPi5PZG99YMwsvtHM9xJJqOZk3e2sYxjrLd2aNXAGGc6wI1aNHv1VyBrJD
IMZ/xKv6jY5GMXzYFZ/9vf/tYPBRNAbgtN3eYA8Z8KFZTNXh0636YOs904434UQJM75B7p5msQua
2SqJKQOg7Ifh9Jj+5y4X2qDyMiCbbZ0C5plCkHcVx1siZgd1Ksfxrl/llJYjlj9CCokptA5b3ncH
Ed7Y9NI21tAph8oEJXkLn26QXIHAzrZycpP8AIzXEp+QF8BRAwPoxK0eFfQOoIRugisl43l+jk8F
tdwTYrkbGM8MpnVmTWjXuy8kj+Pf8drsqHruJBoNtOegUD7OABDwAfbNvh+7Q7xcSAZaTOUr7JkW
DnfF9RkF52LmFmnhGQmuzE/LVKNudetmWL/1c6GhooVDE1SuUPpuZh44heiR8CbUIyMh4THLphwn
1OA9gHfKiR6iI54HPGGfcKliVK8y9SwuAyJ+OPq3ypGUSOp+CK7heQ1fe2vchudQse+clG5ZitwJ
qC4YD6s84LC2g1imwAl587xfTdGNSML5odO1uuyVUe410DVijwT8PTIgqquAT8lzzvqi+SIXtOSc
rttCtz/QOWSh9Xf8aD3E9KsORWSXxdlmJRFmJy5mXfVr/7oxVIVuz3SVtWSFnqQlfidOvo9NhzFL
eWFgrVb1rYVmtxVpU5EP/y5Ctu9O/Vm5KoDbUXEso+O2pNvZy6Kv+ccheNCaCF6NpdSNh0b/mLvs
2RFoqDcpRsFw4F1eVZFPP1GKrD4B93GkMWMD8LJ0QCu9t94ePdWg9ymx7Bb5+jbQUaySlXy4Adk2
+Is03irzdkIlE9oA6ToxvPSTf9HH077GDCJS5tSxfkxQWHhHpyajelx6O7BhUCP4TlaTRbPCB0i+
7yz7pW6SyKozhtpsJJLC5Zeqovb9hWdQUTGxFPaxNnu8sa3QOAUf784EH6DMEHUStjrtofNgQgRS
aJ6UtGV72d2nNZT/rUa7yAuaHpH7NwMfa/yCIGnKzPgZu+Fu5n/UkABqD2312ZUkyFO6hCfeEx3c
y5LlXadJ7YVZzpUngL8LIeiuSnyyYwOIbJNEGmpBUbhL9sI6KGBim/BlVzNxMYRwUri45Y7pnoui
m7AvpobEtLTnpaa4MHwXeAB7xIJFRAvjXW+i0Tcq7Pu8shdmf7eUDHamdSxrt4G9QLX6nb2fPHCh
Sbncka2U00dt6DPlVa49DnXiUgnQsD7pWDPb7JZTMbYh/8juNP2SGIW7VCKOX5CBE2edhqq/yplV
TdzmLBTWTOJFcoULq9c/fvOkNYYsICRd8B1LdG0KybzU9W4R08kkH8omNx1TDqQfAX4YebAelPft
9x1IQxalRVcgScK34b2wieSWjkek3pIrIMN0qFPNa6CuXJhdfzTx4iMQd7GtxEXmQ61i9D/QSie+
ebLvGYQKOJB/r0ELexdg3XGmMkfm5H8lQ4VEbknkaQt8m28LoCId/Wq8orfXLfJ7Y6gygmCn6RsH
QiJGcI/sAK3qsnoiiuK3abObp9QxBQP0guFEltN+ultrqZnkqUPDF7RJF2IHI0mWGbt+xmuBHTmO
2RXkUem6QTshP8JY4gShpcRtP27TylWEIU22twVZPTlS6uY+KG/E7Vmc0ToIbvkKBqlFPWAws/q9
ibCPfhTugKpbvUBWzjzjc38zd3FZRlwc5fN/BMNv5MuyqAJBU4ROlM0/wGnKgFVEchphppVJTb5I
H4t7i72Sbv9JDubPYncptWV84YqVuJmLDcWI374he/KGu+8wnn0b+G9rz04I3Mfd7WhLtzFwCwFb
IxzQFN9Mhk34/3E16hZSvWQQdBZWp5GMxX+giBPin2VUmcbKoWokLhmISfsRSwwsGEpq27RyrOHM
jDd1856SDvG76ykrvGPAESaaK49vWcuTM6t/HN00zCWko24pFoZqc3aR8f7dKIjLLT9bS9CXdofQ
p2uIOu9XV9OrVN8f6+eyTyQxHXrHJA05eftoM+mp7f+yGiOLRaniuPRg0VvuvPBAzHSXLKOZR/Xm
g2nJ3aP1vQHmmyNnIEocYNVzpGZ0lD394Le3mUjd8Zyjavmg2TdJwmCRdMX5dZN5t+zphGZHsYEf
L164WbsFpXudbomwE1NDYSCCrCPUtNDrFJ5RpYooBfuSH91ErCCsZ2RJb/8Ijy6teWNR2PD8+FA/
1Z3tyNRmGoc/SdC69w/h1iCAmkf7A7rGGTNPZF5dyPyU25lYzZIb6v+m65JO996MvJNhwiffc3yB
TQLSy3Ne1pXiRtsGcHNbB21v3a/+oi2q/tqx+PyShr9/sEIzSg3PrQsXcVcFQpWNHFojVAXKb4Pr
Zg7vG+raeGdU2QqG2FGFrOX2XkJMD38XpKOx5tMOmOYvwqb9KzY51DzUlH0Go/rH6lJpvACbsD+l
tjD1kyfPT72CLbvSKzhtvPzJR6S7AjOaT1N/MCOzvfI2/aOkpyPFRx9uVScxdleFCTpI/5WWbYBv
8iz/sBqm73nTywgeBRLLPpOWeeugvRtQ+abTtF5ssO27ILegxTQZUGjP6dmPkrLBwX2xMFqR/0dd
cGRKLcIuDT3lqp9gk5HZNrNfE19rCZYiMGYbs9isT3UznJ6bvWE0b9Kh8cds/94B10vgqDyBAEj3
IzHF6wRMg10f3Y9oOKmT9u6Gz41+/SiS1AF5vXMqaaXrN8mxHTgIKrSnFSuMhDkZNAujShYR1RjP
gGEGQcVGdVPfYjz9Fa6uG9iPpxJKOvMvzh1IRVS8bs7jebQMv/o90KmbuyhkKIDBti8IKWc0HZfS
fWiETV8aZB7PgyLDRVzFbMMmo3+Ako4ShRY0gedE/KPD4lBGmtaTrv+ZJL3rZE3EPLK5nBTnEPmE
Q9Jiwd2HKJp+KqySD+ZiSdWIhG1/2TyeCqOcXMss8fTIzRXDbFejjKr/fptuLGvI9LCWFOJiT9QX
hlnvpDqZw8qKTQ3bn8j9o7tFRRqZMulAB+f+6AiM2ApYU3hBS1Shvo5OPpJI5gWXBLM9W3WU9Xs7
wTqI0x/nTmlN38gG+TeIpkcLJoYTrIK3bUcd+Cnm5qKQjGm9+m1pofhsMSuI4haxWpjIVtXalH3F
F6jQBe2jDlyiDZqV5/y/ZK4V7/PagjANe5T63KeDG0GtJ5zvm4GiDN+fwuiaeTnb/mEOb76wWf1o
1ipnxUsu7ibbg4RL5sjkLDzVOYYp2hPj1/Rsjpgu/X2oVa9L+nvYH+IXv2r0WrtjSkDYiSrMGuSm
FD912DRZIqQ3j0pogVsPTQttF2zoDPvtgsHJPsiyiRf0onMTdoDXrt5MrVO9ndB675RZ08+37CLT
1skasM7b8eGDm0mFxz7slZEDobg+vDD9wYr/xJ4l3KNEF+ooQWuZrb5/gKSDA92YHvVukqAuXPwo
z1vFB9FXJxePIUFHp9XxmuM+7cCiUE0KNfRlrHWHxKI32YiBqYWD4e+KGx23Nr3X5QKLW8Pc31QU
FZtVC+WhKhwxHvFhp2dsk8WE5UslybnUEOqcnCAYM8MwKRZF0U7NREPorIXE+k1+MRsXO+1uPC1x
OOP9PDKNqYTnDTdS84MdLSaSKGwzyLOPD+wq6RQPubH42n0QA6C3WAPSwUvnlMTVLRF6ygeOokA7
9CRjzhBno3vAJ2xHOWHNSZo7+lwtE4Yjrx+Iwf9azA5qK9v7WuLCRJ4YUuPpg4+XuxzvZpVBWP/r
3U5Nlng5mkx9a6pgaMhryD+dHgKOV7Ifi/wjljFcX0nCeZW50n+or4ClaHs1h0GsRll3gwVRx3Oq
Sl4xAzatwh6LiDiiiYNtNI40WwYwrlizVj4r6bHfvK1NhFRF0flAelCRd7qITDQLVEluEsSTM6O9
+2BonNYElBkIT0s78KHgmBnDJXvLQ9LQqGmJinEKkWf8TNJkIXy0ReMzTiiJfKICy2DinWKyWNPp
iBCps704hKHHDZ44frun65fMJO+Fxora9Utf4KPcB3+Y1EP43mq8ybJL/8SVSjeM4nisRtNNXQe6
Ot4I+lFtzUHoF6uEEbruoAn36biVIwwH8YQm4QQpBwYB0nZSPfFpCBXTPoMavsisUWXfbEfi+TXp
aoEhVnBs5zAns+EIksgcGGhn1F7ZaLklGh7PXTU3IFAahokuRFWG0Omt8cmrwLXIG8u4apZRJiXq
2iFvZWrClx6BK/tl7BybjIL1uRiA3hIc9RToaiRTe+HZ0lHt26E4OpR3b4xNf07dltRjH+7d+jYj
mG+i3DT+vpe+inu6h2l+mQXtrF5if+0tHXrcF1A2MasC3Uy+JOuz3etMcQUHfZoPo44idO7/8ZmF
WbJab9bbGptPIyqhHExmPJ7HvcTUuEzvMtlz5CBM7kSMkl/J0oK/ACnRE5rp3FU007w9c3Tq0Pzg
vjLp3wLas8cqW0vgwIFeuDzuDfQ5ELMEbmcdQQBHaUVP20BzTyBSMJ9hcuFxw3XaImwo8KBEdIvv
jnqPDKhQYB2Tbfgtx0jOahRgLD9IABxB8YNfc07gqkWeDrEsFqKLUoBlberyfIJl1PVrek+t56Nh
7yVmGy84KvccLab15hMvyxvHWUM/HvTBADmigJ9LMMRHSsTCiFwWmwmChcFZADN8Lh9V4owX7R4b
NokomFVH66S8kv2kciy+v9audc1vtid3ZKJloIs/v8Yqnwn7AfASw2Tu5LNZ4Nsx2A9imcidfil3
EBySoKOR1ZE7/AJRKghCNeWVC4dbo6+hc8cXKGLykt4KpyPiCIzA93Y6YshJWjqw+NSGMq7zV3Y6
95ErV/iWWdBlIHr83r2NwSPUhoHAfAcq+2jBL46muC0K0OKYIwUqKibEkST/FEUlnt5JKw1JOGZK
ZCam8aNuk2urWCXyve+73c88p6PKGVYdBEaqKj3QKT4LTIOozXtD8rruP4mR5eOEHLaxpITeoeiI
8tyu1NCOW3IViRbBf3v82PBjnM64n6s5zmTJ+Ko0ac8JxQyxXyNE5bFrTbB54ma3qWxYYbmHy78v
vLeDiJVj4OQLRXYoXCAbSp5WOaohO7rI2p/Pbbadfu2jXTn0SioZ6Z2NSJxj4IwJwv688gKpc4FU
RmHmfq7zmExbNuFMRPBgDJXrTBRemqGDHfhq9mtas9/PoSdRiiWTprE7VKJwLx2/uXShKllJU9Xq
/3O1hMhr/9hpTpxs90GyLWTvOwxaQZYv5/D4bQcpOmsgcOw4E0eliNv761Tx4tsBlA4Z8Z+johd4
IDXBjhRbpvY0W2twpFIFdiqH8shaaDu81dqvHNVXN1lGNvMm2HVjyWdhN8AaMXu6AYuj6tm2m9Qw
i48gOQDrXOfAr4wVdLZV+PtX26432Txkb8xBaZPNuo1C+OaXBSoHYKa4Ev+OJm249fqSmjFFylRu
IGgBpR4J5XaKE/886/GG26d5M9GsWq5GGmv3qYNhOWewUfR92kGvnSd+bJFnSEQRwvOJqboOioT8
tc6cF0Osl7qf58mYu4GvZKSNSkMDWIGlnY3NwrfXm9WwaEukz+8BReVvU0Ji04WyQ62ZGlBdrycF
IoK/0lpymBJeAUtKiqDpofxnq+W5I5GYzikcaegsuWnuAkyHWGwAQTS7usghes5++DJGLHmTwR64
xeG2ul0XPS7FM1zBOmV0c1MAHgbbiCSdX0IPk9QYX80OeXs+HfAvmetfcYxnTresczf8kkETcAEX
SK7usAAOUgoh3E0CCC/lOgzLqKWakQu12WBUVkBsdpqBY6QLUH4Kv6JTw7THcEJgDwigII67Th4C
kiqKNwN+WwL7JhBlA627XcBIGiyDPDQ+ptYhMv1ggPJ+RFSVBjAYrcacbtmGp4GaPQX7p/RfOtIO
LMpTBtzYLYWKvvK4TyWhjFY7JQnu0qV2tTB42CUjZFQ6gPUiDhcEYu3VapZN5h4qs23bjf6TBbji
qDevLpA/+Sov4J5YtC7KmnRlMwB5/a3te0200Ftr1RfqVO0wIiBk6pHsnhRl9taXSwWneaaeLVT5
Y08poQNn1KYs8Ua/fl2cpV04zLx/CqVsh7kSQZeVLHJMo38UdRKxsi5586r0juDJET/wGgbs+c29
Hg5nyKjVUAlTBunepfH9tDgskMbm9dmc7/U5MJXF3/lKKVcFms2upeu+KjenUWP95cxZxH12tH1a
TiaRYah0x/qLArKv8+xl2l8voUpD2vjbjvKEqL7/ePxb25gartXYk191vOXhdqvpn7jPaLoxay8c
PbSeQGJJaqOtWJZ8ou1QfLGI7oSq+4BHYI07iXZpmU9qyn2U3miii79WbeLwW8E6TW8gPgEP1pyp
u+PPq0iujY9yU3+jrAuXqRMTtOMNeVsRDNdKCWcGHSmK6ltDcG88avn1nlLHja6rhNUeyyFitWHR
YnVMUJvZobxbdk08/RGMdlajTz2Ruy0tNk4sDrlsvrN/FOIbvBp6YWq2KVJhyGgWfeoO9e+xLQ6V
JXkaZRut6tFBepYkgIR+4waCkAe/TgQtmm4BqW6zrBMZi9eDEYHdDCuF947N8q1DND2COAURhobo
M6c8e+OXjH/18pYMBh9WG98Ls8vn+Vqz5DxMhMza4KNJ7OOzQkJKQ7mV88dojcH7+uh5lxpeIr+9
KO6RgGC1OyxqTi7p53WI+b6HBWpIyKgnR2TAwNrkwb997Wbvuh1JihuwtChw1L2SNrm0uyAC9riU
uoq9gcp4RLQk6rb6RleNPzYGYTei07Ea+lLdwIps0a4IrMVjcZNSL36XkmQdBU0Sf3krK9pcgw76
k7mssk/2pnXX4D2rTh9trxQcn9mBpK9qc7Pp/Nc1QNsrIbHqzwZN+av3Lg+OL/L81/iS59qb+YDd
Hh6a9TOzIfOWtSXHz8bkMmtwFmastWDSTNMOeZxzNh2HezCiLzQ4fr047SeSOGnfiAGFYKZyuNhV
zzue6FDctt2wmMzuuFne7jjgAuO+un/qM2vreMgLG8pbiZqMFmwNjMqkH7lLHLiREun/JcdqntL2
YzwVb9vZfDHCu6lo2nKKpUXHhXRKhLcH/yWk78JixIhJ9P67s3qVteoCUMawebFEXwXgf602gQN9
pa2p0IeHld0LXfMpoKxlOTK4ofijafHtknphoPjDlh7C2ShQfNrq4vfAfpPZen5tUC8gvvwTDZq6
KncTa43/MPctUBwSwIF4ZuA00Ev/wMpfVg6asMJ5UN1sx4WESBqU6WfaNCP0gvFVPjLsMF/ERsc0
5tqQFfKygqLLCmXcjGqFo4+Or3LotTqm0CS3Yg2rWnWCiAWzwMZDmzCglBq6LMD5JigVWHciOh+B
p2OfZR1GJb9AHegeaR+LQAyTGdRgt9WT5V70Qo7Pdi4qTs3cgN4PiMKhuN0qKo3qSRTESO0vvM0c
64MEYERet8kjYKgZEh3yAhrrHD8LBQCUocbz5LT8PkmxCfrV7wNWgUrNAIXajfX6ZbAAlvon2Rk2
R+IHHcRN6wH1vi+bstibfS/foSImazJCRBbiYcKeSRG1lgT/lLA03euuNZjSPLdHPNm4aEy176SA
exoxmq0nVPLxQjO75gnsoNznJzaDxA48wNtoodQXzmKrn8G//w3F/IF/XKaAV0XJhGOwiCOn6Osu
ggUCgps8D3oZvj0Jbu3oN/vcltIqM3uA/6BGdUw6IOU406BNWXi0ujsvzdzzCpUp+OCKe7OOD9Ve
bpYD4WnRhqNOesOSmOGasRBAxXuBblRYGEDt8MWDj4uU5/YfsH9GbHV0NJwdeISOp7RucHKmr/cf
KmuE8B6pV7jEMoFM1bMtX5+Yee7ZFP6MNBtTQSy8Umy0yn2mxlaQWFKY5TCI8srzao2NVA2KP8Yl
cUyul8EeRKXSWjR2CA+7+6JSEVAhn6IzHruBf7lYiMzatFuLZE6T4oyCwy1GccrGm8eZLESC8bxu
TGGwWuRSGjABNpU14LaW4uKeY5C1mAbNLq6B/8n5gOZBbD/4QUJTlMwCuTJB5o/C3mEJKAcW0fpv
CqnxT13zY9gCbdEhe7/yWPeHUnodM1eWWblOpfzfKumoy/dy4qQ+gqfxSyUNAUl3hpobY8kGY8+l
Fw7oiUq2YDFXuAKFT7E6YSB3/WuKqbuhd4zG0BaAdS7M6vFT818yLEZWmMRHV4ynTY4HWXWNOZAq
78xTkgL4Jc7hDM+Ivpo5OngczECQJk04lBot9Bl0N0Q503UtnNGQUim1crp/Vkt3hZrS+DeeLn69
wCk8sYEsgC8SOll8wU+W+d3GLtUZT8pV2F8Bk6jculKsjfj0DTFOGC4c6kq5qp9P1juvasJNQTzG
9m9eMgmfxm3TdS7AgZusslZsDBNjEXoYd9SDLcPXEwVKtIaeja+h7WJKt5HDgcXPCbPi+A0CCOHs
NmcA4GFt3XT/P+zx3ZyfbR+svLWYN6zlytqjrKwwRk3pIW5WAB+YSo3IwjbBdC9L4OtjKT0r7jmm
lwXNnaK8wpcV8JeT5Cs1Gex3uFukzK+eMKQ4acF2FovhibQ0W4y1SBxIAwkRb0pNzgaZsu0LxcS9
Y1zn9Q82ClEnJ9szTRSW8OF/WbbOu1GUk1nfrKrwtP3zJgPbEuOjHlwUiAbA6ucL5sqNTXi85ND9
ID9Mk6e7h4MRe6sN7CZveVG8I11gJFCRpeVerG4wxENUrn+QQOdCL2FBYv1L+FlM2fW+ev/3pCz6
KzdjKcjYR14H++byexWtvUNnIx9qBBlM20Wi1hJAu1hE1JqKWVHM2Q2aEGHLIao38Uovk9HLEHYF
bRr+aVxb2drt2ZeaRLzDZASQs+dLLV7WQdvHbCAeel+CdadUjScgEqHcTg2Mo+9Xxo18b+xO/fRq
V4V+OsQiZyw2BlhZJHuSEHeTQYvhwm+U4O6LBJrPwpRblZNfLCO92bDMEPB9qvDq8ly3t75eU8G7
79axxmKMCxdZXPuyK/a5mXrPZHV1AfNW+mnMmNE60w24Qs6JgDObrO9p30uZj6u/apf3o/PQTwty
FXZ55Mps67MGyMXWoJa55PxnU2RfdqAhHkLolCAUpvez2l5u7+my5QFMVgNhE+fJQmQojnsy+xPN
0feGq4DmJxQRXWhKXahkb6bBDzXfSnMOnasiujoOBjZGAOVjI4CXkQBgnDpPpwo6rn682pf/pCGA
hA+BzxFJ9GouSbzOpSWF0y3/vcm9e8WGgfmFyU2ZNyEgAzGE97BMtGbF0DKtVpj5fRjeVzpPf6Qb
tR356KV0L8YG/o85KEs1TNVsoM9BGcSKnwo/SfPnGRWZYFu7PSjtWWzpb9fygHBEA5kS51UhHIku
CJMchKbz6eFbdiVYbwmp702uZbjNoIZHD0KPHf6adRKoh5lf0J1Ns7uwgVelzS5sepZ3YL/+fsX/
wVLHmV3cOH5VGigRdQcFnJBfMRvB12ovtnpppomchManvVCO6lcAEpKeCV1IdnkcuZj9+be68cac
wrfnMopm+BJKVj/ATbhePr53FHbltInh48H+cbxmdUPZTyddEqFUbJA2t3KjHqm8BiWMvB63WpuF
VqSCvzSJ4ETauhGUf4j7jH3eb5op/WX/GE4zyi7huGPq8G6WIOIb6TrcHNIwqTCKT520cuXYtrhw
KdOLWrEpLnYLxUihfQel1NnPt7fve9ue9N4MQtAeX8wi6zmCvJu9HSBWjtJU77KS2MR4PzW1rnhs
Rzmwb3M8AzWJYYnVcXy4lTXhjBJuivcjBx531p0/mT7Qe6mAKvbrWlk16DIQzgADDlB4Kc8AlYi9
gdx8qekM2BsBgBywxZ/VpM97LYvNhXBQtviGTvkP4l2iFQqSu9tewIXZUoMC4TnYjDnyPj0e953t
bNqB9RMJQeznBqxRmf8cSpkpmn+D0XOIvxIhYCxS/pFhBobfq6sDhoFSlci4ijODOJHVuPFylam/
V7+iwHbDJ2n0D/umt5zJ/jtHO1Fq3x2PHFcntBJsApCCEPa+OpAC3VBatPMIzBQrujJhO19zyq+S
7MX/186YLSWCFlbGNzrlq45CqvfwMQB8f0+KThLOGtOCJyByasT9YlA8xu01E5cnLy3xM10pwVYP
nSn1nnsEKiHgyVJsiKdkAW9EUiYhnRnn4lPKUGLPLa52ysthCuuwxZ23RMuBjeEEuk21MAXOzR+i
/crb1kvKKWv12zwtSJtGuZTOe7VX8B85LfvR9tMPfPZ5ZXNFEm2Psbz/rBAc+bUv17iJniiay4Ho
bw7igKGEYkRxNy5OMaQAB6TqxfPDJrjmAp+7lJLPhbKcZVI0bZ528dMKIYPrIPtZe/Acq/xpaNd7
HTfkeF6/LvkcVM7wQKUVOAfGcbjgu8wKRvYUrDC8zIr5XbCvJ9skgUZTkofjHRjC0uV7VYu+xpz2
T1lzJLKNvxMgE+/elNn4gw/yq3OAPwG9VHdfgppZJxx3Yz79VU8EYD7Yls1t1vyeEiUtHEZ6oPZm
Py6wAdTVRjvDO986bNQjrD3lQchFkC3+CX/WR3kBW55lM0D697WXi13JFNkURgCuh6Lq+46dUnyg
5+QN2mOb2LA0D3wirBrNqaKOpaDL6YMEnv8qlUL053VBkciFOmIyBqI82e2HxZtqDlJ4tx8tl7jA
0ZqHW3LDWyDNfy8x4IcFUv3UoPddfRiPTOb1KxwAYuwaMwYVfLyOsHxb+b/wmzYX+ssO6T6XzBwq
yCszH7UrUwQ8QmCV6IBLyJniJO2R3T0CrBUaFufcbi4rQnr5RB+b3F7GoBbhwjxXOlBUTZuSojZX
F4n4luROnP7zta37GKmGNuOlL9ADPSUGsniTxBL0mXKxxNu1Fg2LobnwrGaIrBSzLTpIB6VOzFPU
iQVXab8afzwKwesDh3MUUu1UiAcMQMOtUdyn7HpPLb8u8pJhglxiOm0Qt9c+ZOkp1aKfVCuLznuC
ms46S/XbFUr+Cb0EmDPysUptJhEGf2IjtCjq/jcO+0C9Dg/Q02X6t402Sm8T2/1Osw/sA9U6zsKD
RRHqG/rhqDPWQwmbMxCuwiO4JJBHD2cqe2poUkA9MBV0JY7UZgvm2FY919uOSpRd0kzzzau+skX5
yvVk6QeIkGhDlkjssygzKYzzWwsw6cy7Q6TLMXGYAhXC81VVM0lJDaYDLE/BRaDDOfrXqeNWSDJi
FM6npgj1GFEelD2u/nn/axFZUnjZlfgToD1umURMdG47D2v9g015BE+BgAX68cgExCWyVqgt0zdc
anwelUdg/Q3/J23Suw4zd3rsfJCdypwsdFIvN9lxTNfk3yCLIgcZn1KawDmUVMtcdkXeRBH1m4Bj
rE9rgI2svCDABbmtcr5BLtt4xAG6x/KwggNVvTajYmCoOgeUO2tTMb4SZVZJZU3S6x47plykOzcA
QYqvrmx3tlj60iTBNq701S2hRku0ICjebbYzY1xFUlLfsKsvyVOYusbTT3PASPfZTgnStghUT0gv
EJplr88lmzSjKVha8Lsno+sbLQv3K/7QKQV4waDPNEQjJnZD9dl2o17we5S+Q590GSWWKKVuqD5s
yPfaJw6k3Hk0TLcs/RMBcDFl01jPyMu1NANvcYGojw7D41nlqTPBq7I25q5OgqgeuSWu727hsT7q
tf8rn2ooFsOY35iTPbZ4hujsmguxXqPNj+Gbhe0eM0k3EVnnb/f/Is8nRINAh/U25iGWgtqXZAM1
m2amtog8bjBwU9ScexOlznmr15m5wMKofQ/au/TmwoUVaWri6UtRRNELZzqCIMErsQOkO83QAsgm
oqjHNptffaMtL3/77m9PiMHOORVXkqY1kWOpc9+QJACJDwLIf3BCejSj/cjxsp4faQWJxronfKsg
lN1XjH7UoaMFROBWi6/wZdq3slVNn3xkjX38dXyqBJIYSPy0FfudbR9+KQ3ZJxP6Hs+n1SH3/GEA
gZwLBXT+d+wiOo/7mxCtrv84omt5wByz4pDg8ZGFUUoXQqAO89WCa4Kb8FSEEt0EpdpeUuC5RNI8
1L9daPKsYSXPWc9wxKnLz+l8RoZTnogk4rWceBpb+/EuZqdGF9/zY6Z3jBqJXBD/7MLx/Ly834ik
zSu6uBra3sQZfvq4+kh6irQh9jaqt6P+NM1kxBHHFc+hdY6FYRrCGKW85vW+NyUqx2vRnRB9Rn0m
UTo8iUkkJow7RLNyS+/qEwluBqtf4dVXqSPFw0lMqqjVM1VENtut3jYtpy0gTLDpd8MltBba0JID
LhNSFZp2mvZHYO0lrWlO8Er5BVjtD2dQ/ZcJVHzh6dZdloko0WRI2Nx35HwO3P3lxt00MOOSNPLy
nI/DAlpBcKF5lhJZ1HIAtBNLUxlJG4sMI5EwrFIRRkNp+xNkl+gyNDPwvlmM2X7OQQGvbumnZGmi
he6a9fThN1WL8sZ/NNrwi7vbVQd0YqXnmy7QLDiVmdmUnXL1iBCNQkSWPrSWPOwfcbfLnRdHhYiW
B8Kw78gwYytEoUXfmzVA1exF812fKkcFFV32q80wUxXZLtRHNQSvMkMgE0B2Pan3g1xDN2Gdyo5d
CoRYsS65NmK7mKNXFgKJ3JcYhtuhxsvsaDT7wmzJSl0p7xE/5oM8BkDSVBc9d0S5fHAW7n/3Esql
TNCjDm9x0D7HaOlXURtbeNnchYZmePy0p2Zh9jYuoI6mBnVn0RD+ltUNbzpl+TUbFgW9AiujRXuQ
yZXgo/ZwWX21m6YgMBha/ZpR6Bpho1gCfvrKvU0nXUPyTaGlZpOiJtYW49D7QdJoarDBCxJ6iM1g
jd6vOv+41/1NOMwuqr0UDay86TBlDmXp871BmXMlxf98idB/myZav43viufdy5G1tiumSiFQJUld
/3LuRDoNCM5mCEODmZXjUg8qZA20sVv/qiRiVU4xZKx8+nuf8BOkVHAFxf/zdzfRet2SgoBhCrfh
b+fgukhPiDFX+2HbMZJOouCWD7CGHwoMODLgg/USTgSI8gFXhF5S9dEpl5irKMGykxg8zNQ0KQdb
sC0ylvEG6n7h8HG6ta8JT7noaEpZeLWrj5aXe+17FXt1keXTs8EOmDNBAn0g2XyL3Nio+TQV1pkU
jmvIpg5a2I4eAfEbx4f7wEtrOz/JAeLXRhdC+cIzNVYDE0Z8hpPgFTu9l14lPSVZmjIrjnsq1o9h
j5E0HKwDLbvjUz+oZw+tQcLny3+laDhTE6Bvt7eBJo+9Uk/0B9BCYU1v8y5zv9Xv88hebk7JTAcj
HYhXlTvBb+NqMoJufW9nOGvrXXE5+cdOrOu3GXYf32OsNl6BkEo3ujRc8VEsUHBSaICIWAeqczmQ
jzhAfGN+UYuGPU4eg6JhrOYyFoG4w6LJCphnZLZMTxke3mmDy84y25yij0p9pLJT39oluszudFsg
N/0knjunfaBdf+yoSe17xH+2Za7FgkR0nUjJ3EqeB5tBMExXyt08FYMPkRa4OkkeU3E/gF+VBYm4
daj8WvYiH1BXssgbJs4tBCi3Yh6G3DIz6f/9U6MwyLPB68TEjp3mmnesJYLTZPJOIcfvJRSnukB3
NJcZXWYkmQae9pKlnKAVKByKWtRu5Mob16V35GFLot5Pmb2niNlGiNZfdv2HDTYxU1+D6US3tBkp
znTsQ9DNMxsA1ymDbBuWOajZTJOq18LEANktDr6et7uuj1GpQYYyZYTmBmv2V8/nRrl0/TvcunDW
i7S4GW/HJKLQG/ab5GleEwr6nBWJhS9bsJuXL7xQOIBwHuR3K4uPTAQG7TJZn7KxfGJ0gX7BHAZo
srhjAk+m1KoHtWBiHmo6kzVMhZil+T0F7U59+k/1GzsX5AI4D9wCOiFzfCwzyeVyBM9QT2wTSbjC
pYxHUArBg/fFcRKGleOh+eOqmSmaorZfWnT10/jG1yIIXyL2zOLijnJ2bGzbP3WTt3MFZgGDXheO
AwPf76C4NOMeca0LGZaFUJMiAYRkeMeU3b5SgcWCAget6xjO/MxaGR8oZJQPNckHApGN1N6KJole
dNDPvU8/YK+9pyWN1wE+fqLYn3HH8lAz8vQRP13F9Qst0qICix65Z5Op1Qjk6FOGKte2GTpRqZOg
9w/ZgoPA1crZpyXWYULJqVhHN1BZmZuE0U5mBqbZHE6CC+0zwrWPvB73fHk4DARcqLy+2JlUlgxr
eN70SfP7B/elseOP6F4q9RsN3QvdolP2Ak2TBVVPSGGVhxfBODAtDLUtXtI+9v0xs5BYspT1fspM
C1eeLPLsyrbf9QO1xYZJNTZ7OFXO+8ExVTx8MyM9gu3TwDXS03VVbzQ47bQDeK7QZQ1Lxu25Ebft
jAh02pFgRg+uju+JiV5vttJAW8IOTO3HqmctvI93PiFZ/xvqosvp3SSVRuC76vQyqlqufB8dAWKg
LqAd+Y3/MAwCKE1t08nHN4R8gs7dHuwv0h0cktUSWQsuqgsJw5Pl1VE8DHaPUPKmmdCVgg/wqChw
wGfgQxiHFAwPMHCkdW2USW3yX4fnEFyOBVkzo09Un4oQFkEYjHs3kN6Z708VwNBsIT1Rw9ZH3C/D
2NxfHxMy4GZToffDrR31JsrLVlGvWmK0e1v79Vz8zNvgbMBp/tK3lr6lm9PiCdfHyHJjwa7HXMWj
S+FQucZ4Z+KMkWUAEHpoNd1igs+g+WEsZoEQipk0m9zZsLcftZMr7FGdil3+5bFykfGmgRoIF1Di
tMzQyL++9cGJQ9C5F6z8Q3gMYSy1i6N4GOgh/JGzYiWaP5/ZVjx8zoOltHkIM1TByNkbEiLJrXdy
Yn/3yZHCcAIRQZq1MZh38Uvspm0Di+Po2QuL7F92HYxc85uz8mqwbN6knJ/8wJHPy+B90bb/RtPf
4/1qkLye0/5GTu1+cbRmo6IJTgak9mCMLRYB1VdWclpLq+SR8eYREIoDDFzUWsxsesk2VCBpkMSu
5Xs5paLJVykS+OcXU4ug8NlHX2Ax/bcq7lII/g00xhgcNINvsOiZWR6HEyEgMj6nWSkdUZq7GWCs
N+zCjJdTygOIOME2hqWp1ZD110hIa5rJqnRQTrrKzN4xQgWehyYg2I8SUj+GScT41+TpSa2PGnbX
0UVBGvvLf6ozqkF+IWmiy08k4uQ+zQUt8Bwm/44tVTEuBnvgF4uRIjLGW+QTvgsU4H4VcBd3m9b9
Uy/6jYdZ6jzaXepHmQoOyHyAUeK5gFtB7j0GSTVqf7HFaoh8VTruiC2W+05RG7T/7z1i/Vb3nI19
pz777rGFdJPqkHGVcma/InIy+Nkxr3iypDzVvZIbTLfpAiF2GegRboCZqYa3Q3dYS7kIvM0ZUvDG
zQ4Y4kR9Zu/OLl8ZmKe9Qp/R+M21Kcg7fuUo1cM1yPzbbl9/OshYxdA+mYp2eqY568k9eSZU/z1D
xqtfnS0YnRwYdiccrYidPg0klU7sn9HwbI0133iV7Q0bwo1PersQtbUHEA6yi7brCvaVx5aCozh8
M+BJzmCgz8XZmKjIQVcJHvCYEhY2tzThK6dg5LsZGtT1MAWUeb5fWwzRvj1rD8O4E1dCN2+3LPBm
4Fl1Td/gIV7+8lRbvl9rva3izXRasHxowEl/GY+k0J05hUVbcIwhVVrKpa6q+5YcvW1Wjk/uEmz/
tqitEzGJPSRPoUJwwU/OpNK2YRYC43bRz+A66g7DkUG96SH4fuMLX7PjEO2NCuWzD2QymnWQ4iKk
kBBMXfWKObDqT/CCr6g9hGBGLFOZmvSNir1kdtXHtClVU86p/HniILK5FgoU/Ep0WWyNZY5yjROJ
vr4WQQGyvW7Q1YoXSxbCYCT5++BzY5bbCur/crN7QrPxRexw2jWIwmIEqxGpkY3vUo25veP0DpcU
NFyv+79e4quj8gmBnBkUZwOXXcwfIOfYIOIkgAEosKMQw3pZBo8/ZVD6vGmHM21K8ZHit+fl2UHI
eoatCIcovVfkKsAPbu4VovH6mvb3w+LkB55kVJS+ugGb5sROhELtKPpTLtIiyD6TB99QQYUMlRd3
jjEiQGKzfKYk5gKswCbdB/fMmzD1bGrP8I9RZepwT59wMId6rI0kp5WPIdlzhF5NlT3aD3Huj1Nr
NjCA99QthQhMQZI5kNABkWGNHJ2nCkWNoBJeOPkgYpWZ0TAt69yRw5yG2gJ36Fe5kj7D/WGGt0E6
qIBjNcWwpE1lMzsrRKs3UhIXxw8I+mdjyQon2JDAwHFalPbEOd+IYjKFz/Y+fZOYo+r8At6kGAxm
XJ+HaK9v29elvS67QREayRKsWd08U4T64QLyR9Shc1HHIeXGik0MIVxv6Hezk4gdXWXUnNp8dsxW
+BL4IO6BFH663DFfAzR4ybz/a/KI2uovpACGOweSPDIORXEuuPxTvZ35QGMDFqAi2UW8vQ84mGxF
f9X7Ci93icJPEUOVXIF+sSiqQHPLdBp61xhAW8ZwAvBkKqIyKARtm3Qy3hOW6bYp0VzkAdLMgPmK
cK06qHZ6qCVmFrtNNsOHOiK6ZwmjerNHpngwKsbZkUbba+5SVe7dkumfmrDLyf7bw3EUHLQvN24f
J7xcpGJKFbCCHt8DtAYITQU03D2mFn8nEylXn3m6CqafzD/3Tf6l0Wa0ejMTvNpx3rK2Ps4Z1l18
V1dJ7LWUbsmx/y9YGgnDvKD/yPwkyJAKnT9H/R/OrW6NIsChZEL0VGf4DIlfATk0i/Af4PjeAGHc
8iML7CYtsGv8I7vsBR6KvhgQlKZ+lKzsatWaOApq3p47jw+z3ypVYff5l/jMakTYJbrNB8iPZxqd
oH481Jk2FlDGMCa1VNRWHJDcTNEZwXBbTGP8njLCk/97L8slLR3iD2rX9c7oxcYif3cTt2yUYriH
lyWNm+Zggkglu+oLX59jphVKPdjTG4aIs4VWjZpl7kZmWEyaL76zC9tBMEFZYqWvc0pSesWUxKqR
ir8vCcbB+mrX5HqrRg07wQ7LjgNOqL4eR+AZ+YiZ73N+10+YW1PbOIXlYwiNhutfETbLahOfbkW4
yzEBXmykpbE6AUuFswDRdrUzNLJ/t1uHPqzm4gNMpCBFjWs0NdSkdk4ypYOLQZNF2gXUOk2EdsSW
lRA57E2he+qWev9FU6Fq4G2vc6di+rrcDo6i4+HSmLd6Ek0qj4YKMhm8kbSggrTKDucx8iBU3qnb
ivl1jV4D0QvfLnsegRbc8VBaB5uAkl3NHZpZZ0Y0wP5eG44MbfNvloVNc9Ats9ajBk1cYGOEfgsp
fIN7Uj3Acf51wt5zQLg7oBVHwIcRRTDexcqEq2CBvqTkLuxJ5LrDlZQVdyMHnACbhiwzh6GhkfT6
xt6518AITw/hoBMTzoSbXN4o/t4hPEGY1T0gaVQRzbf3sZMQ5k8jyCzhGgKLARSTbDadSnuFGehd
iEC9YbA61Ft1+/JqvZr+cOrhKu96LLMpIOe58YQTUS9iMPTuIpxvuLj2xDbKmd21nGAeKYMcvapJ
Flpxmshm782UyGm5TPVGf5hddSQiFRQniLCUkzVIYPCB8Ghq0jVXcsmPpwVDHBNuhYAfvMfRWxSD
g7YkL4OkITr/PHoMD+lbMca5mXTvYe6wdxrrxi4NLcm/DZpJ6O7ZbCRbu4bU6x79hNmJjy++w9gB
AQQf9pGeV9nallOyqOyTTM+PZFyZCHhNyWiK4OtLD0U/MaAWbQScvdEDyejxrkQtkGejjYVafmCq
0PoKTB6KdrVvXF6HEqsbD0ztFQce9fyv/y6sXLzhmL2T30u5FMHnBueKQKByV2wRGllx7eBDDSWt
S1iiosit43im/MrqgAGhvdYHMU7HhmJYSdWQYl4aVzKMD33wWZm1grgfQCx1tk6Ti5FfXFx/DP6D
l7O3ygdtJdk2Y0XQVuySDHRIndIOuQkfOyqu/eqfXhrK6Avb0ia7nKqK0qQIHgME3Pa8nap9QtVu
+NVkJQV75sdKQ1HU9sgduYpZMk8UAVw4NsVtLuxmcCJZjnVKJFhhWDyvE/3RskcYqrFcwFcTFeIr
aFTNLi+ieJLEOOADQjxe0rvRRwX4CfM7tXrgD8P7PcsNmhE4m8u3g6jVN/gj/SIs7m66e322Fi25
Ue5p2jaKCZyo3pGSQAAybDq3cvYtEJms5oRiJs0ljdzFZ1wh768kjOya638/Bfd8l+mPc5KDOQJz
N9r5Fe/FKswCEeBHnDIBxCcHKG6dLyVw5YYl0RzqpBdYmkmOrKfWQb3RGxzk+8eh442zTdLm/+1C
/35kHApw5OcI8gFs88qOexIiT4GAoppw9voCbgJpcawDqYmrCHkWpedelaQlmlA2ehjZNRt0w8vY
SLiJ3427hzDuvo2b6pwNCCc4Ma6NQHuTxzObnnyTfyDf0ntURRLq5j+cioMuCSDP9aVBTsMZH+rN
LE1d33bzoqhwqVNjIql8jj7JfFrXXoPGamEzUVERvEBuBzaiYdgIAswd/PyAJdvwtWstA8H/0UNP
yN/I4JUCEp6v+KOegLWU77w574qITuVNN7AVgTZbYd79GXPuLe+VaGBNqAmUZA3FZUpw0DdgTRtI
ujl67xFQkk5mHrwtdJdZv+mkH5Z54bp+CsUQz1fu/sBka4vlKkOVLSfHCE0KFFBzRZGkr1AnDS6k
Q8gEmgcmsgLKkjWe7a2v0OgzUJDVISh9QWgFJabpBTFHMMrv830pNbIefHbhM8SGKJl9dmOENijk
E/Wz4pL32sSP0rClSDfDJ9mUJboKGMO0q9Swl3VBDXJcbD94G+EOV+kBk1OmOigS5f2pJEJI0vh5
2+VyOKbQx/J4tWEKnqvoVMs5X4PvLNS7i1kvk1THbI9MmBdsbfXzXmqUliwbBf0zRTDQDcJY+iRq
QuXrpcKoLk7zxR9xX7XZz0mIV2ELQwXSbTQt2YVP7OQMLyv/kQZSVEcoWfQaN+33ju+PsS8UAPUi
5sB48DjNjGQLlOiPHCLSaLQGr2m6bdkkUX6J2sTmnDl819VHopt/tzYmaY1McIx6QU3mSSh1Qkr4
LmKQo/Sy1heYXJXw1Z5ZZifetIWmZq7evZ8Rg2rNtXfSk54LVYYUj4937OzmadEDb3EniDOSgomK
9fmwMcIpovtopjvHiDutLadko950M8NNDqskn0mIgKOgdch7yqrlUO3+zDOFAO+pNtxs8uclwsPu
pLK2OGiaI+H7C0NJLBg5NREBQyXr8vK1dUpAKWU/jICJajUPGU+hzrCdpNcROHHEPepRljfWYSN8
UHb+1p1KHwuD8A7fo7XJ2FeLvIsfSJSlFq9ScmkQB1vocW/52X6V0SDiaVay7YyQA8uOaGEhRsDO
VzLKASZjqzIKP9B7Qhz6+uINNP1CyCI8+nHE4pXQPZFJI/wXRep5BNNJw34U2CQpII2N8YZ787OL
DQJikj3tdBQHqEyGhmG7sjToBh9e0Vs3pgixSzVx8PGjBmwe7yfLctP07QxlhQt+s/BMsJMkYDtH
e3kli4zO2GqUH8nyvRdNl03GSrePyNS2MMtjl8BoB4SShVkd5ifEkaIaG8Q2aYVEtlf+XfNDuiBI
6vblG7wRpmRU0QqJD2s7w8paH6rVGGyyKpYIycqNwynoK9AQPcWd40j3KZe5qfq50sPrXquwoqMO
ySYnHUbeKnRiZoaeGtVtw12o9ZnqzJAnD++cQ8C/hcKiC5puzHq/OpDciuLB1pwYoKeZke3oN00I
XL3Yya68r7f2p8pQQdXPAGr98xn4Ea4WGsaZXN3lzXBqR+lqduL+L+aRFYKPqmoM5j9/uEHOGB+4
gLXG7dUuP8JF3LCBbcSem5bnvmwUNNxQiWtn/ny5irN0qa0WPyiO3sb4jYUPGUJ1mcVRtwYkJ7nH
6c2iF3t/62DnwnjSSpmhcJjOf+MBUaTztszLd3KnXVucip4IHGTMs248YMd09rQ5QBry+UKFWzZq
atr8NuwWq/WeLjd7IHoqxACmyLnqQDcyArE8Rko+qv4ycrZ5V5BYpZHqw/Z+3OKQw6WIRFr7pC8L
IshHyGeEuEPvU2C0pcG6leCZEok2CTszF1AZ13j2BgnQgmpFU8KsgkWbgd+p3J6/E3gkTMOodBbi
/0bFkm2LOSp1WzfKaCMxQaY2HEc3RgADBYA73FvnIcYS7a5Ib49LmrQ9b0EYtjrzIhhuFHz4ETaA
4Q7UnQUiva4744SDq3fXfZ3WIFT/nDmS+eHhLPLSVD7c2J1vepQHOv7EY1L/Uac2eI8NwXd5e4vw
lsf0zQibGeOuKkVE3McOw1BHVGHldYXiYC6Il7Hj0tmUDOSbIy457sIVLqO0WC75eTzjXBZQbDRF
LGOjfRPwcdDlQYj1ocL+2pwpCWMq7cG1Op95AAs7UsOS2UObeg9K5rH9EMW1i+lP0K7Yeop0azQB
7lSVWcZT82BHX15rWFESJ6qN+vy/HXuTmjCLr+dTu2geMB6ZIEiRfz+zRx447/IlS/3uuDYnJhSY
2z7w5QcB6W1SSC277E4FrS0wD6I9ZLBpTbnPMLvkeab1DRDaTfp+d8helBXl9dSAJF+zRiHKeBZf
+aQNyenKOHv2TLlYYgfP665LusGcPrPe+ya6J6yZuQAv4wIQ7dWqACVqCnWIPHj5Mo8/9z/4KLA0
Tnw3U5MQVAakLn0dHxSYwYWVqjVaSKEDVYxgu5dmXTv9LOdC4UIxwy8vy8kQeVbe5sfvpyNa8su7
KGHanY02A/lrImaH5yxnaT67vYTqiVnNUgEQV4axeWwGjvxVQki3RbBgBPVRmJ6hsp3T0/FF/CW8
CguTLgIn48jWNvB5eI40Rdj6RuFmNdqcRLwEF7C3aqydb7L8BTUSnHjXtLMLoPJUOe2xQh3S2ueD
lzX84WWJQ7vgrASf4kfkeE/+n4k49UC3ccFtPWhM6/7PzLCiusKcLMVrvKsx+sFyzxWksp5DP8wl
4yHS5vTRpcre8isfyGLtkUg2kWJgD10i688MNlJl6OovDG3f6C6MqJf5S9Xi3YohqARgyQk7mBe+
TFoBmdA1iY/sC7sPArsyPXcgq0FIG3NtDBu7QxyR3qaR9i3SEnKeBIKxX/83f0PMZyYSmUQ6wVB4
g9bkZAf7kOfrOotsNBaPOnpANADnGh9DQ+S36HudWk8pFEN+ayrUsh8scueulTTexbDrN1UAohWN
ITzIiHfQOItW6o+PNpWP0f0W16/XIJyzdwctIfQ6P4eV75Hqf/x9YqWQI93qzXUbIdK5MDGDj6Hp
eg2CUiugk4eCfbBoPf9g/653dWWKeW15986BHIsUDSjVUG8EkEY86WqBTzxrJ50aVaZ/9FgPHUIq
X4JQYcGF4bvKHixYB00hLMmsxbacH5RXOgqAovdoys6xQSYtlNA99+TgPQxRsRztGeU2qawnSIGO
vmK/vlRqrrGzWJSYhGso2+y6quBAVJjFGjih0oTsQ8vHKs1wvURwdAIVzUHIOf14WapLxqWhkYN0
p0nb1U51WCtttTEBFmpiu4ti7jAR0O6f7MoZAE0IWtjGxI2/1pm1jxsuFjHHdZ5tiqBOyDx2+zPA
E43SA6mIE6Kf+BcWphj0+Ck/Nr0qlD+06fj2zbALtn2hvgvaa+1n4//5ZC+4tWUPSktyV/r1SYYL
NO6bFTLaUDOHN0xH44qOKVKk1L8mrPQEcHACKoosY/KPvVgrysFwnPY9CAPs/Hu3XYS44MOkp72e
YfrD5TrJAJZqFHQJb6R223hy+c+dBD/q2/ksvai8HmzRyEfiCbOvVXchrAadIg2B/YF6AW1P4GiW
d7ax9IO0CxTqXp9C0pVDG0ihrsy5eYPS3NzkfAW0aRVa/JVoDyFz3XR971qpz6JfKCTYBRKFOpET
iCFbdcEUSewzuBiJBLRRsUNoRXKEyqU/dWJT2a6uFIRdj2LiYLZr+ZclC2/LrhP3pMyoMbbPaZWz
zUNVhXCej7ZxrqrA5SjjSiOKGotjj7fakouXtwQ9/+XC+ssAeeRL0CUiOLN+UFsZVzayAwgYJaIk
H8J4Fpfg3qRl/WdaMbsVRajtR7N2tmIpoFzMf113ZkqfeNuiuxWEd/epAvl+KvujjzToe3C4LZEL
3L2WaCdKGejmYMSp+cWN+XlyPtvNFIZ2TVOsRgiyl0wpXmnPTZNq/7kZSEv5KxiNGSdSmgD37/FQ
mazXO/qD+SZl9JxneMTPnMPTFhdlk8koDHBFn7JdtFn65DRL6QlPZlLznmztg+UYoUv2iv44A0Wq
pmVL6e951g3nNdiIe8o0Rv0G+vUeJZgVNXcV1hLc2vH+jTcP0WTnxji1U/ri7Pfpo/sWUUZlYCWt
deHQlTcgL/hpIG7e3gG1JjAe5Cu0UGxK4iKtHEThLnZV0YcO3mUgjkwU7Dhp0A9DQ9s7mQIf8PHx
IHG9y8mzYNazXjdPoViovx2rVTXaGt7Qs+ZHUBbHzocx8UnFG8gT5rp3GMc3DQ22Np4a4F0eovDW
j4e7ci6x1kLEJwGfv3QFqTy9IFmBz9USn1K5j97CNCztzRl52VerkxBXz6OVagCjILoUYHh353sB
Dg4EZ2nGPcveb4uNf7ePOlQOLQvyGTtyGoeuCz16Wcvqd+pXt0Oe085hPDQdakyChTHdIYdwV52L
rbe7rbCcF/ToQhZcUPu+6w8pESE89yBvVX+HnXku7RfqjNfq3nqATE41DlpEwIB1gs8QLc1FLU52
5ot1H40LXw6uBaISfX8wOKATXoYKCMAtLK9hHRabDh8PJ9Pcmrl7oLa/7cZiOw8iftgjVXMvp/fB
9KH+Si2TJ18aPq37DzcPdaC4mmYms8iqfPxSfsLl0B3LRC6t8ppZ533d+G9m3txb4mE8xcbI1TdO
dBjGFvEkJTvLYwMSiAc22uoij0tIwHDXPG/BnuJPlmIqw0ylkOcV7FabS2dC9j+26pMR6VvSIqPU
HR/giaACn6bAVc9soaNubuTR2slPvAZ8W6bTgNzJJYdam8NuhFx4RLuciHCbjydtXCC6MglY+nSw
OsrrvjSnczDL6lBdU3Vy6W7ye446AlH1YPF9AD/EZLSOuc+QjH3TJfNXRaivvXNxcFkFND0zI3Mb
KcPfr8fD49POTZhZexGmtB7FCuGZV2FhMruh4ndXsYNEhYeWZ4Ik5vpYRQ+xCGXsyb3bv9i7aKF0
THFwWxwl/mZukF6L2tYSUaW4Bq6PHeGBRxxdaKEriAq/KakeYq02a7Saj2DsXxrNiyyGKUggzn80
xmKngkTBnTMf4Vo7iM4V2bRgJMF9fUS+LfSNtcsFVXA6yzNoPXFsbNH1TERFtYVdY+0YjwtxvJzK
XKl1uNeFlhJY+pjK3JL15cyQk/CZHPdDD8DTNqE3VxLWiuFzPnKe2xMTBYfLHnMTsXsl68I8epBb
FyY2CcPQR4WPfvKlEMz1FssB6OG+ri1OQ57CQ/DhXf9WOnytJQmu81hrnfUE3BtKX8Y5yZilatPK
S3e5+SrdIysw4IFNpUzaFCgkeOgx007ttVITy7b41e8VsLZniIE/03+QH9SBBBT7H12k4temtAzL
s+cEloOmImMMcECTLAFhtDphuWmeWhS0234O/qGzI4l47cfYma/ZDLoHYV6t8BcXuZsq4afgAUKq
3FB/yJNDmHsgDhuPZgHCa8mD0dx4tmabgzFeuY3lJ+TILihplRtXNFHwETDE9tkBnU0Ujsnhqa1J
IEMAK/kGyssBeU27SCbwj2ON70xU/Dz60JrWIfClOg7U7oz1Jb6ae54f3ZN0s58LZb5tkOPcNQni
+7YL89Cm/dBoNBqU+1hUMKDrPc/vdg+YCkYPASbpw3u4/h+mcVIwJIwaT7WA7Wr7qADlGBPuuzB3
aPPc9vSknGm61gC1HKu8iNNQo7wyB7TNjqXJ//fikbWcoE2pmMv6MVkABu49Fp7P/9HfRLP+8XzU
QtAgckurUu5Hd5eq3pjVlnDk6hh+Txe1xUwbqclI+JodKnk1fahbdBd/UjAK7Ch4CutOpxufnXxt
rc/lX7CxaNr8sEwrOXzcJPiJ3lRR+8Ui1uAGZpVZyNOxVLbNOnbA2qF/ICv32L+YxevZT6oa9z2I
CE0dLKmCdJNanvOCfYe4atqnGNffv7UI+pK5Sl1LLeAJn8rUDWA4KZRb42/rXzmnBV1t7o8OoXO1
nbQmWSA3dqOrrIbnt1vjCbprv7EUSLlVh+0C8OpxzWNFGv2PeYL5GWuk7PFnchMSXnQVtAhTJxkL
evdS7Gb9QGvFrLEo2i3mFWZJmdBhnWoLNZIbJlgpE3NmW8vImwdvs83QyqJcgUJMUvLjVw6q1kA2
RGDWtYxo93yn77D884P4/iIPMX0r8XtkBW3l0dm1k2TO7FbnU+jSTPWdEPVUQMYZjBkZxkdYIeEw
HDFIKjiCWBmoG0ubXB+g9KftAF2nSIsMhJml0t26SDEfve4gXwEwpI1x1tieU+TEiK2+K9QOKQTk
F9dpExLiaURjryw9XKbdzU0lD8oO1n8uLq6yDhG6YZWbg8s41lurj8EzovJzyswzc5pQFoFTHIed
NTRq4uai22xrPT0da4KQM/OxFVNCVYUe5ITMCZCUzsT8WzkNPqECUX0bN4TfF76/jU/KzuGJNCho
3KMbzbvZQwZwDoQLm7qVSuE/q1ZrR5kqheOhV0oXsGKhtl0g7yY0anFl0IqiyJRo9Qja7GqFgzRe
0E4kNhax9Ks2vDnUTCyTJfAfvRGPIGWKIvWD3OiRJNss10xr4pSksO+kyXns4svEprco2+qRdQ5t
u/wMxxnKHmInu6kSrBWh/OWsY8BjSTWa2E0PvnQ+zGWPFLr4OaCCAcP/VUhfOSrLMlJm+TfnioUz
PWM+xPdLbU/8jN/fnRMSo7nuAEWWtaNMUv8d6JgdZY5HH4gn/IabphiIN1578SmA3y9SV7sDUcXu
G7DoCKLazEMUnPq0gdVbcVxkPKkCtqYoBYWFdJSM8oh0MMUF+kKkXTp1WtIrMCJOEpEGGAySw2TG
8CtObE//Kv1UmY2e0Nt44rlPA1jd2jeYF0HFbcMcVBdMf0FZo3A1IrmrxnKgL5Z24f7HAfY9nBYF
fYF8QW4PcTAe2/tfUqq9wReSq5p03Op9bLGmtvwQOqdjXyPgqncfbzoZH84s26F7mxg7kHvKLstJ
8Sts1/5UodTMyNv4n6mUJOv0/90VblsOxA0sGcrRGXMwBKdOkJB8QVYqkXNhLzJRdNxdoA3ZqGt5
FESGU5DiotSkFi3VQrKn2fiTIbGehA0d1u0VDOETSdcd2BEA3RXx6NH3OcxwPZMTsHkyderjGDhU
IJrldQCbzstc/iqu1i4ksNeT6Y+AvTGZj13dql8Jf6MBmUcxbI5umt97vTcckR7XvDKUBW1cIXIk
QdGWUtRBU14E0MFoTNfDBT6sRHPR7fxiHbcUhWH4lfNEF2Ywq+xvUCuYW+TaKqZ0vudIFBilOSKJ
Xo4fpjXtDaNZO283ZNpRYfYdrdS1kpgg7ufe5XN5ota3EDmrHG1qZJlPff0IrSO3mC55ZTDyZr9t
s5vGLJLylTjfhbDasV7t4yTbqfyljzYE3eW99G1fIc1Cv78VqkJPhEEUufUZRondcJSTXpRPSrHU
ZI/QZJdzBw/aHy6va15BoRGzU9KSqbIpppPakhrYaGejZpeOSvfu5VlED67dfO719LhN1dCwF5GS
a6i6/iYPRzvttGtqzIe0RTW00v4PJiSi4i/hMR+fur8h07NLs7wgSmT96PB1dN5zrImb5XsRwMAA
Uje5o/nWirrfmiDO7kE7gdJ6fhi2ZDQJEJqYgG26DvEQgmDuspaIHmPzR+Bn8zOHIsQXXzBrvcEz
JeX4FUYTbs9Jb8++fu7s//cVgIm0iQWDhBeQbDvf7K3Dz043/qRVBjwkCJNdmB4fdjTHxgMbSyIA
NIBMMsnCsJL5eZ+MRpSbFVI18nm9f3q3KCmdxYvh8xutNwnit2YOOW02VNT3stQJ6ZaeSuCywf4t
OGU0NFH2paK5LZ3B1uR5ISCHCSQIV/8kxWrt9S8rqe1DGJ9MTI3V1kRXtynyzEutOMpHE4uaaW/Y
cz0SCyocoWOOt3gjjv/SDh+vyiaRUSVQ3MREKcGABz6SsdFjvacwpT8uBwQeuDzJbmc2DB6zlh+q
f2mloblqVi4eM6T30zTepnKMqodvZwnfI9ZZ4FYsEu50lRbu7VI8E+0wBEYYQQGmVYmmU8Ms06XP
duJZHD5SrM/atb9ZlwMOWyF734Fez1kfPou6Fs29lqYBuD0662z2AYEAfzJks5MH3eTb6M0Fojwt
uRvVXWaXeePmIvKxRT9p/gPQw9xnK/8u4V+d+dHTy9rGrAtK2N0h6Dl9HQMSG052KATqo6+lTace
zZNXxGjOLA0GXMA+Z02SrOy41E09PYOssqDl5YTZreiWP2qlhGuHAxR+sb8DvzdWDAF28USsds+3
shpDZVE5IIGNHDQoNNRRhdZbNWxZmNTuJRO5lY8cX8By+6vQmZ4gV43D+GbYsKTlsRG13kDEUBgy
lye1HOJlUyiqVJnaL6iolJ6VDTIy+Ki9PKwK7Dl5MCM7VbJtXIIVaXXQtHYFh12PxOLkA0uZM3qn
I97U4l6ZUc0Wnsulroz+EoFTIyfI59E18uEJf7wgnnNeJoUtcl9oAnggf3Om47bV+otwXfglQZf5
Q11SFSzdgtRd74R6YthDjjGf0Ld6gwKMOPu4gG5Y1SMRsS5CtoUDG9WJwDPryLB+7CKDsYIfNhjD
SSLk5OZB6phLQnLS/RHNTPFoiYdVk8OkyHiqimhMLpvCZkcK459g907hkxYGHG/SwiqNtlk4bx4A
aghB3pHCgOuWACVfLOXzfBs8dk/dG+RKpQpJevpKiA+i419MxVbjOFyGE19BPFR1w0EkEQiECCMX
EoQaP9Epvt/KnWQyp0xyY/nelaghpfoDdcTiDQMRAwhQvDK3Pu/jX2nL7IAgA6L5eFyZM0J8mtDp
rk5UoLbKbOLc+TXoaupb/qoKMirws6VNqfS3ocWD7lzL/2uhPy/YO9I4g5OAXtbnFSILwzAH1G4g
QF7C/6GodpGy4ZRLhAFjfn96qJD+oToo+GqyhTpFPHbyU0gMIovZYKX/lLQGFjPFoyH8czNBXPeD
78igKliMH0YI8BFswKL7VwIVgwt874wPDwAv4GMPaC4vw7RtgO1RxrdzHS7514pwR43EFOcJUnBs
bJCTClYcaYe33dEPlR0m6EKPi9RSpjUgwl9T9Tx/wN4Dl/fklV2bFGlXJbvlpzcN6A7JuqKjZrqJ
6Kfsu4mOV3S+aFdzSZxC3xrIC5u7sCefRfut8blCtGDnuhVxaBeW6+JyZy4cE3NLGdAEte3VmVF+
dGlcVwPDONWC9TpdqBbX9Y9w3uv1D7eTMKfLmqc+ljSzMFmCmU/JomvmPA2B8QxR9c/0WP5RI9ea
H+Fye4Ki+L1KZy4TfkiMo/eeIUmV2BwXMiPDgMeUNvyBmpPuFaIQZ6gfqQSJnJlutc4ScxZGim7y
KvhU1WNntVDM4+maNtB72KNCCkDZERxKK14i3wtDiMUZq4wXuYYpgsHsCqQBW227TuA4Yu5KmivP
+kdnfmL6QGpojBz0LxF0B2YU2E96IA1npJL/8HHP1wcUA5M5r5FI/fdE7iKYGdNxNdwoQhRQqnvL
R9hgyXUOhqkXXjNlQmfmzpw0Lkeya2rpx5WFCMsF3iOt3Km+6bLXLKEXJYcx5m5ilw89O3JihHnC
tftir3lobxL2v5sSDKk00kveacFHnivGeeYcbVD6anQll/3MushKkG9jQBBquLO4UQOcT32ilSzv
b42Glx3ZEZIYqmp3PSfcvR5JvZJey8fSna2Njj7Cf9wKb+BVrRM/+wRSor7Zu7WIZCocB5VrzRXO
EsxQDhOc5rj2VMZ7S57x2Pz8fkimnmruYaEbAAkpvEnEmU30pO38SE+K62x7lxgfKsThljdqJStB
fwKxIxfaWpXV8LGWoNgdYRJKg5cygHCpQtruM0tVuZRBSfjhPqO1dhqyrAxbAdozRKJOqdOsZ8S5
UYY/Oqt09cggVZ8S/PKWFiOCralmySQ57NFt9JKneePf1K5sxpUbPmyydMzwbUBde9Cix22NBocH
5xEyFuJklwDWZkuCszs962P1Szc4sZm7A+0E/ZFhpauw71/8A3v8+QIpWCC4BxrV9KpkZ5PIaBxZ
7su8FRcp1YCeJp/OywKkJglTuamPHpKt7qdtzA9DiOq9CRKZlo84RF/vvE0Q5fYHAvtLruSnNM0m
cYCK7qhKVtgvDyjRB0GR1uZ2hGK0ZiPrx7YuwKO0Dy01aTX5RVGbG5p6WEPZq0uss/kQ+hQk3A6n
1ltUZApo40lQDK4SRV3/vGNFH2QdsD9TdTOO4Z3fipVoIs7MTpEZpUnLnLOG6sxXtN5IvhJWRXFK
Xyt1htHmIHGiKRPuBpE6rrbw/eAkWYLoOl0nyWyLy1v67wmVn8FPKw/QhJ/sK2T53slEd106NrCv
HlujA8CUtFEsMIgIZWeIbZq2kZTeHyfz/i4S99fhpvs+9g51Gqq8wnHImI0yw0Mb2jSFLu385kbz
Fft8mQy9GKXr02HZTF91/hjYfGzb18BObIbAfOBW40m3nJ1Dg18D52M0ZwfXL9bnszvB4fQnPUrg
qw15fxECLeYRqd9x7b9rSpgC7QHsgRlj9GG7U944FZ5mzpZypnOrAqgAjMemOyHPDTadMT03+6c/
ygBMHq4gfNyJHeXwmlZhbsfkS8vqECPq9SXM5bWL+5Ja8XzYQY1z4tQbXDr/LKrNXJ8aVc3J/hc9
7BED8GPXOlAx8SSsBud5J1E3PUXIcE0vNlRLlNGUlAznqMA9yN6pZDvJyUB+bZSwTBFM8fE58CIj
5wZsBZmeI1sUFVnaToFR27C8tmFrdH6IhNv/hyBMSTz1pk+c79CirpotXIrGLkqIn4oTS9Xo9Xnj
F+SxoANHRdzK0dPsCIoZv2hhry7/RT6//SsAc3x26bpo7azlXfvQ567gNBnTjKZUFevW5znpIDcT
IxWwbjEIGKhXMWtjN7k2S/C9c+9KTzxxXGD8k4mX/0Z0geUKU6jYhUUTKB7fIzEZjdYdtBJ3Eixb
dWpI97i+nrhMMHnRq7dCT5vyZORKV5US2cycZ70gultKPsi8OJ0AeoeS91j/WikzL9mfVc80deXX
bffFd9SUNZoacualbW7x8qD3tp0fa27asfMwKRhzphM6EvSGN+1nLgAnflCsmPD5s2wdEVOOvn6b
abYtA3gWwAnjUJ4cZdIzG0u1i84JXKPReEClF+58nHtoq9PborQiAoqUjRj/LmRm8XZBrFlK8D8p
xXru9SjrgkkIaWcZM6ER/KF40po2Xj23/irYCHYQ1JLp3MOh2RrJCAyGc7upwQpyuDFgZYs3mb9e
nSrQMQIejgshvGEehZnSal7Gqm3Nrec6FH5diwm09QSMuN2L4QskYB5cbqnUykzxrA0uWfsAd5IB
bxYYw97BC5AIny+TDpg4YFsrcxNPKJKsOzIhqgTrj8zXTVYi+uXhiKhbVnMdsCFb3A+99fKBVYgf
an6m7sWjqDTTZ1LC00527xb8OID+lz/ADJwY4T3Xm2gnZp/5qUtd9gmP4t5/vz89fjHYYS7kBYLj
DtsMSgQ+1OXYW3wWe5VpVhzpdNNVQG9OXProa6ksNc5+DfRk+hKpOKmjYSWQUec4RnngHxtKqsaQ
YdWmrt2myuRZ4TPYV2pzhQjGn5sAwhqtwGH+G/9UUSOeCdgNk6ZsHYagYT5KbMrgE22djTSeTxkg
Nc0Doe2sLR4tukdLiAZc3XX/Aq9qC3+uIICvn5A4rhuqdQNWqlzDgoOFzzROHwagxrsRZNJNEMnR
46l6NEmHzxwlDSKowP4SopKXIRVTywXms5EaOicKnVVPoCzGO6QGHxjkcCeCyN0Y1ZutBFB4lf7e
pOR+eiQc1S8oMvyPBIAUxOOfIHjAqkdoYCdIAni2AzvrszH7ghL/juLBXc1d1bLlswmuAdB0df6E
31yGTW7imPLrEj2c/qp0xoa/tKrMeBkpdHjXCuBoqR/uGScaDtp2GMyHsk8TGciWc2dr/eLHtmDC
BfHiR5W5RR6yiv4+syV0EgN8u3Sg5G05gGiIi80Wp3es0J6uzuDNFOb7uxaxTAabPHUXJJ2KOsxu
cZrhuNQsI3DY3oVo4OmoQxWyywQypCNTxGgBuyFQMc2FQeUUXYavisWpL6UqGc0aJUWmAKuf14q8
4GeYjcKARp99/TieV2Tg2U9oALRX6+9drMFcxjcIamnsi0um6VKLaX11MK+UvJj+DUlB+xPB7wpi
tzSvoQODjbCR7KMScFv1oCdz5NWWrn4tw4g1mbDs3zycLEDtBKeBo/cM8qDHSRqnh6Jqrcj7xdLF
EcWoWyORs8ycFZRxn33roQ8jwkWF7d93qMZhlZDXlnoDQZFgdhUWVBorucesDlO8A/W9rOnalT4W
5XXJZJS0Q6Mi5aRaF0JsKHfV7FVZPSEeO/AnP8B5IP2MR0SpCgWdnsANuG8F1RA6NNld6UIMETJ5
ND0OvlSi/+IyYvkvBEtaJVAUAl5ib4l1rofRfXk/bumf4spIWe48Ds41P3rMkn1zTU7Ku+P/jRlS
P+9xoJkKQ/VKn3FU9CR0EvyzFfbjc4t9OmbyhYhl0WVCvM3Jzgdt9CVtuwdAFZDVLwzGYzTKxeN8
l4kjpTJeSTWtv7Lytk1sejvGLeBtXg3sDc4/DnYLosCk9HnnNG2k1QbmM53HaU1qSmHV87C+E7zo
7yBDBjT/2bd8P1B1GEX8oxK0sIdy9afx3gc2tc/jJ4euEaKRM7A74PAu6njkY9L2LMpRKS0mnSEf
7LrnJlZ6ex3sG6r0YwNZWKFrlepJ0Zx1YVB32yEQOllKEaxYk+xlxo6EUWdhov3//sfH9Bu89X9J
n5AMEPYhwc6GNCyO016dq3D4nB989WkMDn4/oDXgn4Up3O1RHRzMqk33mcCp3ss8hXITUy7LETLn
xBXC7PJOUpjKwSMLtISMZ41a6Frlg+pWZX4JQQ70qUkfQzy5//sacgktQTGjis0GU6DP2tvWwqwC
EKLJq80TKqHnQyVkd9zd4jzM+Hiytr0xCJRURdMd8JTZqNv+D5mDw0KzbvAA7RWWjEJ+t0Rzsvlk
nWOlVQPghk1ZvrDByU5E3ffj3QZcq9tLEDe2gwJrHfA80fCU6LYBUj9kBxxSTrJ0zM9HmSyNeTWk
HZ5ilup2nFGeKUMzSv2LpTTmmXKY1NufYo61cUDzhPoUNgxEWpQvX5tdrReG0UyXJN7dBZhuNvFW
g80+aUQhlx4BE3EVemtcyW9GYHiMtUQRZhfRM9xPGEGfW7MXqqq+HJWY7xYMGYoeLwdpmRM2ahsZ
V+j/f3eNDhY+BGZy8IiGFsBJY+cwecEfBzIFcXS+LVtDnn45aPqHNS9Wt+N929LJkoLroSSo9I3w
6Hq4T3I2gJIcsM9qa7spHY1hJfrRZIoX5l0FP8EwHof+prm/Isr4saCK08qSwC0RrAve4Bx98zMa
jtug0+JCpZJY7d2rZmEKLy3fuYV0WgV/bmY7KlWZCoLV8+BI8s7ks8XmRK7BVdhK9JCska+QuyDt
dLcifD1TsSP92WO2I8FuUUYVKphnIDSlBz0D6H4tu9llfHqIXjpumZtKNBA4Ziy2Eu7z58KM8arW
I/ALa8KmDWxWrfqRGhlbK9QyNkjFWDdphtdsP0GkskzdeHkx+3WnuXuX+M3xTPvReCgi2WxAr+0k
BZHg/m9Z50cSqGJh+hKlx1BaEHfyFssEpJszOPpVKHQKFBKdnvEM6gloRgAPO+7u4vukNkMjL7zG
Qnc7yJeavn7jm9ALXusy0ytIIWehgZw2dYGYhCaJU8rOKxODNNwUekXh7fKS9mwWCZK/iSzJYEZy
ohUXyl62MYXxkZtLiS5qGuh2E0zug6l4MPb+UwdoVUcFtefTPVwX1NsvZ6i7b/K3z9XzPRs8oONe
D5peix3ObQcs+DP57s1zdhwMR26Ho+Hq8zR3K+z5o5mMmGcRTnQ3Oq0w4My+aQ4auNJV1qemXdC+
GP0i4k6qislbsFDB/nx3BhdfVGXMRwOx/AgVI9+L7q8TF/ArX9pV1e16ZVUF6CRflK7UG7DKMIdy
qxpZmuMgNgbeIyOYvVEg2vX1IRctad8Q62yHUCYan5v9LiBHBGFPuhcf1FbVt8c3tgLGcq7h/s4g
MqDcnnMcUhi+ZDe+sTzJneNXK4LgTYD2levbVGb4RX1wAZ3HHpUXtZ9O8/4hqbd25cqXZeSPBbDd
zltwBkGbC5ijN6UpDrge3Lwj5ZPTIA5pahHbvFr4dowNQ+Y65zDqVvFr65TuIVlwZSo5KWAqy4CP
WMbS4xhW3uSoEUWuQ8HAkI7lVTCrbsG0cpvHaDSx6vGYOVCwYP1QOo7IRcOGHJtJEHPa6gWw4lot
C/Wb5OkCGyZx7ZKEAJ2zYccoSsSlvHcEzEqWBdhJWQToTs93b6Cn1GBkCzEUI3SeDOds7ZrN860y
q9CMF5DD5ijT7DrVVS5h7R6KR3cf05ydOnKNx993dUxaEPEL4fn1xwWtahiG4G+IcHxZTWt8rjpl
s2aI5Q32J7l6MU9jbS/vcIUEdgRLH8X4w7U1OLs/QabgGZ9eCbW6JwBB4BolYt3iGtPIkIIZP1Vc
IagZkIMLPRWxtr6GbLiBROoLtGo7sivXslPSv3lfk7MyhGbp3JPpVFuMqX4BSgHreFaXJHIYcxzQ
l+vb2GSpr0l0hLEUUapNCy7Ip/vPJ1T1tF4AA4gwUGC5I+MeaIfXs2Fp4nZ+nVE6twSL+ML6Jfy4
j9oF+Tgo/0gyo81UKiWlXhzT7slRXOAAmxoeKnx7N2Rxk0Q160eIfSdHNe+uEpbHT4PQ8T8xeN8a
uaCnoqqGaU+oz4P1Fz57jzluvGTpFHjzYIoD9WAU2n1Rf7QC8SkW5aEQ5UiohZ4wHeO7D4gxEVpt
7/UusGDkBlnPASA7A+NT1VaYTcj0Ikg0Tzt1bPKlTL0xswvZpXbZJAuf1WTEpTohoiiRHLLEr2nr
lTgwolv96O6k6tTQfAoV2vBAuIx6wImLwB2h5eq9Z6kb+4n/MnV+0KhaiIRlEK9CflO0PR92PA3b
RH+rlDSJwSIKFJvXeP8OqIrf4hfht+okcbQIv3gkjhyplQ3jXUrEmB3S9PNkBQmXMRlfrMvGpKT2
WAryIWqUUq8iESj9R43KBz+B6JJKMVivW/qz8JYCp2WAgnlmsiA4MI0h2KUdeeZRO7HCjCHFQKya
XTwXV/ye4/U08XGELg8RJk2yKqu8y1GWipGSD7Z6nX2IwPYdkTKxaaPVC0Jw7RlX32Oj3hFU67Oq
mtWitMPEot6WW4VLVYyncwHZRr6LUPoXJb+ZSvYYhfWTEsnnU7MNi35ToRfDbZGDKtlQ9NTK9eel
waPOFF/1DfFwsYFGz6fVRqf+pKa8LxL02amwRCWjLtz5HVF0z/4KL5diYeXG/uL1Dh/6VgmVjVvm
1J25ffAjMrZp0hcbIQ7P61aopD95tBbrjZ6W3P9uOSl1VVKyp674aiZ2wXXe65hAavnu7M6sarCV
ogidqQxIvIp18TMkXfA/nOjBOATvBzQ5HB+o8RXKtpt8JHGnrsbcJICNn7Ko3DEbz/GalxaNwCK8
/xa9r3M8d3MhmGAWkjxPEz29xx+iBlyWuQ2J60FtnGG9sAqO5FvPMiwYDXXbZN7WOUHfNtixOMBX
8H8Kl59vUHW1ifkHv5i/S5W+k/1zgwLyMAB+J2vDL1J7xt25neiH9zr45YUI0ZxXvzDk6l3qL2FZ
1c/3eKngxf9kkKoakAkpcS3d0Ff5YobvPXlD11EK2mCBk+9vPZQxGnylt34qcC2Qqfm4BD2ZB9Rg
FP7i7xw1RpZ2ykHsJ+ATWebun1ULVjLwzyEUPrAfvVKA7VfX5a6I7uV6vZ9OIlaHrHEqUe6bmdtU
6bdCSFmhUA9CEGnZmcINu0cAhDbMDqzEBnNQxi8vSVtUhd5bkHkBYc21983J/klpTYQVkUzfUhwj
yZ3EYZg8QSrKUF4aajcjueDvBs6zaCeCDooopsqjC5EqM1MmN+hHRnnd9+9rBCYT3CZoQNDdxkCB
Q4/NbhtJ4v3M6jmoU4qrbhHemL0vvFPpdFBjk4mx28iWvceqPr1q6+FaG/FyClE61TNKZuEivri+
3WYuqTkBdo729DKbCLkfuqZAhyeZY180IgzEsmTHYhRPJr60zM7WajX9Q75Fa/TOr79EKFc1IphP
WrZ0tIq6z7ERY4N/IF/Vnkf5xUwWVXJDRpm9ZZqWvIWKgNxSwhPF1tdzUKvswFCG/W8DUrsR+1Cc
AtYgbg2yCzlXJTf7R3JxbSgEWKTnWrBpLgCxAF4NNHLfElDo9Xy3avDcAhGohfvqO+CjhsWuTuZE
9cwzmWXRCUFVzJGLDWlTl1ZK/D/oGmsQyBMxZh0AwN+cBdPooUs4BYi+Ayj8HoGSwBJwzdPhXYAO
RSUB1YSGk2cRhAteRfi4QCfKh4A2/GtJUPyFRn5r55JvuGFA9C8P94wZ9U4cEvwXBiaBalshRLdf
F+3yZpsyjyG2mc6SOCeka3rVZXsO0xqCMiNImnyYxj5Gk5a5XYDDVl2T2wQ6aST29pf4Eogs2FyZ
JTplUCWsEsoXM+svLn8wRRsHoNBmJ303XeSNvkwMlEd2uDJwRcbbiFQc4Epbd+prN2cmjpK8H6xT
2FOPbHquz20+xaBK0wIV43b0/KJDC5HBILZ+/ndP0YlCxxTZfRRDgsrJRpUakD/KkO4B4qzU3Umr
3DLCQh3iXbBnC3c5pfMS4aXu3zwGg9DmJ/NP2naWyu9rWumgMh/lOh732rUuemGSPNRf+UscXF8E
vwEP2twVEoSkhj3zbxQjCm2swkrTpiq0WtjmyFLvXkRmNTO54mnrnmXGqlHybWQnBWuC364o5M7+
QPQ1FYyae4N1mcWe+ngh+5bZrcODXMm8OhjOMIaT1kT8CXFKRjZlY+Z1iSKNpiUqlFsYQuYANfq3
do4gKY5pj8jzxivoGLDE3gl7L9bughf30GLX0GX9vGM0ZLyFqCwphAR01JuOzN8eyNJMh4DlhG7i
rNTKJNBavM/t7pie0fwYGN8R4GuFOE0PLlhkQL6mFGfCbxrrqiYFxeaezZVYK1omtHCHYWMT0tNC
H6WB76RYfV+tzqgxdLwbaelDaEy7YgX1U3rysu2tQH1hh5MqjAoFo34smiAKgss1g06gtEYhMH6r
Wj9IsF8b2F8bb+LwtVf9qzZuR/SkA1D23yCTkjIpqgRK3QDw4c1Nth5ElozFDMJL/4omETy6YXmo
66IBrKX49BNnP/PmUkqX7l3H1iyDdwc9n6/waPGGYUWCgK9d0jPcIuV6wbCYc3piLI3bptzQSAEP
bT31oay4r+8301nShkLQpwsaPe6afF3J9OwWiF4bBNZRFuzFT66S/J2ok8S39CrTGAlUax1pNzut
6rOFHULaZAuOskobHT5GVplC8ktyQXW8cxFWw/IAnwWVPLvcMdBsAUOoIpQ2Oy7/R9gs/b5i2pNw
sVnJCK1SuEm+C7UZZPVxPwqMwQIc+5D9qCIOX6Xh+5dMipWKxZm9Gv3EGXeLhMy2COq60kvdBjuQ
crSrhkOb2hQoFus3NTf47VMS2z4kLNZi2Y0xUdTubRe9kg+/LHLvggufKGrht7jemx/bRT0FL7wG
IY1l1uNKerB/2mGsDKby5pqu+thYmq3L0HPEHHVy0Y2j1tKvHDvs/N0G+yOhCRxyzlVq6DD/+9qT
yCdJIxy6QoDjgqtVFQFQv66+wCWDgAHiYotlGAmL4eiCwJWr0Zw0Mij3C99cIaIb6G20szpszRdb
nL1GXzSIEuZJWVOp7qkQ/rGzQMgGvjaemeQVqlpUdH0AJQz4dcFXwdLL/di5967JLuIbVsBlYcTo
BCxYPFti3VXc95PLnCaEHyJ6jV7M3iUSz3dROiFJzj6XXJvyIhxMXtZ9dSSs+tmj1Bva43EJ9bic
yg04a5ecpwx1EWbaoHIti6VX1c7g3Sb8t3yGOGgVpl1/M3xaJrixVsAJOTF9yuayNNKkgT9iNqcj
of7dtP93UZsIFlq7mnL3lf+iwuQuUb/gRWzTYLEBMDKoFsSdb5HfvfqjZYogj/Jt38G5FkfByu06
Wbnn6ypVBMboKLqrCg2AUb0sDMKUEZQhIvw1MQMKtxqlqH0Oi4xOozObBWKFsm/qf86DnOh7SiWS
Z43UjSu9ZumvTZNpZFAccU/sqz4xhRXA0JXrXyVNQ5xAIC12An5/R6VqUm4H/5cc4YymYHQRzO6Z
rQdS3I1psZz0UIrnXcmyXhmJnltpNAD8WSvFJRaGYR6GRtbJcbdZRchuIlxGbRt7ZhenAAiyJzfs
HxJufHMEhDbz/seeaUAgRzJLo+r6KBlVn01tZX8b6TwZmrlQoMohwA6THxHbhiYOVwcgHHE1/3DZ
GaMPKW+w+NgfSJEqSXUIgwnqcatKMRqavWnLtT+xZJv/Nmh8Llw1ba0F1uWr1eGcUx0T41gCQI3b
YEeAezzB7qfqXwO8BHdmAYIkQGrmQts2MNeWsfIlmeKZXdsYcfMuDENBT86524pQ1LtUAiNFP6kB
Al54wfJWyFTUYxSCebyLf3Naj4ZedFwxcp3yWxojQUkZ+7xJw72XN3dIezqfaJR6l06BV5O15TTF
Yd3A8QfQbtod+4aHdnglvUWgZ7yMrlTB8KP/GbwOfQM7acqSOQaXDn0VturHdYOlysQv4yOG7r5d
9N5QcgO3YCms08V9wbnjym/F0IqP+0OwPpDzskH7RAXo27h3Mktx326yTXGq6YkMYw1EN8CTN0xc
L0ZVhm/TOZvfxAnFhHHmFrDIE/FZRboz0c0Ig5eFi22Yhj9tqCxdQL48f5XIMJznchzWmjCHU/KC
gf0Ff8IMdBk8YPgRkSMB9Qr+vgCcSdvZgT99Bgz8D0ULaq5anTh7FmUsg+17kwcC02dOWmJ+dZYE
pNF+vgysoVOtOD9O0JbussPOwVMI6jK+4qNTVYKqgsC+3qUifDNOLLaKUR0tjYB9DyRhwnSDJGKA
EzBP46zqBsXi8xre66GA+KUBr3DXsM6Qa1SqAE0S0vjrETrL7Jg4t1Fw5Lg8SIjY0/aX/e9A3sHZ
jj3LMLbghpb99UvlI5X+fDyfyGJZuV/o24pXGSkpspcLxqTf/mHPQ+ckPsdJAanf65vAXBjqwiaN
I2L/btnsQBBSYLvooKGHINen2Zw3cCQNpHABgLIbO5ve+DeOl/mOdjp2MM28Z4Inhds52dKMTfyL
IR44nDWpOECK1HpTeqKdknu465P1ro5NV2H6ynY5TRLdg+Zhrh0+sRYvytZh8ZPLvUjtUjQxlY+g
zBTl3qWEwMIv6/Uvz4SmaUNxV27UURa6gLoRxfQ/oIdOEA2AQUMJRqBg4x7s1sY/Arql9nQzJ74+
wR/CrD6Ee1YyDb/8aVTjBSvj/K+hOJ4YNNSfv48aa+aj4mKJFNUydwQKzmQ6Z/JG65+QaLZlcs3R
+nOBi222E2Nz3swtho0xP7IGxV5olfgJZYGwEbBbzZhrW5d8skjgpbU+ej5e5iXzaeE5YGIjXKGb
jf2uIitnf6xq7ANUEiT2T8I7dLO6qto7evzqnytIKLE2IhOnR4Mk0jvZIwfcBC33eij1AP98fv2U
gSbIV9i9wPo6I44161FRb2L/M7UwwS2+on+5QWdVL2QoACjwrNlHJALqQiISaYXJElb1Y/XC87O7
fTAbw/nj+FmlbgMPEt7wF+RuM6EfvDWpH9xpxU5XWvpL4vFIZvLD8rUNnIPAFlE5qE/dxoITo3p4
RkzXU5QuNkmOMr65Oo1WwVNwIwxcL9sFJ2X3OWWlbbnVXQr45ARTd3UddUQ4R99XBihbVmsz601R
e98u64xbOfCvF4S7fs2W05gRDQa+IokIKpVulWG3wlTuroYHZdpl4uYJfEA/l5vbrek0lMor6sOR
hWRGk50jpHLuNKxd8E0dnjGAwLbMSLrFAAk6mDhumY47NqEigSNP8VPO7d/PFdbWmWiCxWj0MsWz
WXCPRk5QDwJNap3iuzewCqekh6//+Ws2XQe31eZLw8wTnPGRxaohkDykwBB1bxdz5EEM+im4sw3L
oBwFRQ4ELazlWusM6fC53uuLeQ/Px1BvadWBzKeDmXCd/tNATssCFwD/gx9bXZonMNW2qIN7yTyW
Do749fiUrecVp+cehJVcwUtMUHvwd0WVZcRNMpug2Oxd+JVwQ4czdYyIVRfymEBePMqPvcQLC2cH
b0xnUzB781TFw7ulzivRHFgrvZpyCR+VpTKKvSRoj+1U7PSbkfzOTS6XEZB80lezP6xDdl4wrbff
zolBYnfgUPp426F98+83sHrK7eiZW0xKMmLIYus7dV3y3Ls+6kAVrkANcj2KPvvtHh0Wnxv+hyev
Ii/RQR4xsgqdxIxzfyrB38lW2T29Ssbd2ClnhIjs6rJN1Odc0236cXVS3wnmK7FgtYbpC8QIJ4Qe
ikneklUlV8zt/u18SjMFZCEbQYNxihCk7JQsHaM1sxQiYCZyjt/QlLxMfaGosXBl+FPJj0d+n2n3
I1EfA1TlAclvLkyzYbgHqVA2Rez+odpLLRMzj4RV7pCPDGgV7vmumwtRfl7M1gWOxqJ0njiMGhsO
8dG4K1RmbwNx9xjM+xkYninEqJWnKPCnTKt5VwQVmy4lSDmJz2afJD+Y+/4Eourq5GWYWRp8kQeB
6D+YSECSxmEHA+XqBl45GOvEFD30VlaBBpKWu9dgJAMngRr6MHLdqahdhL58PmpmP+FdSv1+kJc3
3bAhChRU/TE6BSwCRmeu9cdWQ1eNxPIwadIpHSSEUtobQWC8+7OnrY4/aDPmvokxZO/1YL8neLO4
W2XqafHYqkOr0B68RDxeUIfYwCsrJgnMMBsc18w0K6TOs+36TiwxiTBMkQHCQy9GCTkVNZ9edO3c
1D+/O3c01JPKY4MJnwmAK4xj5VDHxm69HdjUiRH4DeQHr/o6WVqPL3S0d1e4Va6l3Lr81ieKxf8a
UgQo5yVa+I4Bm3F8uE/ffNbeIXFtSREfh2ghrvBL0pyb+UDAeluSA3CL3k/2znXaJWAKdjCZSYnd
UTC9rT0nJSoFHKReyqFTW4LrusRMeIlpP60mRaX9nJ0UTzi2lA5HWKivq610QdSQzm3Jaf8BAo+T
bGvYXeepK6SYGruuta+X3dcypLK90OB5JXCIUL2kqpFrEVuGPVghbPnrDLG6GiDnk1T0Aofz8XXH
9Y0p15DWZgtRlRppS4h4Tyxkr/6FEbnjaxSch7Lji7Mby8vNzDt/gDKlCV9T6y025rAWpV9TDjod
Q91wtg5bIgnfMbflNDkFuHiFcIzldSpN91myR27TXfVeQpr7UYjSPG2GTJ5X7M5PkEa26sHOZZph
rW3HVqtPpM7CDxYAkS3NX7bijkC20tU/uUKxb30M4b6i/cf6sYofH9WlxTZHN0ll+mpzZjUx1Ob2
DjAXXIMldI4wkKWHZaM18uRDSTuINFCUz7CAEbyY/aSEOsIYUDb4hnkd+WAD4FOZO4F13aX9P7LB
sxGhSRkUC26aAx+2etvZc8ln+uqBbO1PVnC85JLRUvJs3Bz8nn56ydIB4OhQfR0r11t/PgI4xZTE
MTePQCrREr/h73JQxPTwMmAN6ixFOKuFGJFLhRXGqY3WELoN8BIALPocOBbIxLWN1Q+eoX5R1gJ2
rGpQ7rXN9yBuOyrKE2TC1DFLahU/i3XVXMs8licLhJtu1JqApeYAfkB00kwo3yMMRNIeQ24ZwSHZ
PAQo2/KsYZNYpgBdY44ir3pIIMVgxnZpmHj7rAEiAhXXFd8d5j9FfgZtXO/YWd428VEDhWv5QsbL
xNAKnAbiLygZRlyiszVeI7hIZ+x5JfKe3uWQBdHRdJOIkxghPoaR8gsw71XV66/baVENiV4CFENW
fQz78VUCm58TAsPfa2fzHQkr0CkuM3AMsDMDhDGl+8p/7VhHboxDQtia70SWBLyBPv2G8yYk3F2c
4MCu+ehLkPbYjfjUMktOQAn5/oCjpN+5Tvcs4h/Y61/I8KVeoVMF8IjzSCnaNzmql5B2t8ZXw7Ra
sU7VgKhT3pzIldJ8YufrSM0vdcaG3O0T1Rew+4qubyw+Q4iGZiEA+Cw5kssE+J1i/SVoGRfkFLkM
XuRiYfCQgxL8CrJbz6weYo1qNtNof7D4GCb6ErfAhtY5Q2b5YnE3HtLJ7H9GR2d4yj8JnVc6Ivgy
eZYO4U7qxddU8dhHzXVKLhSlTF/qpUdEpREQRNpkraxXjdiYZ2aVgrQtkSfB7vwjZ0clZ/LXzqa6
iR+xqD41+b4bj40+r3uQCJhdSowEUmPeB7NjLBhFcNiOci+9djDCa4DuCyV2R5St9RDEQg5+HrcG
SDICnAT1fvH+MAyNFjsIuI3zJCtV1OUnDj9TrIhbBZwPSZjFC9EVc1gT6NcT5ZRH3mGTmVkv1OF+
KxMvz+Ec89bqc5tb8k8qjNWUwD9v30ukZo9vSkRiXJ1DN3OHWCpA5y9tO4OdSzmcOLUER0fmNbhW
2z5rh3wtBL/onjTc4HOq79yyByrrKXGsGgGdjWSeATJz4gY0W+qHx4Uvdq+HRYc558I49Bqb6hB0
oIJspFusogy++N/g7KQY1WtnOqji3SCEWB6wDB05KJZ7hmvo7TmaHpO2DgSz1lY6Mp6kcv4H/npv
KAZYsQL+U9TqPkZ/1oh7d+qqiqkoS+x8kTnFE0KQjiAQ4+Sxt2kTu9rg+eHFVN0noX2uBpVyaaDN
wZXjwgUHgR7dHPZrvtHiXax3kRFytpeAUJxhqNJwIwsuC95pQbiZxhgv+zy9nbnTLWz881E+6P3N
9IgBl7i3xbcm9NDcwuWKWh2V+HacdiosczRyYyVUQ3Z9htpeXaHxF34KdVssx85QxwbGDxrGa9HZ
qDlOsMZeW5ZUAqvMGVmsp5/dwcBGdHEjAxI+8udU3QOjcU012KHvd9MlnhhKBp8qFlIi+ArhP273
qGU/FxwLeHQCaIwQTXLu2MQBXGCzn0fP/o7npaaP1ukYulHEApnaBn3h9SFgzuwZk4rr6TybUlyA
QwW47/vhQVQiS3l9D1UyO5cdjuwgqx40Bs5AMyEaKB7J3ffIEQPRIoUFqh7bDHTtU0N5WJrpS/AF
0+3qa8lGfywIvXFd1AZ+LgS6ZagKQFC0/2HWdiVKqC0bgJiQHl+1DfRjjHHP8wettrpZqt5CQOAK
Oka6HfsubHaZf/HCK3yr64MmZG0pFKRSAMGwqaK7MKzLZs3QTXoeTLOMhCrU/gH8s/Jg/X62iqj0
/ZggvhMkn4Fram0tF+Rm2aoj+hM106tOh6Z9qy799jCoVOSL+IIATy0AkXa81o6WCN057lBAZbu3
oL7b5BdGyC9V9riev27aj/Vi13fnMXSqI2E0N/iKMYKL5o4RVxDioczgjEztwOd/JG/K5PsRNNe0
nBA9hLKEqYI551j6iZCkWpgMECJk1rXgb5/uz3a6I/GGlJu1v6LqJQ5H0QOAqhWexjlg6P+70Qq2
FaTYFVJjT57lAFIjsD5jm47Ak275wAv1d02EcW760/z3PWAKm5tsRcBSi1Yg9bCbKILRw5DKVzW/
NCT4PSNLaPhftNK4BuJ42SmkujJnnX1v0P2nHF8B7mnAlUpsGSFy5xTSqEXYm5sI2TF2UUlY99LP
jfKRDHyYdsKMBa77xETCiuA1lviLdkG71sfQcRHLl0CVbth3nzNDNiegJIqAC5G468FMflXQjSHZ
8LaBgmSFK+t2NwkpXUBEmIoxv7NzLy5QVrh5KysTHhFJD0G/KNCSO4UaDGqYH0b2NzOExE9dySaE
hdA/DpGkYvS4Qjqd4RmljJ8ybQIjrjzjcXr9751/f7q7mfxiI8PKkYiV9HLVw4nP3XiUoNXZmJBW
6+bZbQxErtA3xrFEKaCEdJE54gA6RuLYnO/jYLoybuYq0+QnDXIEFZibpzN5ugAlqiq+xGMN8o2F
bKTBa1rhFu+6glulKCV4bWEK+Vn2G4iRmTgnFgi7lJN6FYk2tcc9/xnWccNCYTCldw7dQPuIh+MZ
lIGdU4w8f+P3ImPPGiPImUe5h4OUFtb+Hfd02aowjeBx33QgfUBASkjVENnkhTsgJRBubLqk3O22
ZLBkuKTt3DJn5Kd2p+yaXea1Q8RB/0fAU6jCdwKcZo6tRVvf87nMYbGLa3WhPKbCbiHdxQGXbLky
VIP8NoubCnQZKPfNhtESgt4ANjVeBTiUfOZB9HCnECEQYhdAekents1WHgpmv1NuLd9lUrbEdVqt
TREM6D9PegOhYYjmI3iVuYKcG4MvXyvFzfc1m7R0rtSM+7nWXM8N84daunegl8DqM1Gb2i6sFozp
U4FUair/uwXNa09+mGhiFg1bmaFzkhB4ri4NVjxIFiCf1fRryo9MvX9QHmqKymCb71hy7IarIE0v
B1T274QkqJ8O5DXsCC9CUQttRJFOKx6DcefmCECasM7OaYsJEzKvxvPrEvrQg/SN4yqAMn/As3SV
/YDFLt7320q5NcADtPfoweDn/TgoLlrYSbqCSF7blPSp21b31/9x5lDUgd4cWA+scHPzG355hZI1
6KcYTQiAD5yPSnoWDGLHr/H1oHK7+n+h2sc1jfwYzXvBm/ZGRcEH14sNokZY5Sz8XCrSH/ZW4KXK
jRvVDmq382yxmwH+1uVIjpwxjvvqWPPkGh288MhX55SR0sWGfG5X9cgK5aAVTMSrP/bI2s6lkNUk
E91SuxYxk/5mP5V221HMRzLK3iYRwTIE7+pORGOKqnp5CjM2H285D5nmg6xil34pRZLbzAoOytmV
E0D2ZmMIndrZBHTRqCvUkM5e3Qm32e1I7NqMkMPopCahD8ob8zqoYWctET4IRg96/MPsBZeXbimx
Udsk+wDWF5yS36ysHmZxdOOP7xCGFFTkxbe0WDeOCRmRheR2c5uVQcCqW1N4C8P0/VrOYshvSDj7
dfI1clIYlLmPFcgDueRp3G+QVeWizbnvWlhClpxhG6pkij7rFNTlLXcIqfNcCfmgAWG1ODrBoGne
DBrpgZSAAWrTExkluCaHuQ5Q1sBVH13S++Vg2oGKqsM+gOhN2PKSoCzr1qGuPHuzDYefaKIzOeMX
w6MLNZ8t0Ho0Zbo+1CWObQHUv5e5sf2ocqK+QZ0QreB2rMH8CxJLDRA8YS7dwPSU4/xGddH3crtj
JOJbW2lK1AIKatRW1dRSh36TsxTdrpZUdsJxJjh2zkfSuSImw04P2DBcyir4NRaz6R5B0XM1vz1V
aOaqZOnBm+iiq3EheqhGcUYTiUYSMgyHhb9yfKuDyBtcmWB+3KKQxy+GOOdtz+f534HOWAriRmwm
+igjNd10gmxIohh99kesYXO4kDc021OREXkfSz4L2LIE5zA0rG+mnzjH5zQNtSZJ4+0940voXKLv
m33KioWK1oQvGQtHtN5C5TmM1Bv0to5UPQg4YV5kqrqGNNSbJ1dQQfJBKTvcDX87sUX5SZ7LFMfZ
slQq7p/5wpVKZNjwl/mJcu+Y+WBGO8XJSYL2Oj7dnwVXa4E/NrgUBUr0IntDaWCTBvsv80cmGbUq
v7x0x4BhhPQFHeeviW5VpOZEUAOAQewUy1Ja9yu9eFDvQNt13i9Wi/vegw6HnEvcgeHzvmxbGO8Z
BN/+I6+L3C5wrzKo5XLItwqctKQ4SFpoRLyPFCFoezzAsTG56O92trPB+0iF/DGer66KRmcoN6hA
HgvI0aIJF/uDZdrZe8R8kQvFtKXaaqQcSBiFu2J/S/0UYSHpauGEhdvf/hT5GegMDYBPYaYOp4Mq
0TJeU6S8wIKQgHTdrXh93yjgAx4RKpl5jcAGJLYexW/oITwoOFM7vc2F3rVSYj+U6zSMDMeV2SL1
rwgXjxRgRuFzajF+u7pwkVclhW0kbnW+LtmaeoCY4isEo6hin9sCa86KzFp2zqDCpbAyLvNx8moQ
oZog1+JNvbUXx+rXIjLR+EbS9TW8A3UKgnNzgeozGx79PNUTBo9ViCfKjNOvPwI+qVD97MsvtAw0
NC2i+PYdSzhFcYmXa0E82+topMLSJuTFkzfmDCvhqOsKt6c+YF2ztAbxN80sDC5LQSlTqzzdeTGI
3oZKSTkWQoWdbK8yK4kWoLxnEfoPfOPOiK2Dy64GFBnUQr+U1Hk0AEOAGDTGRkTZnaHztYBz6+5Y
daU59xyKzpWGAP59ghe1LUL0WO4S6hzxkuQqobfVPxTRRz9x6AS3KoYNTML+Vk3QAq+NqTuorv33
ISL203uh12G8sYBdecR0Q9u976nDloraStvHUMRGNzh9RN98ioJznS82GEQ1MGpkAG9TDgX9vKds
dc1cOZ9mGQsXeUhHWq+B0h/DkuBAV/VykN02dxTGykkDq/PmkAl66yk5BliUW3aQbUT00ajKPQAf
J982+GoWpg5BInwHhh+6Xelv2aLFz71rQK5te7pouKegARRrQKbQgpVNgQ3MAJ8+ENdpuTH4ZFS1
9NXBeNDXAOiPCemF4h+VBBluZiN/EUqcHTxUWYSTDItJZIsUZUwzq/7vbbjuCSlRQQcB7YCazSt5
uGhe+Z8GOEvpex2gETKS2e8vrM6qXjydSV/lKYYyYecIzxHsG7rdn4uZGWBoZxY4CMpJrS9nvncc
6ltwcCyMFXgWqajeSJu5IFv7s2FFtWhXMjaOEm8lFGMVVujqWWnuvQ95cOIuXsbBSTP+Y+UKk0Cd
+jQ3BX4SkLhIg1/wKwRrQCZ8GJK3ZOiTCbs5wKIJ76sGt8onTCv4pNGz8SqHfVZwJrjM/LQgNard
gZHWouDF1bas3w3uyxCMNCtchRrdVuAZoE+tn9yU2n14G9abVjxsWg3FVafGSwKJlcSN5jQwkJ77
Fd345eOZUUpPUPQzpjtDn9E/fWyzxj+MQ2e5oXUUL3vgb0xitsaatCgpqsp1fNkosBx/unPL1IPs
iLURC8OpOzPoLG3CLmcKGaw9CNSqJH5w11VbJ6vMv91/TPvr0Z1ydENiK9rdNabpzorF4hgDuOT9
gSkUOL6ALwoo3TFDS82ATKfrZE15npewxJUDsDzIdQDa55PQpJ7yzmDeaohcw6//CSGQzVoRu0V0
Bzc9rUfX4AMxAJy5hR1LPCLEZB7iGKilGeVI863AYGgtcRkWXR4Sc+CMSlXASDntLiMI8xL4aBqC
1Q2rpVtZ6n4/rEUWnz9LGMxqh74GfZ0hpGBxIzf8ZYY555vOgycGystwAmuBBwjLdp0p7W/aKTSJ
0EnO1+brafVqaNmZrCi+U5hhgwMUuxof1mrIpqWZ0aRKxUauaSDmU3M4JnpZBoBczvr/nKRtcB6E
mEBLlJp65ndpFD0Qbh1Prr3DRcXahU/Cc1T/e8Hh0Pa0CLG8aIQJcYfgoA4ELn2vke5FHJY1JWfi
5lGwOhDc7ET2/2LPStkddt1NhIw7FNBn7FLIMkxedrrV44DVHPN0LWRB2XJEoEsoPtJDSjhc2qPI
1svANJ+MtpKByu42nzLA2xRMC5ZHAyKNwC0jfKMl6h02VtiAEM7sbO1CgP7Cz7nBObvcm9xhE+Od
whnAgKyxIELagARbByEY2K5qiBBn3zgCudzcqx6m+ktk9hICAnKTggSNEwY7YUzXkeaMNpvXy/cD
zAWAnpJLcd0FhdFKQ6ILauet90WuUShSCJObCU+9H7+iR9ZIlA3yqJJEkkZgnceUMV9XHaJBtWat
uS4CPbhOFgZwzAIgDx/W4hfD1CL3Kw6fAuqC41sPNwyvpbHg6mBMXvnQXJN3Puz7AwbaHoJkEhj0
+fyLb0XXgUZ+IIgwsI28RIbItejK7QZVe2q2l2Ti6mV/2AQ15xooonhxuOcvb8j1jALa7nm5zkNf
91aXGJxQ9hyzIwOxtDYdevi3lvKDJ7xIdtMgzw4CU7NoLgWeiTV0vgGKJGBK+uioenJOMBUtBA0F
NhkGW56yaRCtaV5/vdist1raErLmFd6XsXl6wdBmkdy9BxKvdKr9bG0yGTwNxA6GWEjEOvnq6kYW
vQtw7GLXVrOUTH23qwpiqHiQkh56ldVOk7QvFyDcimKwaCQc3vzrchmAtebMcEYzwsjE9FXZTkq9
25YYnKOY9GvMDJprEohz3sr6CoiFSttW1SRt8MziAxZHkh9McjiI6uXvo9gq1ekj+PCDsxt7mEPk
sIuY6YxQodlE6MKjepPM3m/MaEvh9+B+nNPF6atmbaMK9hnq6WuMkB/1zWa2N8TUgSbCvseNnpnk
sNNvvo/R+c7ykcC/L3wFx4NQAAXOn6C2FsQ5m4xp+uF+uLBru6Y74skopXCHfMfvdHhTDAdeFefR
nEWP4PpVX1WkAdpud7lSkZUrwkgetRDlBLt4S0R8mGC7nolVuR2IAaoYv8ABagYjT0ZwnlH8PKhy
vJ5UKkT+4spDDN0Ccg8oH3yPagiIkyQ67j7mM3dID++BXOJuDev0dxOCsjMjSrCRHhWjICzBGKXv
QKL1PXR9TMSLt80vLXGeilQC28JFVRXd641Uze0qH3skyGdn+QSi6364dBK+IAg6F/KR3ruoa++f
KLzwuVJeOs4Pnla1BjrsA3o0KylbhjuKKXisTJ0Ha5J60srsGkD5rzFTuwVTh0TGUdCDDklpyNNW
XH41d9YnpejT9+63VrN4CApvE2jZUnkcrceVkA0HUJo/UOZCAnARWybmw+9U+eMlYVm1Oo8QfYyo
ASIUfJ7vklOvhVRAuJ9qK7LnPCiKfptJJp2U4gaICnW9vZW6fvtmB01uJcVEyD3hkRsRfRt5ZbmE
/jZP5Fs62kxeiPiGcUXO4MkTcxxYKrEEf/XIkqnfxzfIiupt6AMmMzN4rZ/s8JwvQGEbTFqiULAl
el3NHudjFsakQDDzVgXZNTTgpUvaE/ofNXClHRGbnyr8K7zE/Ij6iwALmN+K6I6wEfBxtcUKiyYg
PFf5z5pWr1gdetQDClFyYPc5hOgrf7U4M9TiDScQqzzd9E5BasbFS2crdUBm7ndW0t1vYznDCmZ7
k32mM5fg/E8uHGAnsFqVHZB/Dt4vDKKVSpBUTPjKU9+ldvo2ymv9cU7tGHSBoW7939ce+mD5B9ad
a6pCWNJy+BnVQkw9c+AsI41t3+GKldcMx9EZ6jErn7eaxmikul5oJKRy6BIft4TOKfC1M6GeDUAZ
EHWz7s9CaswFJQg1bQK0u86sStEouAFZo/gNndsIKO2Zv15TXHLfkb/fnlS7k/j6iG4kgaba+n1w
DajC9+wFsfJbice+FhPXuhFltNI5kBE/cAheAKzDOdgodLmPVuUxI6wKSJTEmTqwygjW1bxfpnxJ
QwFb/DJT+bwbtEsgiAHJtR60jHL3LpTzjT2S4IAhxzQaGeg486FrzOdsbLiAKMCC+OTjmHCaaxrp
8FsMuAY+blLJEmVAohUUYTzTk8hyjUnO1ruL3pwYt41uUPipmobSaBMxjnCLtLXdAcksEoU/dvnO
QqUJlH0VTYPnyByoxZj3rDaT4W7xgPozOGscAYGyWof4Ky0X7plzy1Tl7Mo4iA8Q/PjQ3o8d7h9C
4kXPlv+mXnbcpzyfE5bBKyy/8m1a7Xvu/0q9C0voHzR5kcclXhdiScF8L1CJUkdnGtDxdkBe2KR3
158bPHWxT1ptum9ZmWFBUUxIXVZoImkfv6iGFjqK4vLVRXSBjfT3rGMD9PygWGdeyBOd3Py8+VqH
UZQvSZzpjk4IoVS7R0HJeLFbNpnCUyiO55/wBn2/UBf90tX+QUvIRmN3B0HnWGeBGCtL5vCdp6PE
E9jtTcjcjnOWtlfZjX3DLt0QsFNwswDN/asBxdyfZbMYaVO5qfrDTKAQkjYi4n8tvmhLaRgYMac7
jrQfh08nj9YP+qQH8GVtr4o6edmX1awUA5EoCdyfBg46tlcLuScK0a10TnIfdJz46Qrr8TLCIUyH
Bxqfwa1ChZMqwnIWo6HI0YE4+735Lmgrl9sIyyrBv6AAM5EdaKD2vnn8DNn3CopcEgwau87KmPQ7
GiYoRTPvt9/AuXDikMBbU/vBTvbxpr3B3/oC3yboxKcbaio1XhBIgMmSA51XB3HDZtztWp6JuYdm
RliAaz7DRvy9sWUoiHokyfyBEhmhdguMrsBbtGWmddJ1pQqjPYvvaEgzuqMvVOjUeIvWF1mmPcbY
wCD+ovXxmawKXVCaBxHAqdwOY3fRuMbN/3rDqAHRXicGovDyOGAKYgEuyIYE6+AJv1/DRDUidZzu
IPHRvm4/wAwJUm3op63uCCs2COU0cM1zhyulUGLlgigW0pQay4s/kqki9jGawNGcpVNUDN7gwbBF
PTC6Kay9myhr/eqPSqlix55oaBkP1o97vzCAZeAKwqlxswz0cxlIVvQLN2aNKukeCN2750DtinOw
DuKlKFhirdcTyrVaLfV85C1OLCOxK7RGQyeFMCtjDOYIsDYtWt1x154oWOTyX3XYemMg5OuNrHrT
LDoMQ8eDwESsZY865RaOCDcXr+/7pf7CDEZ3Eg5F9eavxXATOWNzpeFP2R+voHwnTVXOdV0nR9uc
K4+rADaq8pnbogSYWpSoYFueDq2GPWDNWsh5BLQqc2dwkna4mhpaqbuk9/iua75i5+MeNmmKItJ2
IznRY7KhkS0xOjDn3rxmrM5AHgwNGKuc72nexianE4BA65PadwNQhDPpzjjmiGlMFQh/GfKmh/nW
wT/r1CXsgfo4+kxCP1FxMSWr/qfuEpGbzR6nYVHKrjgbihZ40cjupWHkPfSLqVHd4MHaoHwsd1RU
tVdd4i0+9XSmn7ZEVt2tkPiJ1FWI0viXy1tiQYpqIEBQlHVFM0XdZxal2UyO8HPF2wMMS1CJzd6/
7M8tFuFQXJtcKqVxhVNz/Q1TEFihwokaNY/MoP8oU1lPfYy7phMcUTNDa4uQ5QT6xJ1XxLAR45lR
SqHPdWzIYggsKZPOT4+3Ir8zhMVqRVtZLROeHbPHWPOOmKZgBz9vxOFSppLGC4IA3JSpc9od7LI8
HCAG7PBQPzbv9JKIlTZE9DWtBzndUeWj6P28hEB/4fGSXk6xGiTTbE0LXzK5mMIj6KXoFla5ARK3
U2Fie8a2wnAOc0qp8KpLxxOUTfLQsoAmpu6Zo15QpYi+cf8ys3bP0SVs7a8lxW9M9SkshgqatqCX
eadlh/lTD+lHplu+s0a9CoXXmqeEapD4SrntIpLS7O2lWqRChqNn/HJ6CU3BG7TUUelVp+f8ghv+
l379Xk/9EhXrZObXmE52H93XZGFWI0O1/MfA2SOpKLTuippF2Q0Kz3arVjtcpuWXuilLQOp2wECJ
rfMyzNA7cp7hA1EDCImxTc+dEc5YOCE0ft1F+WAvVGpw5/pLVOlZbeSN6tVzuI2AGUGDrgt/82K4
+KnPrGAmqC4yNssyEyJ8/tMC0YsZp7kuBZG23+9i+F7rJrh6cVe4tN7c+8BSTYnyVjneg1ADl8Ow
/RKvtIf4G+01woXoHcfGv3CKut5OB7FZ7C53mi1b4+1IWNUykF0jkysIVSJqMA/NruibRmIiwxaS
8Xw5NUO9Z0zauQRXxWjV2xk6lKNWJCqtRjDjOIW++ZxNHucYI7iqB1KtrvM1f25ozt5X8JtsgaQK
6uIzAwuhT06mtaK4QzIi2sZQsGYzi5lbScZ+9nYjDkuXlWDKJHVdYm5Kk1KUw0OyVbn7fGMqF9nP
Nlk7DPf0SVAhb9PYm9U9tNf0Yp2a7aYjWkiKE1jrI/ZcLRFMgAgJj/YlFfICB04RR7wekgtPCnJN
mhUhidEBa19nhMHtPqrDsotczOZvfrAzOJAJbRcO1/SkMtrvd6sPsl+zEZbxk1FZYFX2K3CjjdT3
ERfZxOKzw9exELoycT+oosWTfRi5R+xchGrYnSbO4eNHKpw6focP0A9jDH0QGzV4/kpuZkyjQGVs
wWZY2LumOFOfNDFMjq9ZfLQh9l38kpHkCno2dK0zsKh8tD8zXg3L9i1V3h1kp+9GhcaQuYzkuBC4
T/DFrqlf3oPXIuhQ/dNDgqkdL5fV0LcKPe9EI2woh76I8y3P2zIUCvhOleD2D0w+1PENsuOLXPhc
E/EcKj6MvA6Hj8tyukpUEIBEWOr0M0gNzcvgY1BwqUtMV+F8JZtvPdpFtJLODEn/hVTwKJvGHaFH
vxoXKqYXHib9CLmhd/IoToi8Ep1/taMDWB/dxspDN9TCSMO0vw/F4Xmvxb97Y74l9sXCsrx5eVn2
VMAcCw2AwFMYmnxvXSjeLOKcb2cA/iArT5hkLir9kJyM/Ny9f55L8vNrH3/x6cCDluqYlX2H/cUs
EVQp+4ZigQyc6TdeFTOFD/zGwNLvvdxz48cGSJgyH57svG4yXQwF9yPG3OEClbaLGrYTmRAj6Bs8
XxL9L1m49VR2WG1MpxvBkNqJ7/rrlZCLIHOy+qOtOejXBicB8OJu54dO3GeRS11f+rJVstC7Ma2w
iIoPVqdhWdEngF1P4vqoSNEQx9sUxDrAAUnJsNR+OfhIIiJiMNF9zlf1s+nQv5nky7gEaHxAxbiq
GWKQDFyuePqairkx+FnJ9T/ZKR4zLou9BAWTq8zTx0Hctq03AaY7ogIAbjOaZBFnuPLC1NUItuYW
3REoLVnpz/UtFlXimrGnGfY6vqVtDL/64SwNeK0oRXGz3lpbSc2wRkHGgHy7xZUrK3hLmxCXFEMK
erRkmWGE52UsUkpPe09Q9k7ZVTqfB++VtpEu6zxauM8bpoZTsjOBSrMG+ulRptp3R8R+38xiBq6L
0ueUHzXHdjAXJuYRDr7oa2ZnEraeP/6HFipJH0l2jvvBN8GUW/tdoO26/hxRsg7CZMpNiyJ0TUby
H8AgA4Ly/TDkMJDH6geiGu79JNVcM/MPTTFYMuCzMMaUMQN7H9GnW2klM85P6cIY76zJkHV9N91r
p5esdnHVQVMa9IbwwSqTQUexZLEyq3dc8G0vOeAj5eeF3y3PE2B6EzyRbh+f57TZ0OkL/O78WWIP
EpeISJM3JlfvephdQcJJZNAAu+3bBYrgzksHFZfKXrl+O0OIZ2k5/kwRxjg6mF8/swWVA8670XbU
D6WUPfPdYUDE/ecwh8VipesooQk95wRmxU7Iy4+bcROZHGxAWVDVlGdzRhDPwXN1Fbs8qWx+Pc06
8vTk/WBttNpR6fwRMcP668aq07hs7BSAFnknEUjjqo04QQioWw9mzTGMyfcm+9LRZczq1b7JMtPB
V+kBDiNHuG7j9rbc27AzBuGq3EcU5gOilt3lSMBDkderDB6fYnUoA3BVLVCaih+Xvn8ooBxocZp1
xcI3c/7jodwcnXYMt1bsD4fhIKYIiN7jMnZyfhe1o3MpBcEY5OBL3nJDNJkc0Pyg/+YEQgc34GSH
qfWpgBu7hmc0G8a74v7840LPuMX4CXpXE26GWJeN9nTClfZRItbbG3Zn8Fmy+oCsssehECQG+3Mb
1q6yPXhAIx6VEZ76LPFQxgh2VjnwvOLbHELL9b7srEFugNhVhCdBlObddX//5sXR78vuVYA4FO7F
B7w86ULyPN6OLPj18HRPl4YqXd9xWZvMdDyoT7Jflu3hqofpcvcG58fy2rctxeuAMp+q89o1sjM4
UCYwwdqIaXwKep5XV6SXqdOH7LtPBjG58mcQCPaNMCyZ7RKA/1EqqRK4z3VFzHyE6hDSMObxerMx
0bQSyG0CrzfkXPhVX8u7bAzrlwjTZmOZIM8l380ArC4M58ZyNjYUkFJjfFUVVl8STs4Cv18hB6sD
9R1siY3gSeTk8lYU3xrmv1Ai4KtmCae/k0xTmIqT01rkaph+S2Uf4Mgv0oud6KP274X+AV30O9yi
mRmhNZH9tibT8/Zhzr2ZriD79ma2wNpMhDXCFIvPuWN/2+sKao0s1taksd8lPaIK+zhOcHHnOUAR
mSGpVaWpIHQzhP2Vc5uYXRVMr68VPeTQy27G98d7NUlSrT+9E2vNS8j9g2mfajUsXFpFvVVXWdVx
j+1sE2jfJDsQDIpbA7J+zWPCROlBnPpBu5cCErFknwecX35LOTr0IKTcL5y9otbgnLXiogHExQAG
m3WwjT6GtEVL7ggtOee3OXGRfXKZhqsGAcr+6DrYelpS3XPdp/N4pNxkk8l3KQ5vYsc4tJ6pp1xw
/mDJ/SUn6koNBv0tQk0dpkQbJUDOMWAECvYDWlPu+K4CDmCTNxILu61J1hXG9h5H/VcWrA0ESCrI
aO7XGTTUbW1un17lhxqxUFZhW4cfL/S3yhQIx/8XGRyg0GTcJLeOOiyRWlHwu4isdO5LLzjQppIt
idCfurjRwg4EBsz3t/PG7xOYFAlnsd9VK50dIzaIdl4GtSawMwnf2bVJj8Ql8EPxp44gqGywXphi
5yisG9I0Yf665zxw1MVHuILPStQJNbFFGRnv8qawpH/jmhamAF9QDZZmxCZ5s0hXhY2qojmcG9Hk
26sEOMn3vU1b7BsKQ1CEjPrV6JjSKSY/1rrtBLnATW7ThtqV9AVwJrtg/81EbbPxsigitHOmF4zE
SDdmvdTkGBOmixuK4JUHXhpBCKirb/N3pZC75deh3uXShVlSDms2EXcqN4SDUptdNi/xZ7EEATs7
O5QQFBX/IYVIsUcoY6B0Q1SueBmKbnGP6cQ490d+OUiXg06gKpgPMpLE2q676lDWyDvbTyhcw14b
nghNneAQzkStd/4RT5NsIH0hrrMYepx3suc8Y6G/fquWg8VboEF1y0HS/fdlZh3cqhk8X02sSz3g
5Bquh/NMCJUBbERd2HCIZDyeZ/tqZU0lWSxI8h8r0KMLz8sa88jh1TNhFJH2BasNFRSvE2bXI/B1
36xvUHicb6lFpEpQwSQLSpfBU4lS9JPlfpLZvZq7evRMtzHXqbYkvt+qBYnoBK5TvJBgpPb2DUH9
P+e+klRcp8Nt8MzWVZOuzPNxJTj9cNXtAx/EXzHdwnWCan4sTLQyzyqj16vB/iWZAeOXtmi8DKdl
YhvlQaTHS5Q0blWjY6dOIvcPTjdDtzP1wMVJVXEli8GmDyUfIwXv+zvnPevtPCDmitYuKZLrsla5
uovzlEbpWNPLx2g+h0qaWRIonxzmxxWvOAe1/5y7oYN5mz9yhd3ySVxkiBxSxXSyX3qmMdM5WStw
dIaHca3oh9aLd9JtjANxIRbgJaIQw2LkIw/IftWHXZVg650+aqZRPB8B44C75c+YMWiK3VV/wajb
3khWMCL9oDh6rlFRSaOfYfb7sw9u9AZH5gTtO3wO9Ve5FN/xg/2+52LSF8bXyP0BQmXEclCNBcL9
UWBahlMBwuCqsYGgRbaiXcf0pPAP4NauFdV5shIIWuIRrWQmos3IbSg1V4W84LhilZGSoAwQ7khU
YNe+4PvzJ/jJ5KK+d6W25DNF2G8k4Ly4wAHpvI7ASU1BAsVV11WBcmDdQXuXOrLQcq8EBhQZy2FI
m1D9/Ndpa9eLUwadQR0JR3NBMJan0MyIqaH0unq0RrWnv3XQcVi6yZ1c/XNve/4ic/B4pJ3iNEhe
WL/rHT1TFVt/8Peb6wFs0lYLrXXnRe3Je1Lxsv9I6MuLRCU3nLa3BXoxWs1HJ0kwwfZq5rKcFDRq
ial3bAc+W+ugs6hw1T//LKEkiOiVVeCJ6Ze/gWV6u9Lqqswgo0y/rSDV+/w9dQCeVzeXW2WhQ7ja
9AjY66o2LPKuunO1SQRtcBOm5d4jZXSAr9ebBF8U8HTy/NwFr4u1ypH9Wmp86f7DuGuMxH7Mn+EH
6xX9Lw9QwKe+EY75T4fzttsVTaYcRfJRC1tHpL1gl6t2QhwZ1Lu+KP5XBI7KfESh+mUNY4TRmjot
fn1D1BMvVBF0pGIYJ+sTADNmU3um9HqD1rRS4+cRZiPlKsmlNdBthCWrzd/awvlkaW1+ctLeZwwB
BP+N8O7gZNBHIVKA//p0xmXPNj9+XkDlbSNCWKM8LExbaajlM+P/vrnW6KC225y8IlgfAnoaTcJ5
KiaCtqf4DCoE54oQkxl5RGOlkgAJOp7plgUd4yWyGpqMQecb98hBqBWzB1uq/eNShMuOLb2qBtJJ
/A815CF2nSrViAy1jfLPwhjExwfWLt/HCgrsaVoS8rMUsViYmvOrk8ofdMv4gcw7yRtaXEnUexsu
88VaU4fdo1u494OR8rAYXHvbbe49gX4BUTVERngBQkixJyEgJr6lSMdGvZMsOfqDGfIyY1V7yFOz
KnIyNE2bUMjpvAws42yvM7BGnCPMARdVczVuuP2C44eTpDT3bK2vf4JL/olO8GeBjdMUQTTUqKb/
zH/4umnWqzvup9c4w4s2sqQqSP4O1VtBId60bm5toM7n5IZ3sPVdgZgcUu/O/DkLCKj487f7p/7h
RF0HanKPh4FSPWRidceKpzK5qhEk8bA5RuEde++g1ezp5s/I1E6TRrVAZAyOA4pbg6Qq1oPShOQD
/lBDAlv8BldVpZIrZaoUrBdFCWy4nej/10aPmfnDj52LJNY4GX6Ug7Lb3iUIjHHkL7hX6a8QZROh
bFnaWwkKE6QC3QwSuV7QPgWVKUoJNsg/U8OvFSvPXxt1F/OPvfBbhOOK1Tj4Fc7S8Dg+ymGZ7tkQ
RJZi5S84AU5xPY6QzrPrFD4xdbzPfHalenjRKwwNy2BW9fnYpRBa79MCFOeynprtInyzq9reu7ry
JFHiOJzRGlSGoyXVUyjUbxQVZ1tzC3WgpUx/RWV6Ft9N3xHaZ4OKftoOF5xE+6wPkwWjKxNXMaCu
4eB36zROTHx+Gc6E0m4j5Y0R0t/bnjB3+mw4jUT0wuj/UgQO4u9sgiLycx0SbtT6RWqGvMuExjh4
xEzdKZabxIJ5O8aYV/X0A4WTQ7WHIOqYcginoGYimWCsgSRor8OGakueggxnT6kxz6oSywZ5Dk/g
Sa4NeUTJdew1x9ilA7PqKTD+J1QKA1O/bZhsvTxO07kHyh9wDpKDnfpgcAlWJftNyuEjiXgdJF/S
wTGEONkjyuIAMEiGKbRkLyE0mCp/RgMDxt5PNfkzBAbs1JgQylhwDez0/6CKjfhKOzTTsMUuX8hJ
n4SFbzozylxvi9LXEmnOaEWKVHy/UtRxMgMC58xlsM5eXrhcY8GIrwwFe3ODIe3T3zm/YEmHk+nQ
FlD8LgVjuc4IFSlYwaN4odWUfifq23NxB7Oa2LqNp+F7eSQw8854fhZxdFSBzWZxRpVXeROfZYaB
ogOGlhmjBKnxT2ZzbIqViQ1LilWJSx/32E3GgqYNfQQw8t9YKBd9562DSMHI9LUQKIn2A1w7ZS6h
6LKSzqUPEC1JemfDP2pmKOlzV5mPnFhcol4+Au9Clg2hIuXUNmLmXGwhrIy5+1WY/+quhIUr7EjX
WDkK+/pHeT+ENbVmcOSPIEOOMAan3Om3pRZ0KAj9bAVXXRbmrqvLIHymcbZMH1wz7cTWFqMYyFHm
gamuu0mInQc0gD+EfPmxklfOVdEJJ8F0qvrmS+sR49ihExN9Johbs9oFpUwhZ/2+K2fgfk+KSEuP
ZZaBEUWxUUmssjmbUw9rRpJKiim2VgwjWHNUkOnVfnDIxeYOohoWQ4mn81KILCHd/ZYDTfefuAWB
mlb4LscUDLh97p7Cnww/DYY7YpM2VFoK8vsfRWHojahJKcbBoCicUDuGD5H3fbr8nGgwZXObtL6x
0gJSAItuLtVLBeScTr4i91J7B0XF1H4eFgo7LFH9a6DKYg7KRe+yYyys8xTY3uKVrn+6xkcBy4Gy
T2g4aZ0k2d6DL22G/qk+yXGuaY1t2YRTFDeVcHVWIJ3ALk9Lb+ArVsUUJ7zBJGKjlNyixyL5SkBa
wjmwsEdENFMe4GYeR/T2PP4dnqxg6wcibj3UWf4XxTcHJuEg9AffLkOiHV4L+a0K2eQxdRU+fLlv
9NBgfEbQC3guUxapaoK7MIbegWYHQRcwPogOuundr58TuCvXn1Mazo4icBHevBEuxOaqtAR2QVfz
IyYZHJ2D960VMFJ/z7D+sBo3WPts/jbsel9ZIqyvdYcRuLf/54iWpJk+0XU/2LgF7m97eIsEG+tM
RQx4A/zVLZ/XdpSp2/PQddEv23t0Gk9xFK8V1ImJOcvzQHDR78oTZxh6IAumXw2+DDFzbp8RgYGz
Fxu6Han54qhUDP39BpCZZoiULLgdVv4RCK9NEvesxNRewwgawx2RihmCJHpsB+yIFwEduCF/qdjh
k2N5BuoVQEaRbx1ACdMf2DIT6G7e6jqQWhv/P6pZwn6EIpTjrF/+B94U8CKY11KelRpxGAh9h8yn
7UMYbFcBoJ/0Kz2Rly+vlloMdUWMDJx3EC/DHefSZTdoZQSRX081xLr0FuXO1SBG+k90hf0CHIpW
o6lsQDG+LQ+eTelHBRbceMME6hYyO42nK1LNS0DIqqFO1uQ8hQ1fAO1RZK02u43mdHEAt4761M7f
EfEcVMDdkoagElCYlGxKptZFgi5Dv63Wt4BlrU4EmDa+WdM9bv/+uaM/M5d30nbVRaVV3AeU2Vtr
JvUREY0Leq2zG7MW66YpOT/BsoaqX6X9rnKlH/yWkXL5NnhMw7wnHM1nI4HLqgBF8RrlR3NkE7gt
dbffW1TyVyg+SqIHCPBNxqFokTpnUrN/2QDYZkZSaQXfLI0S4uGUjLWQlqylIm0sK0Q6FMsd3pyu
/iAzCQUWuv1EH9GjIrlCQ2D6Kma8A33gGcvYr5WRC46lZK7oiweje8DI0Mgs2vqh2UE7Hq7CgewY
NORgKZ2gmpvKqCZK8xtz/Sh5vt5P/zLcIkoaZeYxie242tDPAYhVWz/7/gnK81kJGxRoB9Apn7O+
25mhafs/Is+NyhwziDb2GXI6oreZk2ho8HVfpM/Tv8h8SgGns3lSog8zf7GhZoEpbFeTsNQpELdH
W2SApS75nTgW9YKFvckJySQZiIOa4fRhZUuLtN8XzASfzX6vhb3abtFG+GJUzs2bQNR80jB748yr
aFvOYEb26wKN6RQboMbJgXSCbXDEAD3Ij022sSZGV6epnENtnJroTcOtKoIRE+k7NIlZqTLA4W+/
j0jJHLDJkH5uaCItpDsxpaPbWL5RGtdAqX+kHHFiEaoG5GGdOaP3yUraA8ae+w/+oOqCcH0ya0DD
8IXi3y0HkkOCcUb2Y05NMHQv1kJg34KG3iZjr1FvlaX8INGumfc4OsNDPd0yHZfm19o3a7FiX9lv
XMIN1egdCFy0Nl+GgrmhI01sDj6iAbbtwbA/csT4/VdaTm77lY8U09lnuqyxk7HSHjxwusXjwkEv
Cg4rKULxJcmpexWU2CENR/TjXsN781Hw5VrjLcj4LvKl1QdD0zikhx5kKNa9KOy16t9b1RG/BVa0
W5vY+4uJ8qFRY5UbDIqToYYFiLYlp/sTsEwj5QjrM4lA3nNMBabS6KLmdBA4qE65apFzKnZ7UgbD
aVAnudAZ9t4RswYuklmGoEqaEXyezrF9VQJMDXmcU0T6RIgmYYY7CTc72Ku2WFsUmioqzSze0te1
RqeMYbxjMALoGatZrfjAxVuUKKk2nln4suVl/sIEIvCjRzzLvDfQ9pCqTEEZIKe/67ubezWm3e/K
19GOwDoBPF7IeY9EmXKzQ1beVNiQPGBU991kqOzKblZKOKltTHF4+7BSvT2eAA1cPeysIctj2Yxd
l7U6K8pdf3rJBWV0VC0HT14nJR2BUw/Zl1narwupno46Qy2efdtZnzRDJDOWRWDYVmNB7/yGhHT3
mTmlq63xlnHaiwGL6Zq8dMq0n7vY8g3h5x5znGubBQIzNRMSNfrAKzyykbf4ClaObOSxlfjd5xrF
wtxE64iq4CevEcd/mKq14pD3ld7tngYOUz4AEzu/YJ+Ej43gQarfwwF6b0AveV+zdclHBSP8X6qp
Azkw5CJ7br7p2IutTKZasllkzujyHnD7LnbgyNdbzev9ChNWmzv5Ow8DCK4rD2QkIW0nxr/E0r+X
hqWhVXchnxgW6UP4jvryYmkerObNjP0RDYfSBDbtE8bgIqs3ccHNRaqOisXcFuKEqL2u5Wx3tfVK
yU0pL1YgZnDJkU7QIDzSKRGtGQlEHar1LGJft1D5LeYnkhgR2RGDqqZdL4R6NR98KRQs5nNgg1D7
wGnfoXKQujiSIBznU+ThJIla+kvamIcXQoJCssGGBrLMpm3gxj0PjlyEkLHCFz2HfWiDUe3TTa2X
6b+0MvEuAMbXgACkJlxyFt6FO9CrYOKQvSI/WtVdlfONwS7cNKog7CgmwNScJAeJtMZRuGHUZ8Ra
3Lje3EsHtQjb5IxyrpaPAmABjn/MKG5C90qqTJmRVCmkhXr+uaVfTwjZSgSbpEM4ZufoxRnSDFd0
dz8ilpeiQn0zI5SepeGFH73AoyHo8ghm1z/Yc+LNtieUJj8WnVIVlmqyFvIZQY62G3W4INt4AIo7
N52MHoeF4a43GDBK3rJLAygBCCCIqAeaNlHGtz4nYTiZ4qJ9VNebyGJZiMw6RJsakVowjb57eNYU
x94S5I31bAh58X/8CouTOM/wlRPEwPEEs5IR92eDoMU1XqOyo3I+JBilmd8GDewURXpiuPBxmANJ
SDIlUlg8yUw6DiY+id8DHL4JHN23V8c1pG1BtHEdZwjKGNX66QfYJm8eDrW2RZS+08a1gFGV/PXy
VvakXSWS1U0mzLMfHD/uE7GvsGzUrK/tf+Svk64YHL16R3Lgpza65VlRYjnAQI/Dt1mSI5pjMtG4
6DU9ThVFO9JDjJnzPMm+3BFVkxjKGWBY4jKoPkzplgjiNY6W39YZfakVAFm+v0lM1JOdsSDve7/o
AAImlrteV65Ag5KqjK4o/ogEuoAA/wG4Wjld5L3IUCEMCothWJTy9b2PYWeNqbD9lwKeMKTUIEa+
yp0Z4h2R+ZqWviNR01mTWpS4PfQd1u1jH7qicIDCWkvi8DLl4eQrKFYJMRGSAuvJmVJxOUmdQmyV
cwbIi0XNo1a1CHX6Kj8omQEYY6tfMMEmJ7YlZ+nEevWARCJ4+5f2mvF2OVG+Iheu3SWW62ymjsXm
XwvFPCNlbpL2UNTy7gpClyeBuFhLvn44ZXletYnWUaVd7VGHFruzDtaGZt/WjjuVZUVm8Z3CCg/4
eumS2ln9jcAowKlRo0vV7ExYHnN/20FUKszQHrnEL9rFuh9jyToBJYwomeXWoqkkPuYnPV92ppgi
mTcTw41ipkyzPvslLNRSZ3mscxCko8H0DlOCv3AO3a+MEh7uzD2jJmU9jDx14sqMK52Sz67Z8uyE
ShqK0TtzhNxpptJxheIiZXm7BYMb9OrU+cGlQQUoivoGPQhuue2rZWuNYrYcDSh1rpZclsNcSdHc
sIaEVFubKYSQPnn5oUAfZrreFXhb2fQ6ezc2epoQquVv2h06umH9TsFV5kJr6zv+wc8yiPqj6L1Y
IfPoxv5XFuU8eWuL5DKbb6oGFzU28FIhvSETV/HbEimndZM7LN07dMXQP8jOlPefgyeyDtmlo9ln
U0wL+FXw+WFBVUmtc2hyW47t5bOPTuJK3ghYPnW+2H0KHPmL1XRfyIhTE4SH6ZnrjBV9+z7T3RD2
Y6y9eH0BBvcBmQhHVxWcz2joKp2cPqjTxqa366OOTbiQSGJE29x/xYBvA9e7F1ocxfAN1yya+gc5
KMbGSOUYLhhH4VLutjaToDomNMMD6041KrmeyH2VFOgKmB3nkxLnS8Dh8BQ4y+JqIpZYbEbTIUIP
f8U6GomPcc9nlOfSHapryRsFRu1m0ylsW57Qb+N0Ku3byzX2bgUYo/+dCexeLh8n4mDIFV1ISWi2
vu5JBXacIU4DOuykrUK9jV3BpWl89tjkX2PbSXr6QypQUApqR4IV9yjtdcJRgGL/eqVG/VbPLcVp
OpR6MiXPZjTFYFcgq7VAgZiXMFVQKnRAhZB2pse48Uc7tpVjh/llUpG6wt2oS9ah4xPm82Bsw4Zr
rS8PKf0tXM7MhupjpJ7B2vOoVku7FUR80skRGawmLYFUeP2CHjR625usPIns3cHGIt7iHjufCSMR
/T6PQ1NvEH8AeI5WbGQJUvZkisdUnH+1r4nyZWGEgHSRXEtNIwKMz2ie97WUEJrPErg10iuBa+IU
XkY+bPnhDoqBvlI3ygpz9k1cs1UUBhSAj/EpWO548YlKqDWip+Ct6JUxtO69To4OT4r/cfDq2C1S
vI/gy5M9jvPFQ/iKDz5MenCmIi60yVHmd1VcZpE20Xt/iRez/aoSWlMfVWfAw3DHXvwJFbicqftN
Qx+lUmpSZQBUHax1thfQbAOXSn6MguhN6epBsXrSu34nHNMQierH1Lwmxp1HgE2LCRw2LTS44kod
FUJLW+CiA4Juy2HEGG0epKwlLT2gmB4jLGtH0upgR013z1KN/C88ww+/EMx8WYyIrMpu7Y978jF4
sQblXXcwIGm74IP1c48A7YgoJP6hka8NQRt/AqmCOXC6yk9mxrK1PgWctuvMPFCwGeYUmGSwmALP
F2g/QfrSFbIgD7WWL2cZWf5QhuDbQn7pqncG1QWXc3SQYe5tEBk7HxpQFXPrpfC+S7hYspmJFfnW
/T3oo5oPDzOsHs+EQLwaewCEXyBDHA/HT6HMMBVt1NM9rWlfB/ExbAlmcjnWbHJuOwbCLLmMriaw
80z/AK0ucROyuWR6xFh4wmdPscHmlc58H79TDhAG63SQf9sUcsuaTGVSO0cuXPJPZvwY5vzZHG5e
283d01IoXSZkUGlHHDnOSKAubn9Ufnsvb5nDJlkTusgJrVnLlPAagMphpE/cjNslpdNLn/zUMr1Y
/9P1WsCK/5AJdyhmZj5nJ4+7Ns8TkP+Wa70gdvDmA7M6ddeBtIv9Rx2rRafexq0G4QVQ/180IB9w
jdIkj8jadUo7HyqWzcnjrXjnis1LxlW2hC0AA6XD54WL89MuALeGx888qVa1q3IRy8hjHF53YB6+
g0vutSXN7hEq8AqNRKKx0HhvKLe6KsqzZ02NpAjzNKtJeJop0SKASZpUaDCiZct8gyrmLmHNFvkX
/h7nv76FHhJ4OSB2MR0Ps+3qutyQZkhPSCB8ESerxfLueo5Cxm/fLavSgOBLz1HA33ihD3KSiLO7
viELOHNSPmjirQJLwmubnJTCZ4On3t/O5VtYUo8xzGJFn5VA2sTMWCxyBB8VTfw/yDqWNQdFWHzQ
q+38KpySgiCkruK2FZV5cD+dmkL4G4I+Gmgc8v8chhfTITMitFkSYcIXuFVAvLdX10wQ2YpKlsqU
RCUOvwlGM4p6od4xV6qtWpnhD0aR2nGc6i3Y9DTwVHWv8fsQ/OCuha3JNTNnloun4MgB2TDm9WJ1
+KDYM/kg+9smMPheHKlvavflAAC3WCgpntsnpqQ2/56lxl3DMGaP/xJdroCN4cybhcfOAtzO7OIi
ZmAs6eC9O+hu9eDzUB0euSsQlxhUMMOrhGXmC7EQnKzOdAK3vz2sIzBjIM5STJ0Za0gtnc4fJnuk
nDXpojrjjzKvNtrN7Mi7pmcGs0V69jDcfAAT5gc6JKqFcn3RY4oRDO6CUqncLwf28D9x7vks1krB
alzzLPY36A5tDdKQv1FdkQhcU75E0yNDuZBO5DhaIfGm5hpS6BlOYJjz2fp8GsAZEhDKRS9I3k4G
OlURvCdNPV91yOBWBW7k2zSwMuz7xT8Ctr58husm+piL+ijUfNj+Oqzb8giPfJConvypIkadeQDX
2BloB61k8jgCL9HiVfZtf7HPKm1rpEc0zWll7ijxyvhTTsjJcQgJTsrmcWd/wsZdc4htcfHtgjzq
Pn7iZjghedjl1/9HOO+fcuaCeRl64RQ3Hlw9yCTu7/JQsMyiy28cJ5jY6uOH3o1VHE8LaEK59bkQ
u13VManTCAG9aaYfWj4RF6jRHKm2RmKUkRkL8pDGmKPZEmgHheCnF+yxg3weF/mTMDTu9RdspZbF
Ep8p17pOlHZOeCm8JpGjffbsrFaOJVWX/7cZWuuLY7ap4iPF26lV6Fe9yMxtH65BFHlQPO07BqP6
H9DbhGs3jXx9HJlaHZcdqS5u8vpfO2aQrZUiEhOQ+1+usobWRR8MIYBGURk0STPGl/1AikCEHF18
W3ZwTJpSurvjAzNmM5ehhn9mZHsd1iCoj8+6KPsbI9xxW5rUjllZCoGjYSLUNb8BB8/1Pt7HVNOI
7Isio4Vc1g/5KNZATUGNteRMZmg5IoPkzGRKoPRSUls+u+e/gm4/ef2TKMx4g6tIx17x8A7gqz6q
lo42F4hikxsngnbivVwC+pef69HbzwlnCBimyvK1fOet4zBiyi1jQMZ3mEi1teG3RC5G4UpHV3Pv
iNHKrXO7tNnry8FwiDOcxCZkVuBX+e4PUBt5uiotSC20uhJcXhZrA7gzQrdc3tBVehbgjizWEjag
tyvym7NMN8T5KKIvasMzrFOzDvg76Yazz6TbbDeq6V55uNHCuf/WZw7qHb43gqgTZ90PZUHmcTSd
8UFDkeMrp0d7Vv++ydM+YtHu6ub/ytC2L6Dn6hGBSC+D6+qCVLfCb4G1JmCzguZktFtAiZbiXXuk
eIODP7AQC3CWIkZDC8mXHSUGjCwVoWf/V0YgjO0Aj+gP5MgYo7/ihWMf7B4DGom2NrtW5wps+CKy
NpMR1p4OWDO7I2JmqEldQWLDlQ0kVsSC0bMkOHV3hoUgOLoN55ak1ow1dHUJhSZ/8UZ3pSNzSlkG
0P5JOlVxsoK9nMTXs9KbxmFRfpWPDKT5A5jwn8Rz0KBpSyBsbxIXo44XhqyYERm3MeUcvE7VwZP/
O2/3rCyyVsVShR3C0e39BI65raYFtAkHe8ttJGlx3PEn13D1eRpGI8zQVBhkTSgyRfyG/xgPfwj4
kwXeQqIBFRblqggiasb1CjuEyRIQA/64Wetw1ttf2BrBhd3ZmbiE8QwMdExIZZtiyMI0+xL5Ca5V
7fic2cAOhaUnbod+2NLmYxS7XzW6suVrtCHypY/CoGnxHmsR40d63nQJwS7qJAUJlv2zE76y7x3Z
FMVV2kDapUiJa1rHEDPQBeHH0uFMYYgm7j8p/l+IZqiG1rplOawBRjBhCMLZuh7Tq1ZEAVJT8e+s
RSvfz4I1C0xD/JXcsPrJv8+JKllXWKjEGOQ05/1JD/t2nXz9Sv0x4KW40Y3SAV5duEAU3LLP3m9X
stxbFPqvx3XzKigvn550bN10nENuVH/ISywPwQOvfUZaCntaL7+4G8Bf1KiYlJrS6CKA3/RkSm9N
bRFZeq7hCFLZFSeRYOO1MaE8Ory4oGhkKa3GuwjL3okR+D37hIszRk5PAE5OV/aG77AYmzLH1I/Z
hjOuhzzKqh9aQXgju6hvHTR0ZNxioKX+QMdlgD41enX7yDAgu03P3uxG996oSWkA0GeYuiebHbZZ
56QtAtJTsKt2NABREfuRMmezLpYK/rMextdM9sZy2MnEsEwOBf6OrvdcYsSCOuNJKjRzIBTdvdiy
6UyXHAF2Gm7oCUwRek00YhuBY6nFNmsoo7WAbsXiGnpNn+fRTyynEh6IKh/JlBKk5aHcjoHfZMqg
2gkcQMd3DaPaBB2flddsbGqoqw0u0Rzdzsqhf5RC3HeZO2vL83nyu/zkbuT3oYfpyn26ZDeWsoio
sUOhQ9ak/jDSzUd1EZZ5e7WT2fhf56BhEX7+3AEI6AexttdsP45oknJtdD40T+tC9CpuMef9djKZ
R/xNDG97miEgOQ0bU/TtnsAs6d00iFI6Q5KdF9TdVZVoMH8t7U2xstvPqhOzVDHXPDcH4Jwcljm1
RRAYr7HHlTub+KyuNiAO1c81b+pCMNeBZfK7JnYSr2LHgNfR9CjHISB4ZLX6l4t8gMvIXNIsINYM
pcB9yEyZ5RU7Gw9QYxphktzSwOZb5cw8U/NaH1H+RJWkWURm/kKbBI6R8sd+b2LWmfiITsAo2YVK
OXnCXmMM2NbE+cJQ4Uslby0QfLqg5kvc7MuUFb38xbcuCMjoMTdS2c0+A6F2qhFF0kW2TuZJXko8
6pwrESNSF3qMD0ISL9m+Q6i0bugJjf9AdO4r7iEkvenOPwPodrG70ualZLGE25KnzYoZ3pF7Ans9
Ntg4y6UCHTwjzjM/UHG2T1DfQJbeIDFe0AkeePP5kDBJ4KlihUGnHnsL7CGN+yyH/Tn7kjrf4h7Y
uk+rjhF4KR4OIcTM65oByBpnE6oOmBPCZG0JOgv0g/PN/tkQ6MLJyVKdCWnItL1rYrjBYmP8mapd
im93jQz0LQSpKHUmM8Z2MDAaoOn00d8RcU3is5OY3J/hcJRkQqF4Ly6bVxnyWdcDauSsiZEmYe7i
G9LabNKU7UnMSVnYQJjKMIWCz922UhVKi1oAlq3NqCfkK2wdBg2SW+ckDMCaGeKxbP+/gxUDmN9Y
m4dUBqgXu//69f7teKgJvxqTiGuhV+xgEsueYs0mR4NGuH6T03FjwZnR9aSySqR08Hbfau70FGq7
4ALj1WRIxzyL9DbGnD+HF0iMdmXSbIXBZ6/FVCgTA2r24iLRLta+bV5J4YG2jkIa3aLbKu9kes6u
KtNhZ2inUdgmkRbbepw5y7ZSIgiP+46/fzApkEpIOmRdeBzO1ijbkJyHdCOl4+sokjZQkvUPh4l3
/EHyNIPy1pAqagdguR6Sjfj38egzzN4r1Co4rn9bRtbpqw4etLa9UUYF3TqWT3CEH2kmMIWGIq6d
1z1S2jkSJNTzHm6bDPEdeRsS7eE2Vjl+62Pkdi8cavcuCUmjFRXCHtI5OzCvCLFpHSlS8UBt4c11
tz4PMwZur9Ee+QmRmY7dNCcdV+6OAeavcYD1SGtQHYsm+TThYDya1hEwcu3RZ5k3pdCfhUfGwj+K
ujH0JU5OtkJgGcnSixE2zCB08UmTg1irZJjjM3TYQx3+ghT67vkcsMpJAOPlTWFL4Y2pLILCtKbi
liu6jXoXGfIhmt4dVJ4J8FnnqrcfK3ZqwxFe8Gkpm3yYzMLo3TCCV77Nc8F3REH8szsirZdqiR0z
FAgcBc79AUcs90w6+Nz3NApCh5tsH7hLY0GpE3j2fZd3cm6vCdiCtwq4WZuhwJITT0u5i8MzOVv4
zgT11W+jv1euXilRuXHxV9zfLGYHD8LiDpQFZyzEq0R13BXLaYi88tO7lJl+RL8mXS+K+BQHe6xr
eD8J74qPsqqNxAsEZv5jcXM0gy7uzJorUiczBoRaHYOSnrQ98pNyhcfoyqa8mJ/f8cv3ORN2ZIvH
UEUKAsA51My1Ntl2X/BV1qBhpwl+E2XRWbMYy7Sfg8qgSqWvuI7XL5n8BFl2Yu1AFgdMUPMGXXqI
p4NydOv52FG1Pw1Xip/C9owpoPtsqyAjamhNWXV+c+whXadM3zpSAmLf/HrAVGD1ON2Qv2HAffVJ
O7eIKnEWz/TUgcl/px8GOIoyUiAZosP1wyh7ntR2t48vhY0MmvafOG+6FooaXccmilmvcb/lYAFc
65aFFPtd6WnavtAubK68eLrfAXbyYtu7bDeCsMsyOoKbv6ailh+QXI9L/zaum4RmlXYW2gjrTmmp
bo9T+7zFJ0DOh0hgEkZyvyLJ4/0uC5AA+E3V4Awan9tsLKg8L6fhRcoQSla7nv7L03JFyHqYwQm+
h848IEwS+2/5hYuI6S+JmjmCnpvbfSxtnQnwLfZ/kdclk8LalZsmZaRlA/bjeQxpFP290vHmDG4v
ef7K4ZKwJTja3PGTsNuXZokPll3M23Pe2TZfh6wBQzjrMJu/sG3ExBiKIdPpXbBfrvbLcJetU4lB
ogO8gADpJZ4dcqsyu5g2mIg1u8xbdIU9keGHr15YbMf+u9qGCkgFrgDaHyFxX1sXMDx/OraLqpZ8
IJIkXXkpY6kmFDIv629dsiHp+r7cvxjMOZ+2lEKYyw98yK3DeWW7iTPqShTgEkMNCnAAmUKwstXv
f8Evtj2QZ0fBu2l768GfBJqLAPlHLtzRwBd2A3PTur0lsJQ04lv8S2MuE9mTZxFamrQ3zjQou9Ky
nAYGp1POH+lBv+NkyeooXbJ9ELBE5LHLiWHlct83lC1FORPUftShHJsZ00mYbLYlRz8dzuJysROB
eVvwtjmebbu4SSlrnmkB37XndXOe0Fn4CDLgrAUDUuGEhtyLtr0sUuMfCu4ZO8rMDhJ4S9z1O3Wf
apuYfjDI97aYccqSLZZKJ6Y49NIrX2rqNMTr5bJFjLVLp9yIegCAU9nya2oaYanhobrwfV5ut7hK
t1mz+v8mA01O4lj1aJRM4UC1WwwSasbTWtedJt5v9yxE8v/PO0YaHpD+ir0/nx+sWlo18SF2VFyE
Y6Nfhw4/ZxatPjeSi4p2xFPgGIssfSMVwr5CmFKQS0xMO+zsXXJMT8h+8rpVHkXq6zChhb46Sz11
7sQW0fUwdKIUfh61t+APU0oKRb1i54UzQ3R5X9Nxcln4DUNYsxHH6W3MVgYq0qn8PRTwICh9A6sl
4Z3YkddueYnHsp1Rdxfq2+r/5ZrsaSY8RNmpq0gaar/JA6HrO4WtwXOMarbMlqXmuFQrmnhkkkNr
3SxCauKkt3Gjeywec2gZZuAGi5olnlsoV8ag/v45F1TGRDq0zGOl90z8n4LbWbd2AulHapDS6/Be
gwJYvWLyS/pqD02KtgBFo151k2pygIMDQAYvVizOwn4MYtscRbrIiXUN+GwGT5DW9ku4hrWCU5a+
q3RPzluTQvCWajyY+RAGgI8By0p9jn5sM+DX/M+jJSwq7aQISM4sann5WxrDBXSaJOay8otLNluP
puwDWdqgup8mbC4ZgDWbHnma7rfC27cctjLrU7aoJ3fL6+rR3Ug3qgc+5vEb4RL/Y3XqeZAmWwbH
L3FxKqIBpqkvsP3ixMgg4e/8TZE3bY3pZa03AI1eIEoqhPVkf12vBcsiKCh4QWGeRWHwtReZzyp9
6ldIiTSbf+UoSDYDHU7fH97G2jrjRyOmJeZujRkyP0aTpgEE7CMadaVbz9OA4tSwwS6g2bL3G1B2
YJKKif0IMT5PeaxkrXGjS1P8jooDYcs3lstTdH/r4Am1bGOPu5xAcdETDA3+QM56DRH5lPlO/TjE
4hbba2KS4DzfRuCXKhtOByggrRKU4kzEtbq2fidmninXFzkA4UPseCPeefg5tLrPAXz9YxH9iMTr
TnmC8nyBhLdH3h48QC1nyjpkx8YE17A2hweeG0pJUijU/gRaUoBHFY4V1HLL5D+61wEahS6MexpR
txYROEYScnGf5HUwoIoSuyWIzh3hlGBvWGLeDNhFFsRU/ywFjP3A6BhIPpk+GKbcQ5lySeLMbg/p
T2hmak8wEGGFd2W+ECUaGSV9LcJ1FEKEQKwUWnRZdvbds376ib3q7KuyZxCKjgB22gr3HD/mlavK
MsCkjnrjPlD1nxNrl2mWL0FZzDbNBrPA408ZuArUknEQzwb0L9XMEVhKX8x1+8Xlk00RPioPgE/L
2xQtG+Wje7Y7EAFFswBzhnfGWE80yuqtXCBEBSTjLpsMcURnlDoI5wqtAmV5LEK/M3VikcVVn1Eu
dlJ4WbO1OBwZo/2JzMAQNimKQSKQJFqOQc2Gl6isZ0oNitQgxAPpbmPWTQtAGtSgB/5eCwq3L2w1
0Cvaa1OQfun6X/CIGapkndd2tU0ZbBVhHaE1JDVeoVL/0NZ0s25kbZcfqEYFm08VBxvxpSmIXHuE
b9JpzJAVE9b1UtqkL4v7u6ofNc0HERizpcecs4xqNiifgPQyH+9/VnZcoMD1O5sHFv93Ek1nouXj
hLdIo9u5TzGzbThKz/quGuUeRumzb02FngJn/ijtGyIZa5G909ZnQ8r1XXrWH5Y6CWW0UEYyIfSJ
2rDsLtYNZuJI+ABs5DMVUZRguRWd0Ja3OqgNoKkQaH4XKO7gSEj+g8vXwOQs+rNI8LsJOhBXQn1g
l2V4o+dGzsPpfB+0+5lSGi/6f2VDD6OLKxqwh6nTtydaNawtOwWJvS10OLU+AqeRA0BXMvxsExap
t09bbH+nHBMHYPMhvMcsMrr1ZP592NGjTF2VFhUraL6YO/ooT673U/MLpKufZqhac8sRmK+ScdDE
7EmfG/SwM+DHlGejJiEOOeH+CRX2UeyaQxKX+An+y/c1f8W6YKErVwb4t65ohg2Chrt9tXI4cGTT
0k5rMTrEcs8NOFQ1TWw/XrvbX0qyV+VIr700vdmrcwdcWUG2V3+ppaphUjNfC1HOaCzP4p4GdlaX
iWL9ofWKg+ddxW1RrQj8eGxHf0PixvIC98NjlhWHlDwQUNtsmkVyMSKYVuS2PAg0cOwoOeO7Wrxr
3fjzMFvFEYp7KXZ1BFX0BYrFknNxL/wBGAz0saFfjC7COA+lfLjKCiWjh1UEq6kUMak46SxFHRtx
K6yYY+5T8c6/Q2+kFipG34JKKkREPCagplvkFec13SpBYddrfwM+Zo2eib8qEJXXqvgAHSpp8+/c
4rS9R9RWYdaO6S1iNvcEGLxp2umRMNMsQR7vytaS0sJ1xfz2NTdLzc1HTCSgiZ+gnJnaGfTHQvYk
URon7Fk+STNyCGTOYCWzZWxMY7PUxlTKhb/ez132G95QvKgQZgLMkoU+SbELE/G05xoSQGGowwtv
oGnvOKRvzu4xlkwpP79kqiQuYyH4P2Q03CvLk9CzD715HZh/WgN1MY+oStmjS9VJENzlaCjQVdb1
sQM1hxDlI+/5g/ZqjDqyfYK5t7JpIZBdaqVFK2mmIkTXRX3MP4OGYQ3cfDs2mQp6rheHs2Dm5Dv7
FErkSAg6Uon2BNHbTELFtE+RobNFGiy6yI4hIoXqxpmxGJ14+sVcIV7RzRgs0kDvEZKF6Dwc1TXK
EbtWlHxa7XpLOxk8+gp17wBonc+G+rrxKoJa2wsl8K5VFn7uITr8IF7L2XhT9/OTnmdImuwbV7Nc
e0LDn+PVWC43XsyOc2kkgBtO5mug2wFL2/FgTKoPcrxRBduos0f2T9z6u1ka5RTHvfvJZy3SYmIl
mJVhDCPu1O2utTWqZ046WwEnGZDeEzNE9AWJg5HsrnSeigu4nfzhih2SdEDaMHWm1iLs0g4WS3Ym
zWFcVTFnvmMbjGdBY5xfkyn7mWxHBMzuC6ZhXeY6fpZJA3JA3YA8BSFVFnpw/FKrIqtjKaKovV8Z
G4RA4yumfdU8QwHN6FJyUdtjxY9+SnX3vyMlc1EfwChxWWp0X7cOzTSbP1MdLY/jadKXZdgWXPea
yCX8Iq6E4idxd5I2tSjjJN459rddspG+5CSgOhSM8fxhjGRV1POXudt3EuEXXEQjaBoBytrVZDF9
rQroKdpjqPjtISg+A5RRW2dp/C7wV/CAnPyw/gYRFj7qJebPp5SGdRZpzi2sImXVzLGJYVY0SZ2b
1Ld9OABFquDpdQwHsGBuoQ/JII27S2nI0htQa7aTOLskwcyNhqtCGOtHdSZxzV85ySueCXwXM4ja
OvZ5VANgER6EMo9axKgQT04sIwykUP4cI9uGWDnxyU1J1Z221uz/Iy0EZfonLbV4PIWmQ/jHeVWY
Ctaue6pK6gmFVBsV0Zp6SNs9euvrjYe13bNkDmILPB7opiCab7a1HhssRRcn9kolnCcH1m9hTzOA
/CtG/+ISYlRFJq6PDxBswR4B7wMtGOLKK/sqPM6QP3zjSV0HSvfN84apDbh+X3VLJPZtofUw5ldu
4I95Vw4vDeL9GrcKkooJViokBD2mJ8LHHE0sH0K6hwrquKQCuH+OFIcSspqxkAbNW0HOkdh6Y16y
OyKrUJ/W6YjlfMhioorCLM1dk0ZznQHBuFIle0lDJVuADeELULRPlcDx3N9iJvtcuVF3Ze4NJAQk
37eHRp1ypD6X5n4rK028qTqebUxvkCjFnGBUrFBoN9HjWyRC+3tIVhc3o0aGKF+fxWmcCRexRqYw
Q7PCy7PWhjLJLXaGZyboFH+BxcDXaeQQ5VNp6Ju25hgdEpQwcZAwPSj9FVFrucC/R5LsecHdCA88
E7ZM9k3lFrXWihL8bmvsKx1Bwtb2SrC1wBfaskTIwATwn45nZrmw+BTUDT5rHuDfd3IvYoWvIIaW
BEKVayYpV03COAWpVk8JevtVyZH62eeY9MxbsAEnOWcmMinBZRqaJm1n2tqMABLPnQPb5AHVuhN0
ZNkUHMwZ6m5+20TxT6h76qJY/8JYFlVIMMvRMYoZBcL6RXfsuYgIbXoiwqj2iyGpq4FfGcJPxpmh
o5/7orBuOD+SWUI2roWRvflIj7SuZZk3kPVV+EBijm+ssNl9jW344msAZ+ZQfpPeyJYzZ76LT3sv
YLSfUCbtOFmnPpigUNSv71GP+IOF/Ci44/2MhuZNMaOfHUgmUoV/5Hqv8NfSJ6k7nPg5uQhLt3pl
4Rg59fA5mx4B0/T2nPAah9PTUg+MxVigBNTPgCV7dQZNHqtq7jL/EeySJ9cZv4MTvbjhRMS8Ft2e
6VbArHsFyhFTUeydR0dHoEGypOm6enlyNlwTVn8HZHj4S66MIMJ1vKfunMrvIBOhL+xooEVIZkV2
hDZefI1tvAFUo51nFisny5O8yOx85rdHpzpDFabMx3eBqGTioFy/pAb8nVlqIQauCR/M8xmhPmDR
5Fpl3AgHrro8vhUjBlDLcpCBe9qh990RIpFut3+sDrhHti7fE4SPRo+xkcLgXVyLFA8MbEmxXaRi
pH2D6E+Bwx4Rr4D23PQjMGcQsUlonvWPxsYB3ve34L+JA86kY15juge236Pun8R8NuDQknB9lGhH
HpG+W0o9pCW93yvyxu44J1F9pw/U/pl/4BSQBcqd7rYbyko08Q7yROtXwofVBUJhzcd9h9Mx8bcA
14SLQbuuZjdohjcKRWJGIcGlZxCKagtEJNS9M6oNvF4xOCvW1kllZA2PStDLgNI9h3s/R93Icl5N
d0g75MBeHTZVjCRBeWbxy8aIbabmIgWWzqjRSXRO1KQMDiSavgIDrKEF9kPoRBcRMJHmm6+v+6/d
ZHt2WEW3rTYBaULel2lxtv3WbQo1qHOMHQnIqYZKXaLmwnByYWKdgeGtpAB2oWaCQeOV0hyvvY1T
N+ywg5+DBZEHJmthB1Kqx1nBaOxS1tm5O/GJh/sxXTN+A5YCuPzozXAfn4Q47ED4wgmV5aKwkuk2
LN3/sbmc30Ap4O5DSZR36+SIudqQFlyvjGxuMqB8djPB1xLBSsaodF1Ez0rkFFMtzftKDkN32C7B
R73HCj2r4plQfmZRpWynhCK+dpkUz775SHsVod3LlIgR7mgBqsSeiqDl7S1dJFkIYImmSZWcq/+a
7gOItqRcf3g0BIHd5zUIdfBzNMSRz52MJ+NaBoacSNbCQT8sxQCoqxFfhqs9b7vqPJDEHZjXX0wo
PcpIBz99MTCd/5aN+1k2+zVcy2gomghdHD02ptQqF+3RAzmEkkdSaQHNP1ZAyCvEGLZ0urn7EIHw
5puGGBcueeqpsfGwMHBwF/WRyrfrqnJRmzSvyGoz8R0xm4EKZI0cTVZvb4ikFiqDS6Y/h2gTJPmf
DpGPji6ZxyxpWO6L0JwKDOCepD5/AZn7U3UqKoJNwxMKoMxAlKYchYEJ349imZIqHqLnXqRokDmc
6oivTKyo21Nm3sRhorwpdjru97nukGz+qceSkIm0LRT8hroZFgNCnvTRg91/aZW3CXWXP18574rw
Y17c0PbTQqy6TdovRTjSTV9aKHca5e0HVJ4Idh1OKAt5cWPa5b9kXmcj/qq4T+RkZWGeFyC3hDAS
IljYPBSC96P4f+56laQVLPtlCXQBoy1lQXullxXoYxlxCz/ncK8+nhAN2h2VcXUUEEguShrx31yu
NCGezavJJAC+eoy437d+TCMPqjEk8CWSpk5z80ZRdZ/yo1b116EcKKQc++uoLZxtljEvi3sYsZvw
CoGlUT7hy7CwYRb+hbDrDTihJ00sULbPraBLZV9XXpCWGG68p1srkdrMD/78+K9QYIBtGp3sCGVA
1C0bXyQ12y6bZyV70b60ety3idP5kEhKpruQCUMI/I0YZJCpI2jnKu0HI5A5aK6t0SCc04DRuIZ0
VLaDiBQjE8vngmrCGhMadpStVVu+RroSamTRfsPKGiziOT5VNWPIaBKOAjDxlI7SKmuxIX+n22Xl
/ZwQGgEZxPzZp8no24E3054gCliUa50i4s86pFadoI1VJsC0Oilshc1h7yRR/cRSnpa+U80kMxIX
hlzfHOhI1aDm3rFphrl0IBtdKf5CzM0jRZH+ifFS3GRORZ0gIXLNsVVXOtC8E6vtWf56rYHNFpXy
8ypCmE3YJ9646iKoZzoteR4BT7qlgzwsUs6fWT5Er+Vmz2nQad9G7K+iukdf2SKWnrSIkj2AZ5cV
XvJ0H3KjG0QnDVE6qvowFIWh416zjLJtnhn2p6NzUHwJ0ZekEOcrufsbqsPpppWpzxEPgRndo6t3
OX/g7GuVcYM/g1Q7eE29du1wtnICWXUNg1+CebGx7v/0ja2A7yyuQ3CHJRrMOeT/5D2drijpcRz4
4nB7TGheChfRlOOI1jOsJtMgyxD4jBbOSQ6bmXx/rJ5vUVRIq5vbWjarXx6WdKkxFsc+j93xECOZ
2ZTalCaMiMKgFyZqFk1gZi96czvOQge3e+A2rwVxojnWIZB/qTwyMGVs0brxr9dSw1LDW0tUxGm8
X5oJaX425VneojV0vg/WWXwfVrfwluffcQn+dapdBKfRG2RsEutMIaXNIJf4/rgZTiAgWQSm8urZ
6s5n0A7DMzeZWRveeaBOe3ryBjQciNhGh9JrMwfedrxJGy+M8SuEQj7CN1rbYcA9c0DwVxq2Swti
47UsdsPUzoqRJzY8rd07Mlj7p5yeZ6JLlY7n3/DM1RQsHhe9CvxHe+iPditvDOOFW+9Hfbz1KfPg
SUu8iHNIJttUHq+XwhZiU4lPZQ67ks14S/B1XKChUW4uv1VSU4oYfWOX3TWeiVeo8qQaM2nTY7/X
oBGoSTXwr9hGJpX0JnMV99UQSURf3radUd4GvZ6QCJu20AUEHTX7gdSDaQRZtY+zO8ZGQC92Y3xS
PZQj4OW5qq+zOoYUDmzYQTPRjk22P4/i5o7ekt0Gf0DCB3CKGmqhwMqptU9uTRAsvKq/woYgxJXw
eS+4FeDM+9nVWznLSGazwG1FxF3puWoL07Dj2V13u9P3AfQ+1KeykX1CXlzVJWOrwX5uAjErSGnx
4JMFbxR3aCyvv18xPB7/Vz0WHUHPN/q9Ykyw5amMzgoXpwwWXdeLJXTHrJSDCX2H8nV3qOh+e8Hs
lE1MLzwAsi2WB26kezHSwAwQCQMmY17krlq4nQGEUsXS2+RepN4EeygFyiq6J/CVC+e9gHGbWTrS
msw1iQrrMaLAe418YghtCoKa2Sd0Jl27OBUyGNAc5B0Oj4MaQ0HKAviViOeraySXWFjX91fKoFFs
4SbAGL4+PFqKAKotLMJ3pgEAvQm1GE8KjRCc8KgLyHSRwWXSpVtnmmsZbQqFiCWTE/HS6HrTJ+bE
dxgmQPnfspngZP4TQBeyhXcwBuYYsuSyZ28dsBb1r6OyTNmJx8wk3KWo3x3BGZ3qhbwLXfIm7k6q
/SqPm8i2IaxLe4OAMRq0OdqFBQbT20MjwWeG5Y3Un9FOrIW+9e/hzjZLwd4wJDUktmxEDA5rWIAS
53hw5uoAvd3Za3xRMovFj9743dfkcMrgACLyQiTVghDZaqLOMiSQtmJ2xc4NJrzNeEBfiUtm/2at
7ZLQEfIWmblgQWiFvo64oAbd0EQuRoG4i1/dWQZO0Uy4WTPyUetM8eSJL/uJ+zXHJMs2ByjfTsYm
EVAbOjcA7wHjDDlsqpY7FZNmEeCUx8tm4OfJxu+fI0hPIEkG4QL6Z0D8574PdZOrljv/qwsP+Q83
tQpTGah6ktyIe90mv0iubiuAbCyl+9dhO/f2dSKLwwIuRVLNWSXz92P6LEHzG7OylGftlREhaKAG
dlCcEfqWGPP5guiKD9HwqJB9plfgkTnbZ8eYxvfSSGQUd9P2T8exfhP5CxfADF4lVKpaLdu7L0z7
Pb4hDAYGE4JbSaIl4e1uKU77as6o881VvM09T0HEoQjdQSKDW3y2RZDE0lxM9EOE7gaGCpyepxmZ
VvyPJEGVIHd/1zuYr8JBJUuUsM6NpDNMXJWaQjJdv25KTMKwzMS5jl0cxVM8z0H2OPAfRoaY2YPL
Sn8UZ0SMJvyKLttTvsnL24wCKFXkl2aXOmqAL0OQ2DnmlkXtl3eYrmYCN+MtsNJATuX4R4c9G9vY
mj0qVPdr0r1u8B58DOozlEK9f+LxZPJtOQN8GmaCXaVllrtDku/s83gbffJEv8dm4lBQKzvM0qvZ
fiYGmYXgKkzbxP1hkEoQDnBNXsmtLsJH6Q5pE0GpKCGv9b/0TWSTL3hjTUr04J5R5ICE2PpobsHs
p9LiJYaRZSFrE1kPFElMNMvL5lgfCddtvmm8fsSeSQ6o1n082y4v5XHrNkehO1yQO9s6p2NoXqu6
rZEDhmM6aU+uYjC2JZMv+G8O/CYZZkRxFGr7UaO+H5GoZIn3XLMUVwIF753ji4pyigdeJa2Un3h+
GwrZ+7v9LoGiD342wxuScyzYXlnxALdPXaXB9c30pZgBSkhIibrGLxM9jOMmmHMU56uBw2QL1MUL
5DrODjiNfWk2z6RHNb/d/lby1tfwDwJvoyj04L8evkGx3JmKTWymiE8eM6uA6Siag2TcNI33x11R
r4TcWmVZRZebRIu1Ob6nttNPA5gLY8umpgva/j9pt/Mi7fS4wJll/tnmwD1HLCbGrDu9HvzQxqN4
KctWe+2PHk/hoXzz9Ycta9K5dlApeu4qMZAWLsRb8wAPEBR91gO/3j/XylV1vMtGOvF9Q9/+1SBw
DDVxPAdh1sTszDmMBezbJl3siuadsdK7MSRCzVBpW7h497Fqd0VqQNgR40riXmhDtyQWJWSCXnd+
Xftc0y/rAw5oB3tQfFOgvsNCd1mXXo8eLB62XrXce1lfB0wbsIKKPvhPGCsqeGh4JW+xXms5mVEP
F+CdNjXjQsLZemXic4a/gSUH3DjmkS5GwmVIn8RykpDTLjVH9FE6AuYP5r70muUL1bHSxTQGwA+O
ytU1yDV0zJVJD6SZ+uv1Bv5RlWLOb32HJLp7NYh3dw7zRdzMlIMsJjSX0tcuLFPlAm2hr59W5p5a
rVukipdFoNC4NGl2wmy1aT7jUBBoTKeSKVGmmjTPhBL31oAB1m6jmhhcIYPlFJ9o3cgXKsc73gAm
NTaPjAQerOrUdMvWXhl4WjVY3xSLehoaREc2nu5IYHY1G3GKQKImk6BCm7OtSa5/J8DbMZt9s8nr
k8tPkF9A4mEcLoovKXC/nWdiL/Hj6BTf1XDAqjuEStHv/j7cW/hKoX0Gw1sijiMsbpOpAJlIJT5e
9nNjd23u9i//7PXoWpq5uUL1UWxbt6bVnUEEEUa92Qy/SsIdYqA42ErhJ1Q8/P7667wFlAw49QNZ
qlPgdeHMlUSJF/vAot/ggosLbTE7LSQipb/wjA+vruhQUt22CYguJeV3gOqA1HFNmWJCnb8NoAgv
yD9NZhEVODbWU6JOKO3Xa1mpVbsVuA+WdyH7s695nASdgodi+O7E9XMpzGQCXqOS1LdMxMrOteJU
x1/a3HGgNCeuPEg6L1ePRq6lC4Qmk2iSguP7y6W+jrAXWmw2mCFxAmUZsJCapPyxU0Hw8deDNRLb
A4p0BHcqdPq+iC6zxu69InaKVK2SeFqjYvxZyr8+SZW1+JOXqPl8I7VJPBnQU11IAkguhlHikO6h
5X6ygP6s6x3dYper4L9uzjao6hTcA5ynb62VsgwAvdkyBhIjS3hNW+X5gxXPuLB4nHYungw/4696
IXvtPSUE8VPl2P5uLNfZDz4pie7ittqDwqbwf+kFbwECjBt3+JVZ3VBgkLHqrS0F4GB0UgO41eYV
YE5Bjx3+Hy5qAjuuKpDX61js1Qt/jO4Gu5aIGcXeIHgB19RtBpaIX3PwA+aWlYGbBVPXVVYYTKvq
g2Rmc6Ygaoaxvued87Pwwo2xY1Z+uMe18wW0hu0mIwOwRPgsicnaGGctKSt/B5Ao+y5F3HdZc6ci
+HNlHpyHHkxDIBiJRGWEBhnbCmI+hljvlaSHypbIxytOM5pJOQAhBhT0sCoeCJCgLXndi5Y2yzyF
eu8lHNUXTZHuWGk+blrFDv9Qnu3FFI6UXAJdx94RB6QSIUzTTWjWULTVoxHDV8sB9AGlygn4r+v8
xatPg1sboTAGfJuqg6vLJShriBLEA16UoFDBQFbGIMYBU/oHxpwf6KTXMBm/kuQC2ka8ekeE2dr1
xzogwXV1vqRjTmT3KYNyz9ooRQtPiBxrt4azwFtTHvNuZcXlPjz4ghHMaxbbfvTc6eyxU+Q6N04s
VjYl9M+/bAYtxg6iXW/prL5xFaDkMf6VcchgHygtQhZoGXb/5gCowFqO0DnQy+SX2nYQ+f4BLinr
OYLbvnURkGKFc4VtLu5DIJxiR4XfzQWfCKLGMpycJ2D7TUn553bZaYkD4Yh1xqRzsfsdtXPij5Us
eEgPIwsgvkFDJsKGofBZE60chY11lvrSm9/bgZQB01Ewu7CwFsO30bAXYvVSVk9/4SMJ1PuHdEun
ALW41MtsVDxUDosAJVXuoHOIcQ25Dh0TIwIXsZeqx6CfDv+WRBQ2GYtbdywcp+CJJsiRvuqE6gl8
sH7KyAMZ5RDYlYgbx3auygwDQGHqAuI1J05Ihu1t2aDfBi1aBLijHQZVdu//bC5j0n3HOTGFqAHg
ODg1j5U01qLnfgPT3AAw0dN0+DYq7Ft0SLu+U/gO/UUiDOXnlL+vhwoOr3r6q+AzaAVJZt9ctihs
zJmHH3WrOmGhZyb8sJfX0WcMK1lMNIGGMrJopblvn3CeeGxGKQam33gqHrimS2WUCZroYCQAoLME
vIlSLjYK1fXCk688trB5e8alT+lxsG/1XKUsqXnd2Z+i2CoCS34jOs1j0HbmG3roNxf3ko43UIK/
MTLyxMb0iv2xfDrX9RlYoSFLEa4E5wzXFlLt/nRuoh3s24xl4D+iUV6zdKieQd5BmNLnOjqarNPH
MRCWpl1Qz4odQtVpVOxYeei2DgqiOGttqzcnQ9/NDkZTtitPAoT9KIFEIj5KyOkvDA/pFBqQNhUg
jO9z6x6qRgNmycoJtrhyQkMPp4XmAHZuYmqV/gfGddUIeTePQjK0YeOqKuRUATOiBsP8/WdSzq+g
SdiRrgxvrzZHj1+nvrgOrfCceMpvpoOz12dPKdkrwJASGoQU8R6uMW6TSt5bHIrbIMF49emsA4zI
1oLw5CTLBCnZrTnKKDCHgiUIXmNQh+72FEFA3VUAQgvNOD/hCP/VOB9mWRg1ncisjATWARRffTlj
nGuq8RDP2deC3nuKIcTPoWUVdCPwJU3anTHu2E9V5jJysoCXJb7xXY40DqQ2pYApbV8Kf+jnRwcH
ttHnPk3CFSWPAlXwgB7kOiPK94teR55ztx7W8dI4Ac5BTlxV4CBmR1bETznhG7xWX+Kx6amgJUVm
UT90Uw+cQAiiLSVes7jPdOPjy2I2JqLl89JDq+06U/Z/r8cdvkkNonDf+GN6zSJWfzdRpRRgowMo
A9NL10FEl85l1W/egev0itPuoTUU4RSyw1fKeE+Kw7r9sQow4R4GISBujVLuWKbKfORNW6VYGh6G
lPFxHdtzDE71M5nZfTMO9+hoagfluauAYQxY+rkb3vK+TM3hVUBd+ctH/ojzkOkYeb2KFB+E20SJ
xLvCIOu1guLlvKtxoDcFGsH/XNQ6bmqHJQfkTAIRlrYTyDUrIHxx84g8q9tlv983mtTNAuUcx5NA
qTUJxcNoaADDn5CzUNWgSEb0WV630hjnuCGlUsf5jWKfFXFaXPaR9fnaZuMy1bI5Sre8+CRP4sZq
hkxSMrdMwJAyKYTCYtIY3Det1GORxbRApSpPoSY4jcCWHuiiMmkAmdCedkrLxpSFI9Rx+m8R2gkH
Bz9eqUi+X48HlVEaX4eyvkTG1GHwj2P/MW4BUDgGXwfEe5WZHGVvF34lZ+Ss+r7TLBW9aLOrta6t
3pUqPD+K8k5Sdv5moDL5scZuwKs++6Qh2NXe7Zu1NTT7VojVXJIiVnXV3K8E74gMNAXSTlwa6Dm7
V6dY83P/12CiMdMcbIRei1cmrvhPd6g8GsQr4+UvWY++kCirXp6GkURuOHb1AYccLMfJugXxHSmq
93aFz8+e4PaRWLaoUjqeINQgycFK60QpSaqbAiZI/hcXLHsLFtcGhJ2BkYbvUBkE1RawWk6A5hwm
sYdYYQ9+ME5EwaZDQdCiewJJVTQdB8BxtdLae0WghwdWi9IM6OCYKxTb90pNrT/ix2aWP/bQSKXb
vgQ6a288H4UJ6RB0kqobHVKzgUZa9CBsjF3zHOPnvHgwnRFxmhVzz2wsS4bV91GtiMy6TQWdalCr
j67so1OfOAKxMaJwAljzk3lxiD6XaAOdptnCgiLoren11SHVsRH3+pbMlKAaoafi0wO07Shn4UaF
ppyWEIbG9Il3H5hbOmYhYUMiV/PRp7tJ2zwoRTSKn7CKWm9aL10QHqu1Ow3GwonZAKz/AoSBgAtX
HLk1OPXlu2YmaklHKnuV5igX34CpzyW1FW3POVpaPhwZhyGESxgY1KJSmt9Q16p+goNQRmdNinN2
KeZVLn6M7N01ax82SSICMK71uCvYQhq0KZtEhLITDcFMZ/Xs/ySrEb/8vgfBbpbWhE9RaA3V8U+K
r9JqhrAAOCj3TuxIC6UP9ysmcy7mibCkVJDe6lNjiiSGauaEInJKTr0QDrRZzieePhlC+wUh6tj2
ghUFfnIKBjfJcfsNKKeQxx1aUuplma1h8qdWUXJNgSQpfXHFm+nAcy3JGleF5u4IgE9UWgiTQcP4
HtvfQbjHsJlquukgVWUTUoSoskdjL2Cxi3G8lkrhZuVLqtGGzqaYnfCODDJd9xc79O9qFJ6F1p/I
uCVF6fVGURCNls6vter8e+IzMa7rX6307KkQadO9rX5VENQyRXfxRZi3Q/xgrGWv1mswZZPC9o4l
qTt5DvvMWow7C0SRb5ku3ISFYB+G7vlx9DRf+m6ZGfnrmznqkC8k/WQOYMgF3jDsZ5stOCcbf5N7
opbYfhU3tfeK77FCZ+HbAc3lwgZLUThcf6PbTRkU4I5/EI1y94KzJMDs+nHtwx3ncJYwGr1ydtx8
isqI2Z18ctfmeINOrvFL+t18YST3DteZTdhv0vikO9MQZer6pa8OoDzJ+eDwxInVZrI4xtnLZZM2
qhAx5gecUK89mx1pvDX4m9z/QRh4ev1AwcDTfcWARREKRGMhN1OCmpUdzyZvBY5y8NAxNaPswTpU
/+pnL87Fm8/KitUfwMcx1jBiFNtTervPxjizt98RUT5ZEXdSSgV3y4EEuZQHo5DSzWRkImzeYjVv
Jz/RhuuadkaxcWK4AfZ5XGNx3JofNITgkorVigl/X2c65TV2hUOKRFpxlfl1xf/axFle3tvFjbN8
jq9tYkBVZ8buBW7tlrG8N0QpowoL8XH5OhABG6Eu7GnIqgRn4iBVOnN/wwHeDLrWYpHlZop9D/9O
91yBegd8lZiJ4BjOFk7yVTieQojCKeilaJvN9ct6sHVI91YSR5vwcfjWcAH/fatphqMMtKqgFKJz
d651pvgkUGZDSfz0p3LTFg5fVwRmiAAG75WWnoogu8nEYxJ0wN/MsvXZe+wClV212AZAcXwgFFfy
FKOukUCDAivVDdGxQJt2+Li7Y2uEeoiIl7S7PzV5I6klA6Lvie0i1OEGf+8rtb19AB0jKPGyasZR
467U0CzHK9fX1lRJQ5R3lRW50I2/BHm3hAgbqWG2ho5H1+MLIHXIeAcXPuQ9FSzjac9dcd2402bc
o1gShC/0SIRk3AvJNC+ypukItcDax7/WuKLSEz88e9ynBtsiv69SPNegkcEE/DECXb21yfKu/L+3
mBqFz1YlbNpf0pA6XVaa1FPNDJOYRrH/HqVvhwiSL3AgX+mQzBF9iILyOECbHui7k4+7tu7xELA1
rgpSCTPZUCTYZSFxTDZMvKa5yAbr5C2aulAeMDRJoOyIdpYaVzQC8uV69vhZI/ZwDabl234Nf2jI
Nuex2B31wK8yTiFSEcye0RZa7TUPhvrvjGnKrSuTGZ9ExlP/OJqs2iGbiLUU1G4GLeRoxpOJm1Mq
PyegdGE6QilHMeRacpohIhnXeq2A+tc9W07nZ9OrFkCdIzGrXp4ugJ35HmhxHagV2s0fNAsfR2Gs
1wG5cTL+2LBul7tPcHA7jUtbeYBqAl6ZKFkGKH96p60woEngUJkubu1JsXHEmO4vABqG4Si+svco
rTHfS7DwHeN5D037HFjJWOmVD6sjVSZBpW51QLvh7k2ZcTq84+Kk5ISNdJQx7XR8l35LyN2mpTZ+
CWALY5IXEvWQbzIfRU2Ocx2jh6nCBABVI77HBe+4oOUbUfQQjf1tWnam3D89mge02ndblFDbFeEW
sRNVf5OUm+wnZmoeY9BCeiT4yY4Y9rR5OdUfyTPiAb5MyW9iPlyb3bS1ANeG+tMoGu+PTWXJIws4
O/yqmsgxU4v7dssRTdnE9bR7qhNE4tAXhapVuz8rWGPMmE3V9gWPD2vveWgWWHTyMjlmJfUhwyup
lc+RYoQDEqboaZPw5I3CeGP/qFcJff92gqqbMttsc3Ic5YfPk0fI37G8ZTqxVAZT9DJtD+b8Xo/B
Tuow82RDzE0phPCx3CpEGI7uRl+OeF2JW7BafA5pnI0JLL+e+r2Oix+S53hYy+Dr5zJ8opoLiRam
OXSn7gqG2dk6fX1J7DuLi91ScL22Ipp5dMzrhf6wEmpvMlg9df2BvqZv7N0tHDKIT6MQqrtmJ5BG
lk8QCG8inh5k/2wLYSxjxOKv2fP9AM9tUbNsR+aAIgK2AW4/JU8ub7ijhgKFREkjBBfhNjWniwuM
ULW7FaleJaQthVTyh7sClR4N+MQWd0RIHayI7z4QkGX7vFJ6XmSMGWSjegptcWr9+R1aZ3wJYtX8
qF15KpLTQH1BkZSlRHZpJLEqyhb4k+Ud64PPh154kpi3BF09i7duWQWr1OL4fTtek36V5DhkaKWK
6HyxQHukfEcDhkIQ/8XoksTE3iqla0Ps9NGaQtacJnHskdm2K8cR56cDdQGeclUEU0joQjlgW7LZ
iuSUMTEAQJujazJHYxHjhk2vyWhxeC2DcRtkY8MbJaVQUrjoDgBpyXtygYFIaNJnklcEVDhmrRGy
8DEALeI2qAniwXZtVM8IkUqOdMxJ1n5pH7nLGonG+p/NxP/agwRdb0wvpTR0+1EugnGdQCPWQlm3
PhM1d2Eu4zMlWTYSpNRH6LPJAWfpiQlDCfQMAxUKLS76jIBs7Ul9cFGWcY0P3Nan36OeFvItvfBc
kAjzBvbFabjw4tmzURr+HEY4We444CZK+vUpqUtyN1PlAZk7gzSPmcTeAcF6gb37G5C4D3sggVh6
3FWMs0hCFwbX7Ix7PzzX3ltbPz9jpEM/gc1m4RzSjoq2ZHz4K4zlVV3PN8OH15vBZdlsuCVO6mKy
5S6x8XanhwNmKHRFkTiTmNZKCEXa7Q9N9CBT0tiu7sUcCk124Eb/BCpEyD31AjdIQeOjWO2L6ppd
OyTLEicXGS/FM1JQF0RbivuPJI3OTTdLUULXD+3pldNZe2tdwSyPheOQI2prqQB34GLFRDULVag2
6OA0kl8psWBf9Hf8zYFzeXKlSTHhpTsPFKQi/P6CFbvXxDezvaJAO5q3HNO7Z5MFZEKwQYYlEMAe
HUD3vbWXD9zrpNjlQlMgjCNZY1a5rxDxSlNBZRizuLlcsBtlMVbzRxXAINZ6cqfXbGT7oTpLgSBu
d6wg5/Jw+pHSSIUM4gkEDdi0znUlx3ZDNJ2t8uNPalPw9v/FtmF2cCKG6nHPCxZ0yapG5iwBrfbF
caHBhG8vKP88I/6XE+ysHrpTSR3u0ZbCG9+j0mvHCdK4QH3ONWAqh+sZ0IvTJ0/Nkl5SqKwSuwu5
pxSor/+FOy/HcB9vLyjhp1/b3kHe6g79iuI7zjP295I9Pcgv1s9TCa2pDvwyTDdQ9KV/LNc5QAAb
0RXUv5A2dxzHiwsPbpqUGPFohZlkwxgGuCVuxZAU3mavhK2cQlU7LxiE2xD5IzroJeaBoe36GZTE
5z7uADwyjRy1Ur364HT7pCspHrrn/AarD7VwZkMGTy+GPhI8HmQKZDYOW0Pzu8dyE7daarqeV+O/
b+Mk3mfGc/oRSFLATEysysM1x0wFA7Tq01pd3njqDdc936XdEcxpTcTeji+ymojK5xBtfXVTBl19
72JsLZZYZ/H6myr+21b2tH6tOyU4mjD+3nHzDtDllxt69PUVAV9jLNIyuW6GDUyIHKI772tB96Tm
9lGEZvB/DViwzbo3eaoDJXSYYOzUMjcMrU8AoTJgfPPeS1968BLCrkvb+GoUPWuB9S9KS7miaj1o
UYhNxo2B6f9BOkrYKwLu+UNRmqYzv5p1REucIRdo8d4NTMCZiUF4b6KSynqWxh2I+RSvec59EHlp
nfKpUukbJugQvl+GISsTPLCqYKy7pERaaSjpN1Iin5u9TiJi931p76ZNnuSBVbHzgojZl59j5ZDQ
yN23TxwBjRPIYXZU7WHEcF2cpk2ULNbFXs+JI5vo2uF7T/XmxR/j0P3QV1mHhAJ4rRFAupye1Lnv
cJtTTGKX9LMNMcfKB+8boxGbEqviMpUVTN09vlJSocAB4F5Z0lw00rmd01jnBiper4TxgOAeAU6b
eiqiYclda8vCeLMe0c52m2VKHnHvdiZi29AqPKK5PtsCAhLKl6n81PMwQJuUm07eFyXk/bNnqom4
2GD2gB1w1bn03dq86uiIgGP2eTME7eoSFrSl9B9T583bm8chyMJ0yWA22EjKL97Ct499fQ27gngW
vh4+VnxhFM1IS9mq3V9rVQlEkgc/BYTBerIA475ldXTOczuSt3JDXMO56NYAm4VwUT50g53kAcxO
atDenSNqxuPQIcLGbwhyuUv/APjP4Y1PNNaabbFD2lv03EtOmn40l4+mKjW3zyN7uT/SOjXBvzSL
KWCscHFR0HNxkkVCEPterNq3OTl5k4B+AHrBFpMPQ7fcZzPew4XlW+ACRlDGrVQuUkvcYZZAFLXh
GeEr5n5+Bdl2/1KbmnqdALjEHDDHmoCIHHYd+lgGwwkkeJ5FW5EJnKf6j9hBtxrvUodnQXJCNfL3
ZKa1iQ3ZXgzjN9N25pYSCasiZB6WXewskpJ3o9AzaFk+7ZoKgwp2ZUTgQReFHohgQljxsRS2Xd7x
fUV8iNPUTw76YqpqnwRADOS02Nk/qqAhsfcx/JvYdrzxlvzz3s7F6XVhtq2RcAKclBRk7gCIr31Z
rHzPk2nSeigYVSJCvp9yuoBclNXZp4wq1N5jsNMEqtYJMgbvKYG5Lc2F2BguFm2z910wKtS8JjUg
+OH7B+YjKVMMxGl2m1fPmox1M0/GKDtW40tUqnj5kazFUFkL+MxRhyMs3NNlmyVEoNWI6fJpgV4B
UPDzHhxFP0/IPJKXWFPCBkiS0O3Qaz3UBhux8BIPFqYIv2vI+EHhoi3/+3VBXEMV8eI+jhZe+Z09
uvVUL4C6HWCIwLSHyGUp4kxfnDSI6WYe/s+0ddGDeDeXo+SfIwxm6ppL0c1z6NymmcOYQfa/k4O8
OT43J0ljQnKiJzWkT0jWZXO+jWLX8zm9ZZzkX2dP1cq/xR5JNDBw275RyNpNFZjY2JjntydNTVOU
0W+i7iwaq1ME0YBk3af+n9OlFpk60iSGeVRLaIu9Za0m58D8yssh4Zb8h9qaLToxeqR5gUHldkQ7
7U7nHB81VVsZ5K30axL6cmHeHAeBJGbAnf22wVBHVZCIw7sJ1877PsHJqkCkWkZYmsLEvn7e89uD
0MeD7NOh+0luynvTdnxkz8dF7qC9nmMfhtBhmm8SRAyzWF2mRAx8kJNbSs1czBojNN4MHqZKMhfi
rggzx3l6zlGNXeLj4HC9f5mIfBlLWwiUUKoLRrupLxH3NkQMWZf8TCv0X+A4/z4onrfrmk8fOcjN
9nM0VxvpLMzaS+LFtyzXXsadOZCT0RmixZVwYuIyjCcZ1gRnhYW8BlOgmsHQ3lEPXuh7ZsVtlTh0
thdhtUAIc/kg8hP8dTP5XmbjTxnqheyugUK0FZWJX5+kztaUNo6d6iTRwW+iVSK5KX3rZrIpbQ3m
on39CELVgLe9kFi90R5Gg9sOxTzuna7rtkKXumjbfxYfGVU2zk46NWmLIBv0/ZeHDaOwn6d8GQB2
7GOaXreBk9oO+NVpOQflHHX3zOVg3l7PNAlrbcXGxQspsKcnX7G0Cs3PM2+T0QKDxCsHGWnZzKc6
7kZD0htOk4L6LIUy7WrdHtzhrtQb5WS96owSSum+jvkQWmB7SzPNx8P1aooxS0KqMIB8cVHWBZSy
q5De0jXUs+xDos6W7eO01GDF9BSy4ogK9sR8LuhcMMbgp8tmBo42jku3hyY3dXHKMWgkzUd9Oogs
b9BMkUpHaQumvxRwTNNh0+ZkdRsDDo71BFu0k02OrKgGAWIyBdDL9llGz9MDSq/WpbQQ+ndDMG4y
zox5v/9pl1NZSVSzVYTfsoHC/hDBnH4TsHvHVzp3muWzQkcilPXn6eZPw0MxCf6dTam2X8JUvJFj
5TxuacoGFZn+u1yUMZk8/6sHpQjarFF3F9lAObC5c+XuEZLOSSjHjm2IqskNNLT3OCGTJvh5bSYT
MPY+Zo2Rv9GaVbKq09DLzMdo8/7MF9x4f8FD/vm7fw7gHD769j63wPIzBbbWDQylFrT53Q7cd0NB
syokq69CRgNz1RJo1i40I7qaaJcVyp4pWQKLvY8Cm58UQXDJFLVT5ISWIeia8Oq05UPRJ0P40SI7
idRqBKfnVR/B+KmcfQ3M6NxOv83wD8sKeU2DcBNq5CpMeqF44OuHFfrpov3c6yEGpQ+3r8QLbLFP
7t/5zyQGJ9YbyoP6/nafB791cugy9Xdv+7hKYkfOrXla1/uj0ROHoAcPCbD/ckh0eDYD1rrpnM7e
VYyJzlOmoTVoMU3WYpaGV7uPQcRxu4N1DarAUkxIkz7WWGm3zL7B8TsQsKtxSlgW2R5fPDMBZI4W
VLxUBUYqtJBLdg0Go+wSZfz19pRYe/8ntkChroiSc+DolrQJN7Ps37orC/2ixvxNlpWCOit2DIL5
Ajy+ivoqX1PQqHUf2X6ARht+OMrAqogyc+p5akfJXm5uq2+s5mDyWGyPpohcIZUF2dNs1mLREMUP
/fZtvpb9Mewp+lukteotRQypMWZw1VX/DEFCTVbMO3Xq2dgzxOcPR6Uw0djH49BqWLd+kWPC7EoX
HGMx7iAIIKM4lYHQYWwp4t0nYRtD5UU55jun4Ac4YzgRrjcDqWiIA/ZRdXCpC9qd2xxLty6T9lZY
+ctM5eg4t3egBqbtTHsyHi+WaMCvQk+mInhF9GUgQE8W4ghG0kI7sbaRiZdkEOVwjqjmTAqdzVm/
FASgT+ICQQD0IlsWmVFDH1oFw8JzuLMXunF6nJcJcKRQw0lsUNKxDkKIceb+THTXGiEN5h+BYZWB
sW+W5vb6AwHPH30OFUojubf9MucPAVhA+bG5GztdgnRiFtVlVQZs3H91IilcG0bk5xuMf3bvwV8m
1PcWazS6VxyYZOKvcVe0/1IjIJRX5jijT7bIkyRBfTQqM51UgXOtUXZ6t6FzZtxyBJaAEFSYgX91
CPABUsOIdKK4WKMPBum43y6qnCXKYRRsvi7uaXIVDpDFCSbnO57vAPB77Y3iKLBFN/z+ob2MSoO6
x341MKtrDTjxG1S7Dun6pdJ6I300LmpeYnaG/WY3HZg0NV65a4IKDAEPCiaUb0KcWPhYuMOX5i3B
VGEciQ3wa1m66yCNG7+0NBHbTcbDKWFqv88JbEnd7qq5pB0L3taUZa2LGgS2vfHHiXGqaPBOplzZ
CwX/8+096fiG09xgnqoNNC3sktwvd1TCpEnsGa6iS2TT+/TpyrZtIAIYhGJHhGXpNwKEoDgA4V4O
bQIrYoPH5vaaGhASssQaZkpivhqfo0pi5OavegD0zFpfKtPtLlu1TJs2ocUN82nh4YUldq4FEl9b
0uidrZRCB82CuHFxO8ifAuryqRR8RYwEVm0QLYsZpE5XMJOkYe2zOIQJcdB+0QvvtOXE+ct1QSV9
xu3n8DUYxpjQPzmKrD7++R3XZDnFLTU5P/jA0bOn54xoI83v9qycACCtCFiZSf9HBiyYPS69WM+h
s8hRLG/BW5IMSGoWX9+UZGPRYdDEsemTaW9AnNP3GWHPtwQZtHW7ifU7enCFNhlpB6Swksck6ZpV
C4m7Rz+WbTscyscRAXJFRSf/eg5Xf460p0pIyBBCvTTxa/bol2I6Z+agIN1Uojd6dQgLg0T5uWpq
4f3Sp6JjfHqUaUPYCnBLltAsi2FdpEeve6H+urYise1sNpFlcSLv4nSItW0ZxjTCdKOCu6ChK7M7
h2k+1gkUgfQCMSnovSTb13tXSb1gynWnJVyGMw6Li7uuoS6Wm803mZhA1L1YHqGnMWLLCai7aMKY
Sov0vNw66pUxpZly1GwZtegR+VJCYqFWK4dkstS4NqDMsPUBZ6/Dfi8P2npqvNLU86M5Xr0q5v0R
qKeg3estVyFf2VHyXpRZq7vCrsF5+SBgM3gcZ6rRKyWu24hRF3+Yds6qPcbteNRBcFdh1dn3H90F
wwtx0pegCGHejuilNtKBY3MFph7M9/GCkhuRyjhfE4JonzTkdJz9CvUbrJ57i0dX6mPcG0BG695w
Yp0w29nxtZi3gU6x/bKroYJaRstV52g2B0nVyPDctmX0Z7fQ+OjG1jZz9SJFdLDKfnjCf1a7h0Ff
UczOeSC1zUC+H2oNho1+eRHGtxCZm1eZ0iOlNuhvgr8PtG5hEq5MMuyVsZE8aXOFPbN1/SVp5QH6
8R9+3BeOCnPP3ZdGRjC7LcaPIQSPrNvgl4xy9PlqvhYQ3h2vTfbo1ETgIPrU9PZlfK1F5tf6pygx
T4fbt0s5C1ShY9ezYnqOxjOMmZaTnutgTVma0YpQEZBk8PtpPtWNYka7+uRJnJAGbHLsk5BZDezz
vgdx7PbFpxlA4NZPje2QGiX6tVBNj1Cc1rGVHlU2z2aDQnHTW8oG8vS6Yi15IeQmtQxEIo3Nimuc
fxY4dSUAuqxOAfMPV5tB3+1MmMiePcjYBkBR07V2SSk1QsNysssumc/uq2dK/+A1YnfCMKqOb5It
uCcXBVtRTPFcqsnlT0Fb3DSibZxuMWpE0rQq4elQ7RlYX/Kw/VUp6NYSAOiY7yTCDvJ/Dg4RaaJt
eiCKO57OeFUZmx/3O5Jk7sC0x2Ij+ISMKQUk35JU4J3C8ZbISIqcNv5bF+ZDjxnFNJRAONlCgQnM
DHEBEK6zQpWIC7J6pdCXNOhrd0ZXJtz/LI5E7otTZma2xgPhP+4ElkujvLVhM8Wvf8LpXnqDQVuj
sySll95HgxMFaA/TgG9bEhZV38NzkE5jVFfg8A0qck8kE80g+NxasJ6yks87kHZwwxVdtW3sN2/y
hjy65qqAMPDJBZN4+lAYlN0+oj0J7iw1u3nox2GJ9HfrAL9zTvuesjdajhcgf1k+jIaxIhl6476R
L4zuK4aSZ0mPG/tG8FmAMGB4R7smerZeuuZS2x/V8uJEuhnQEexBUkZk8ye8LEB183XQckdCzXu6
Lu+t+5H3evzv7IfQutpehRceZtTDLQRQ3LP9zSmpfWl70OBFXnjoNWFXlV5u6Nx4RTNfXrfpBmIQ
o2MhhqsX4TUHYsp113wIMN7et5lBxvu8bGVARpUVdjuDsqHl0WfNIXurYJ7dr1t0/7zMA7i5ZZek
ZvamqOBGYUDucguWXKywPOIzj4wCk6uOsD1YIm4Lmfjsle2zwVLisafqyxzJV5j0ARquhFxcP5vd
zcR7sdi6AE35856C3rY2gMJYVnsz83Mrdstu5wy8dPfnH+VT8F9YkULa2IwYHuNjhWuav1aAW2Ee
vgYmhV1g5EKsuQcFEqKHiedSR8yW068wccgLQ6abjTRj6zbhA293hgr+NvuXwQK3vBtkgIxSFWoB
GYWh/DRnmbWL6dZTgw7JrUqXnQoP2kyZO1a5YuOGH9rMhLpdEONp5sbWmcs6UzBFcgtKq7P09St6
coelCrlp8fU/3LHCOXlzSiW09RCNPdOh5J7LouQITa/rChtgUa3R4k0ESUBPKYABFUnhg6dUm9DK
ODrt85nlQVaSKSqd3IGRKwLTZc7bf1kQD/XTmx7mcZoJCDCRmakMbRqBfucFt89BvFqL8V0S8iR2
HMsGe0CJLqxzqLVs8WmztpPguu/sDVun79M178sSu8qrdWQEOo8sd+3xddwUXQwjT/TFdRnO+qtO
9pe4+ja3CvS5kC3JzNj61VqU9DT+mqhZaUAq78ACMNrswy3E8FxNK5tOAEFJVsjzQUGA+LOeN+3+
HnRqHlxxr25dL47Gxx49xszFSEb51ULWR2WuMkGtxLBTkLrqCUBgyXhINhdA2xQXHcEIPtcclJ42
A6t1psLmFAJpqNpT/yueLS1M2XWEAyPQL6+9TYx18OzDYSytq1teExTdPSbBYQqWZSffD5mDH4BF
FVXkeoYLHXNqNrSvPIFZh9fA770nQFLI1JPUmZPTIZvVZZHevt8fasINRMXEWmolLCodgmSTh6/K
3jPASPu2Qcq8kuprBr7HyFMHmHINWI+93RPdnT957QlMafsnAHCjm0BWAdYMSizH7mFztg7snip0
yUyLYvl8RKn/dje0o1ZQ6ncCAQ/P8mxz8Pv78FDFLp+4DtIVByFoh9LnvPSn4SGd2MgFL8renanU
Ek+5muZnYjSOAbZzuby3YzVQPWKJybzsnXuDZcwGFPZYPpwY0P1sgQb4NEfOS5cX1cSkvyjqaKPo
43UHnb8DA7IeYhq+Pe9ylBeiczgl0OL39VV/0tqsh30L/vk43ipRuFuhqjRW+kLuL2uvP5K09xsO
O5qEHe+yqhpt+rRYV96KebfVnKpLannsFjvnPj3uqVJ13Tjq376tXUscEDHePQjM9n/jEIGl3KiB
kUqPAoa605qZ6hP8O2gHtYj1b/85R72aZKo4TR+iQgdTQN4PRJ2dv3HyS1BYof5VgivSsCDDxyr6
Jp7KbTbiih/LrvuvI375+HIe6qz3L04PthGSbw9dwwgOequZ9LL2LbeAAO+/TdoS2qqAx3DiAnIZ
/Rl1H+Ya1th/+sxFKlgSQ6S5dTlTaeDf5CntjgLgLHrZJ9flP1lUhfh8Ow9G0J55hx2OycX+ka1t
zOEPfyeLzAYs6nNHgsvl2SdFamdpV85dZ2/6GPyc+/s08dTLRNVuJ6s0xrKKixFgttc6zvpm2wZJ
v9YINM9AE8idnDq5ETx9YmGfi81nWBaO866kOvPlIwhGIQKe1KQZnqyEX7jG3Q4XGLq+lVbWDvQ+
Yk3rxWZ8kmNBsxKDlASKhuuLIeidt0f8kga+D6qg+UwOnzTgKsJ/vbazgjRAs2UKt8jFKTcc8pEL
4sqdsZSy5KC+AwNpaMqyrvB9M7ePftGgYtu+vUQHv5zbMauX/rRJ3Le0mGCrJVNirBYAWt3FXT++
NrEeoF6gfTn1XQC05zUBeyYzYJ3sD6OWIA60raSlU8oyDSm5TOOjSvmkyRw1h0zjuuvk8aQfTdqn
ZWhCNM+pUaHfbXLTw1COns5lKxyNwRHKNQnYXUGcsiDAN6Eeco/4xMRWvV1orjQfuwptA0Ag7zSy
yUOoyseS2uAoxHCAKOYcZhEsxO50qL5f6T17Xkgo6G4+3yFvPIOcVB6L07gUFTnugtJmyNg88Fxt
dyBu1xDE0qGFKzuRUDHPTjTJ9T++W9P0xJXz9PlmJvMbFH4jlNCtVjABqjsPvWy9AQNMsboXWSxE
cc+T+PWA3TiYWSIRYVenf73DfNrDOmkciMksM/LRU2vC5YBZeTWEcMNUD5d//lsIf0rv3Nt7OJZ4
1ES7y2KHVEmcQx5+dJvixLc6voASn1dAxWu6HIl2caKDvh6iAf2nNU9EqLLHnLenMcvGNrYpopXs
/UcZi6rZWQpE/a1XZJpk4iO4F2hLT+UFHajkZfVy5YyyQgVxVSbY4XnK8BGiUgCZuIsrXdPbioyA
scrxzy3u1RjizJcAIbh2SXKz8LFBmh+RUG5leMGRznXs1zEBkEUK38t9Fl+SEW2a/CIEoahm+nEm
AZhefzxVrebxj+r0aT49B3xm5bAbtkw0Uzlv1AYx5pmMn8LEyLaUGuskeNaDnkUi0D29bxMhYcQJ
1RhNMvkf7cTRURHZ1+/h+sJVMwwXkmFR0bE2pJ/xwlH/r15a90ZD6Amh6obwmQFvXQpTEnMcf4NV
BWhItVeMaOYPam0znjRGbIpq7TX+fgnbTHkzniIUrzbFpWyH7TKSIGnpnlQg+d6Ae86VIXQQLUf3
be6lSGBe8s0fzbeagAD7S7nqFKYiM7RIoGghqVnvesDKm2T9FAhbky5o3vBC2NHIuyqkatpxhA7D
rlwNnLt0brCL3rLwkKA/Ry7aaLC8cMhSPZorvBlHNsaW2WQ9tB7sElQfIeQk2z3ZFWwK82QGOJZv
Bld4O5Ppmt9b88wzlDtP7qtgfg9Efibz9cXyu4VPrDwP8LDLkgLX4Figi+5Z28AZRhX200cja3V6
Bbam6OBwx6jDhWPRwdvdArSGThkKhBW3lHffKJ/iS84XdgEhVJtYqb8peIR3EhrO17jGh5pen1Se
+68TNAuzxgYRwziXKVoZDUdmDqiG4CaL+J3yVC9s00YJEMyg2JFAu2cyx3MpEEHdTXzgQqd33WOV
fVCTd6G423lNyCTlqN7zVAMXcNQNU3B1eF0kp6ShOCVGdUWU4F3SbLoQlfzeKOGQbRzxf4GubK8i
qkmzmaBe7djjkAtMHfeDmEpXNGhiGLa5s0N1vvMG3qUgb/j7mJYUJw9cidPXQ3KUuvmYcBVFD9a8
0VxusTbZUrGkBaW0TVIqUYXYx2Ez7HePheD5wqPpeYJCELeecGS4RycSiMrfSrgvRuxWkOedcYfd
4Y0i1xX1FPr7K1+mGmyZuAUxNgurdiPwL0VKfNihQ3ZnowM6wfscWXfBZNxIxfDlEP/cBrSRVFXc
LRhxbF+ZGm1J+gRx8fivi46l/s6trKKfOrRWcWEntNWAkkYHR19n/ko8za7Kn2rFPXbSEDQBSWDX
x8QjenR+w9RtQJ6tHZYqLto6hF0eUCJYvKD1gTFNQPW7MS9xrONCxlFyaiI7QPNPGhAEJzlNo51w
TikBUylwJZ9OOim+vPNnAGrNwV4OGtL7vSRv69zr0Z3t62OWWEmd7mmzK7nUDlXYLUV9t0ZsPijv
XLOSmb3uYYmpHw+r5qJX5e52E1p3Km3qfQPqFZ3Trna4Z5AkJbTQ/2xLbo3c0ydTgXfwsVMsdwlr
zCYfjjLDdZx9N+WO2j6k3biSQwcjEmQauS/i3AArLwRBECwakiKeEps0cXNhiapUgyqopb8gqQzA
djIhvd2LRms01XUXJHaKTo5OD4JKAX6MgHwmN6iK+s9PW4UdrUJQ7t9ytCf+eVz0YOp5mbw6m5d8
HLBe9lR04XQ084BhCO7WGZfxh+2+N9/64XRfyoH6rvvf2Ho2kh+wFN7Gqy9hweCaIV1H07UYydkO
yjU2/5bM8JSdPbAcUqzzTxp7zths2QGaDFvKoURlNOT2c2yw6gQtm1yrGZt0IrBEyrKzVnFF8Zug
VCSe2XpWjk96/QFNB8dmWCwhdg8DW9KVuIKMxIEbw/zGAUdgm0VdVO1laFHV04/jXQAV+qSU1H+V
iQwOvy8uCQMSSFbgyV4oBii1CYlzoU7RomaZJrd7MhZx4BdmNiPr4ryBG3ehecWdI5y1ijX4sLam
jV7UWAgPB8O2K0K2lb+eCZK7pk2xlKnTDGAwZA7pF+jOVhkbXy+EHZ1VR+P8pi19M45Syix0mnh+
iBTBIgOjpyvqLxz3mmCMoa52dsDkAiMn6u7eyFj8CCwZnf1yV+9jNN8Oe05weVTnI89lVCW735LC
gryev6fLak7pgyLFZSpfyRbo9fptQNU2XqDPnmgkpKqZIpVuRXFwrHtb5sTdbHYoWRr6UVkcNiBw
PBI/+XGRGBgwSgcm0Mi9qH/KTzH88b0k9PHcrqxBcviZLb8rjm50pbSP80sPpqlwOkMwYvyTW8Us
Qy6hoiJhFZg/BElQsKKADMiQuKdoW7JmFECTQFDzbttBmcbbkVIxuwvKY3ZAHpFgDQCpwRGAJ7is
up4ADMTnFgqgnUw/SLbD0idUk5CS9mT0On04oiXIfcRASx7MBSKrBBxyp+MCgVZprBedqwza3nV0
2UvtZWZWv9R1XPYH33UkNpj1iiUYiU6xxHTdkCqv/Dx23vR+iIZWdaYkLZV/GY03eIiuY7oEkDxY
8WiM4ZriDqodDadCPbV69r1Rd3MMtJrb1qg4J67NyBzLsAWi/nXl4b3PWx27fZwT1TyFAS5AFmII
c8eE+ulavfqYZuBFbdCUnduSzwIWL41Z7jXLw+MAIMFc8LClL/ql4FguCj3UeGn4gN+hsn7UmTxV
vwImZa9nJAE4U62EZAm1HoHtFGRpJb2JoBT1JPZEwnva1GuKeNwcSsgmOMrCaLpVl2lF0Jy6EUpf
xJHthByUCW5ye7yemmQRP+tAgfXYMu2vmwAIjtAM6rpiW1Qe8KI9+srYo5GRfcAiKlmPqCU/BhtT
hufdYKzDZERIYoEqRrNWtGDNQwTo3eR/XVdI/UR3ZhJd3YGF6h7oGP2KRP83CIvExlNr8SdIjIsT
kMOnUUTL1GYQZ96dNbvmbniQi8RpqAddlnmqpwhxEnQfFUL1HllGEzGT7E/NQZ8afLT7iRS1Zulk
GWNwJbgNMEAtimRftqZhYWkeHQCTj5oQOaUpRM2DMV3F310HlDpVw8S47JNxl5BpXDnDs9s9B0iF
g6vs8qLH5ekWE2Ht2tBSd+wViXl+12xerYB2q6tWltOk/gZG6womjnSCKv7eEJUnL7Cjy1tN+b3a
QfX84XYDcislNph8vAIVjd/stnL2aw4iqeqmdtyiYmv5qEzRm3F213i3R1+aAennhfVMNMjktOh9
t+hD4bWklg5WtVJODjbbdZnDGybNcOq7i0zrU8hVVbbNTJ1XmUi8aVyvkEnpWXyg0qqLmA0rzS2C
y8HUWXdJEitmED+7ECkjsCZbeUWnUkdYDw9tOre8Q1MJjAjiCiQn5mVHxVaOCJZo72UNX9xoLx82
fxCrbqBQruMDGu9Ydb1s9KqFn52Bzp8GaOyIfvoWf7GQO6EpPF1tftftpC1jgFMJwYbvFJgNQ+Zv
Xd1VdJXzV3CWdZneKNHNYSFTeWv4XNdIK/aUrBrK6s4xKS12t7xS+Bt1dWreEQxVMfYlCvspYBmg
ugdLN8OpNbBK9BW4JmRoVeHXbdCux+nfQ1cOoptieWIehocfhKzKEm5g5pQfzPo8o9ujwlM9KxWa
QAf3C6IUXdD3rV7kq0gxYPMUbcUnJc+vlBFy+2awc3Jfs1CY2vtxFLAk3gnH6H62FHmxE3R5PYIh
GNt6LwwNgMkBh2bDk6OoNfbhDlZi3vjK7sg8Z/6PJ/g68had9dt0IdjafWMyOXQbtyRVl79ofPLT
vpes/0/C5H5PZyHHjyzkTTjju8q6pZHy1wKQGQzQqDkz3kVSh+WQkRpQEvXXq1E3xKOV62XhfA/S
/2jFHFSyE0vz3qVp5YuZvpCRQN/NHR6L7Va0RWDawudJKWhDbTLrz784+MnTyGvLe67ywV2P4Isb
EbFgrtAuG7pcmoO/oE12c7MfX9WVSjbEQ+IssGpI++FD3nr+xKJ6XC++H7ASzIBzt8DDzmETs2Sh
mNPk/C2ngWgzLDRBTQDwNHRNED46PlE0R4ZScWvhtKm6Z6TFK0nwV2iqGuu19zxuVRDRuRvs0BAp
eIzlNhgPdPLrJoJa7gUTG7VSkWFcnMB8jHLJRMLpVw4N/hpOhYKIy3uee7PMrJK2dNKL3+62osyx
k+f2XZ6Nt7xMAMlRz6rk9pO0XdZr4WeAkrODFkoTWv+XB7MQU/kyMxMEtcS+4tCJAZ6I54RbyEmG
ggFzB7Oz4+qWK76cwPI2EkKZ5iTEypSvrHfDbV0jTg3Bjszu9xHaQLh214hnulE679qidka0EUBU
pOgYtCsSvJBRKp5Z2VfxIh+wj4PyhNDruPU4Hz5gvE2vZPKmAR4lFszFXPxUm1ifYy5WHo26Q+pD
rRBqROMdTjf51NGzX6oLy1s1NCzIVCSqMVZwFqNLQC4s+xsT9y9QZrKamsnbHb5WlArwuyDy6mtX
ERhc4Db+He6MSVcnhu8ljIw9nS11nJ9OQiIqXmN5lqIqP/5rBor/bFObuFxUEzBDjTHk+vezsZ3o
BrYplnfOZ1T2mhUzUNesKvknG6M28J3HCgmFk2S7D7+Z2a9LIBCPoWOIEgKxVoe+CJBrR7FsWuPo
0jF5B6gfIjogvDFku/4SNLQ88NHOXthMnqdSsuCmZRz84Xula9d1cLG22WtVsFbmY8i7JLNx4IW3
Zp2JEFWiNcybQHTBYuEiUdGvYVHO6d/c3+dB//iz0Rr/aT5wRiwcu6ZGrYlsxHOiorTCrszNwNh7
v7F2wOCuIXa3IMamxcZ96SVsN/TlbRWha9/C0YFMXtAVZhnvEsnAWwCbjx9j9YJYomVvNoGVm8E4
Se/ed16RAd6Tr0nZY/37dsEFZSk2Hn27oIf88mObEA8NkvDOU4QVtZJDRqrBUimHRv5JM1DYP97t
VYxe7z+7XH2t/9Mva3fVEMUO4L7Ewk8ixzJRRe9RYbIIEJUSjjoAXGWK9rZkf18ESkhijYJT4qlD
n0DTwGv4NkrEidUxQVEZFihwld7+kmUfHPNSQPlli7hdzBHOxdETwy/xRFk1VFRSPNqFxr4o4x+b
BORsJ471/REzZ5BEBKRjM2rcS51qBAovpGJwo+ccaQDcdDESGm1MbHiHJDdumoJVEE3y2RKfpSwL
bmyzLg3zYTAQGd9OUFQTJu64MAK5/pYrsJk5psNumpkVu/UELDqWG5REsPWBHaLq70TIdz7q2lin
pLq8y9F/oqTGIayQLgBKHX/Sv312DzaPbxHqSUrjexXvOl9UMiIK4ucrukwbSbYJXBy5RZ4xO2Hv
iaoO0FEBIl3NVJK63RdYT6FjRi0y3Orj/dUgCPA09OGB0b9taz/Cx5dRnVvq0ulxu2U6KlnAHqGr
LQ79nXj5qfQ5cjV+o1nhuZticWRd36MPNMIWGmyH1B9QFKY6yq5Hfo64iHp8HGH8eVgzlOemu86K
5o3v2u1ZcDrqlEDKN8JbVrXsDAAJERP5IR6zlTtDnfSyxtBwySj2lfg258pIimZ+n5qICSAQ58mZ
QKY823+nqgahEej7ABOUzqYlz2rk7I4b4arMyrT7Ljc6NUeQVSaEB0DbAtF5Ie1lqFKpitf72lzx
NdrkXYSU2E3wXobd2PJ/TpEquRlPCbE9e5KSlRBYDqIyheQGrHvmQKYkybtNCKN2pV09Lv65WxrH
6SekSkI0T9nMCqaDjPEPnGGKg/ZvIf23jjuXoJ7GBzcFEOiUA7pi2P7JwtTZWGSH9b8WbmNOfcWP
CQUR/d9WK+A1iBxQsboqF06vCyz6+Y8ZNyiqoaSRJtrnc+wujGh5Bo2jXuUJGyU79cA4/rz2SI/E
UjiG6SRV1SLvo3AZvK07qvW7wri2SJXu1pkAotXXHi+u+T7zp9hiIZlPn3CgCeTUjSvo7w7BKP95
pOMqbHwgYT/KMTpqu3u7n/kXZsAl+A3MBOZF4opJIjEDDxH5n0HaDhI9TGGR3sf9xrpw/EUcUfE0
4ObtojrfW2tXzDfrEpPWF6osaYpTbaWwBvHS1Aq2/8yD6H25gcWQzfkVVKlI21HMODtzTuE0hhQd
4eqF8weXepV0hC5NOtnxCEPvhfPZQwaZF7XIPoFyJ0DVrdmecbeAhNow5FVNi/f7Xjoxt+9BVGDY
v/2Z2/f8TP9vocLeY3Wahd3VVM59XgimXcF7BBvl8amAIn/58Qi2aT9y86Go0/FHmNEXgs2sPoZV
3wQOqyFBKsT0hHVsLBFr+LehT9RPweOrFOPfnConRk5ZJO92IkrCWO/75eJeUWZwA2/PmF7GSPjV
ezJZxTx9zVyFHtcR5j9Op++5qYTB19Sy3WlgNB6RAfumSfrleVdTlxBz1W3+6GaWmOoatEtIcXS1
goT8I0CLmpmuyxdD0JpfGCoFHPNiiGdIeRGlywTTh8dHqSou6kI/t8R7fZ9UiVMYGKcmndtxL2k2
KVURDyNsxVc639oOXSWiBUlq9btcSPaUrGGYHgltU5/vdutJTjtOgPjfFpZgVsqXIcP3g4YiRQdL
bg6fS2MlO3Ta1YfWgL5FJ/ECPEk+cCxJ9eENm2tIt+TMZfKqg5VZ1EyQqmRg9qTE4fhhXlFZ/6US
XVLUZ6ggj9kd1NsXr94RGiG+ykSgl9MDdM0YtUVo3FKFWdxK+MBKp+df9t1qD9gLIN+eyRwRcdJT
NUzz8Taq+f5U8oOR/BexAKcuGBPcn4msUFtWCkPx7496idbdIBYpmQ2rWaOHir9v1e2RkNIYYwG+
1EmT0PjPUz9KUHs9nIYA2TdYuZcXwbwNNPKsBo2NSbMr4yf9NCU7EldPmwGoKEFzNGKhXlGaceSS
+wkCQBrSizR+Pxdsb7MfpIUmo6ZW/i1A2Zxjn35p/B1GJQIoVTltXdPwLE79mUYh033INfUCTghn
nSELReiaPqYuAlk3y8rN6FwLuxz/nN4tsH21AqyJmnhuhcd7pueLq+avB+A+DuQ5RjXkjmH0e9Lj
vF3BzP76G56MsEjtDSk2TjFqfozTixf78AjmLz9enNwBrIU60R/KwloBFIguteUSgMpisOhmlTQG
EMyz9BlBvEmPjfQohFsiAusxY4eq718ATDLUf21pX7rHGlC2S2qKKIggPMnzEEoSK0kuByB8pn9+
eFLjV7vZRBqoRx92jdhhhdmjutTc70YwZLHtb5RxHKSfL/kPwcBaUlg7jde09tdc5X8mcfJv0fpy
i1NDpxiO3L8xcQb9A3w0SzBPbjETK7DDAr3lpf6QxkQgXtBL/RAX7sADQ27P553TNudXaFUx+jI2
ygHgsC8H68kqsA==
`protect end_protected
