`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AMFHcUguJNyRB27EsXJDDXvgepsfa+sF5kuPtVMDDrKzGug0qI1o14vhfKLrIiNG65IY8e68Hg+6
PWF9Gh58/w==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hstu8NWbOaafLHc6VDTQZya9B8AZ/6GSRP4dnUgEdpnRwVc9AlGAhUeYZfYuX0H9ccrUSK3Uzvpa
2F06i5/xjoeY5j/ppBg7dKDMlIO6qTMq8zoOCWYPf9S0yzqGSnbkhNqS3C3x9eHh2rKBlHaHun/u
Gyg4NkFRKvWKJkupono=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rbYWSeQ3muO7VIcUPxvBNSfMKbnAui0jqS2B3mpAXwGEivEP8oeGKyv0bkU2+QY4ICc//ofeWGpW
KGwLYE7Aw1TgBWMo5XFj/JHZguPA1R2LfxSZ0fVM+9w3Xr0Eslxd1+HWC6PXq0ZZa2xgEQ9GmItv
Qi40Y4lrbXyp3zOzaZfIXfabLdH0BchLaoE5DfFwtrYcjFBPfnwG1S2jGSBBqlYqT1/IHCD80vju
811T/3iIrwciRj1yb8/SNQC6dDwnpGhpVdvVkCnhTE5nrMO0tbIfBKG51OjXUqnLQLEXGVcaAiyl
164vq1g8aFgvpFYwjao3z6LVRZkN6NncSsO1Cw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lfk6FogbBop8ZAB8hwwNZJdynisStSwTz+hU9l+ca4MW09f+JnP3Pw1J/tJWg+bsvW/Hzfu2d9H6
g8r/B+Btqcl5vVOBmuKiinwbVqmVEWH5LjFek5D0apWKCWgQF0sgHb+KSR60beW4XPq2ylt+yJBp
IOY+/PJ6zn/VNkKV9ymuElTeME9VDFYW2a3wU118zb/91anNqxudFdmI7MiChlHmKzMlcrWxxAAk
1daWsvRGSWguKSADUdnBayWTHep9SI9w/eOLMhIPzkDoTD7gxcXzwY5BufH08XkqG2/UZ5+xSSQJ
bjJZrLtCuDw5RAbfxGyIEwPE9XVZNOIYuDSwqA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bjM3tjYQ57+64mUkuCAC8dStVCUIMc2qBJ13vKXBpT+ZeYZEnSPRAetgfI48b6isXgjtzmZ2Z7pg
pU1YyFUDdYhUZ/vCPsb489sLMNRv4d00q094bieFIgKXNd8GVtqcx1MYKVDeS2JaxM4hQv1gUXvK
WNhQgHPugyzoie/zj2M1Zlk0EOCyomtIj0cEFV8YqOPaHKb1zpU7Cb9iWKRx7TJe6mTexXu7qA6i
09Am1gISBFXfNoZqi91X0q3FT+rTFQXsHwwwllbegTvFxhiZZKD3uL9RtWtQmoC/mX2WbwIaN03v
xMMBmmE/Y6k1SsKPeNo8lfqksSMAynDrnadTdA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Vdkw5v6+DyKm4yWvWTuXlmhbidZF26gcfo5EN5DjPrGbtL//Xpiars8PW2iXMiQCutHTMMPFLCeq
bSS9FZpaE1GCFiZrpj7e49ftZlFAOSu6XfjVvchMe1Ps2fAL3Aokel5WewMa/ydL2FQh0f8ytf9M
ChQPPH0glqeBojXSADQ=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EmJebr7NnG/EE1koMmRFWUGffc7WTQy+/es1DIExJZFeIeTxqJ5iPcL3y9LmCy8iAS5GK6Dvp/yO
REXFttgUtkwikmXyBIHiXW7JQeXiEoDXeuUZKxtwdPMnyiyJUfE4MfKdxTrl7plLrz82zmcOOUYD
KLAPo7pQNh7Bxw9Uhcx1RlK7CyGK1HRO/9f5uB0Zxg5y0ocmNm5ZLUhBscayZvo1qr5nDiqCO556
H+7WJCSjEHlCVsZfcS8pDrBqQ74Pk1iJbyP4aqeQIyY2egxVJwraTBE0whZ8Lz3KNcuckgVJ/MeW
sD+rTvsmPz7AQ9VXGLwNyUIQhzzDW4sJbqJtOw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214080)
`protect data_block
d2ZPMg9lV9DYrUgqmi0P1LeY5wzH9nHZhN9VJxJ6QMSsJp+9KAZgeKM5yM3ANPtNpFDN/Rifm6x9
k3HQbtV50EOdQfLGxvSJ6TeRJegU5oyLW5ulOn561rITU8VWS5UEKMnrW+ykGGE9EtEeS3HLMx+g
hUEnzMA8kjVL4I0v9dDPpvtsUSdKxmBdydqH9n+tpybIc0mVD1CYy9v+yuVaqWfHz9WqTsPZ6eLS
6cLtiIWv7tMeO16yEQnjegZPdtVI92Kv8+dlXoWgSnn9hJI837qbuUuV8uCKxBGSnoMhnK84mmwN
xKk9MZ8PLrpW6QtcdqlCp8JSWuXPzmgEPXOR9ZRGrG/tRQTJv0mdgi4rPtC0PuhlDpoadHZUeydW
6cM22l5nW67CwevtKvfA3hDLcNR8nxy0iSRtvEBcZG0ZOiPO2yvVobVHIyPWEz2USYQAgIfv6QZO
9B7lfQ5qZWCfxkehXHSciPv8uxmEsGxm5zLWmqiVec3H4MaESiG4ZRd1wrfS8UOSpHCs2QN6ru3W
+5LEmPiojArWKt3l1vqb0bgMfl4LMY4KS469FcjKgDDyPSxe+zDMrPNiOJYDYGyTv9ujKCKE3V3s
2MDk2PWQFfZ9VsXLRr5CzMB2bk6QpT4S8/5Rym5UcezBGU+rBB/8RDhPfHype7/tFUoLoc5jBTGH
ElYJPq4bvn2yVaM/G8UYY+NzF9YaYp+ozc9nn14XluxEGRncq3H/3vbC3BfoCfvdhyWxZ3xYQvLm
tbWuRXw+7pXpuAB/0nA6kQYv+mMQ/KPHrpxNz7L1tk+XKdvqzW0EItqFx5y63hSHKQow6qOf+qbk
9IPrHNZRiwbMjhdhAUsXt+5+KbfvBlGmHcsrXAD6UwEGPDzA2Os16huS2ZDwx89iHan7CvNxIJyd
urxCtedhLm6svDFArcWWtElxyQlE7lMXZUgZRPNfBOk/PF2zbLQL/K7HGBe44t8a9O+KTPdrqWSI
NouzgSrgbEC3Ztw5NzELKXazzKOHHaHa7SOmbwx1NB7pQnIQ2ZgyYKbeSJa4XpQW7JFKMKb71o3j
eHAXlI3ay8RwMo3YqvS+XkEEWAtBRhqS/wrTPFefiSMfN9Yd8M1icoQ63tFo3WXU6X3tAOdu31eA
fkc10Y5W+SKcdPJpaW2R4wXtWV90WMa6SRspp1qXZdPQ1R5ItK5+V96aHuMTHub/LwRxH4GOLsyN
QSFhROSGSGrGIhllWQ/lIJl1nax1oeuvExfKmg4dUunCKPPcVWB4PfGJpR79BXU9wDPUCsnGOQ+U
VJwG6a08oCJdzpoPkrOZwJ1IQq7AJuDduJw/77lAlZrzNZCNTlPOgGD4yuTuD9Jtox2XzyhI2p5u
yCthkxYPvthAlTpF9ZKl421GSo7SPlXDAIhgkt+WhncSNKC7k1sY1hxtGBAzquA5PPYONVt1Sw4x
O05MSQyVYs0/J26QmfAkqWy9ikwCrU3nV+sZCpkBKlJRCvOvlpLE8kWrN685F4ps4GHD1oGbOTj2
IGz+b3LOSC54LUzWNet8BjMfH7vezKkmCvP0XPSQbHzVJz7nqm7T7B2zUswTxYLf6gCPlekXmVs/
gbqwiglqoxXopG+ONEUDLRAFgfEC0EWPbU3CKZSg1QqyQgiv1viLoDhlT2x/KfqefMXW3VVhUV+2
5CJ0l9+euvvxHnh9a0Jl85orZaNjiuiO+vXArFByuv4ta8G9K+OuJYeS78chVBtVs/Zgxxp0DXD2
L4PZwqjjRyOnwi4TA3yMTfmFVTfVzmkTb9XD+JbvAMDCg9ZYeal3nDyMHghUC05lTyKpr5/e8945
YgLeTasleCMSk2SPlWwSCcHWEet1yO+gjRXgPQNKh4DGrdslPqNwNbRxqPE8xbwWz1gy13f6HWYo
EF7Jg7OgZR8C+t8PfiwLYJbPFinPDg6a3cGQLIG/lvo4FQcz+/ee9ghewC9CotyVzuUHgrusPByB
2Bc6g81Igdw9WmqsUPXmkCwfUIdpZAY3GHoCvOUravvDUMP7nUwp3UVNDjrGQaEhXAI8b6mLEbtT
zFWgnAqjD2/ZLNdwr12pa6SMO8gY4KRogsSW4qc/CFVLzh9KJYTCLZdt6+y4lJIEVVNav3skW/OW
UVZ73bnxcLwx55W30o26Dk7nphdm6BNTQoZNt8f0t4CPrXTQPvNZxzEIxh5IHoclbxEiWiKbMIc5
oNGNWT9o28777Tj1LtnczA8UZXtVTe6knqn72nTX6JyukvEa1KCLYBRdC23a2W7EOV5sgC/bk4vT
2+5bRQHGzLg9TBRVFB8uASl9aACK7ij5F4IFXHZSVd4aYMsze7H4CzIVLXXd7s85NuFf372rJUH/
G5nSnip7Ezahgp6frj5ESKx92JOCan47YsrGe6zOWWoLRjzqbW+iyuJrvV3Ym1D7aKaXR6j8j1ZR
b7xGrE8p5Sfd6DzHmHL3PTlXVYloQxg4prnfvavf1uOmhgoGA5zcib0wWVxdR0borE628Mf4eoXQ
oFYChD+px+jw3h/34NVk2xZqEUdbrgHfrS4BgNXaTzQT226Hx/i8beios2mt+afHV6UBGfnJOeBp
Csv/YolTqAZ/VzKVmd7Au0F60wVCE3SXaP9dB8KKxIzXRgZTqm5NSVOH3yIYTQ8dJak16EZZeito
OS+/182hhzXrMTNDaLHjtk760Bas/7G+DxrH8/EwVrIcMBDyVGM4zsEJb4oFAajrnz++Un2fmRPj
IRilLXEL1gX2j/dCd7hnESlHoC+OQRimVLVe+zs8aj362l5a3yglV1IKBuE0YQC9/0D7uFU49t3l
SF85ByYq0bU49sDvt6+j/rZ7GdCn70yMpduna7vO9bFRFJjI+rDGWhjTG2jl0Ov3TFfCvwoou9y3
y5Sfj3D/kfu5jYuizlt70Qt2PnghxmNt78NOoPdCeLciEE7cLoKtqJhzhxbEjIJK6vQe7fdwHS97
QH8iS174cktKnTfX+hXj9X0ZtAq9dI8mim14/jMqYxpSg+Y7zhzDOEBEQTEI+utOvJbsuixSbiIX
s5VhWwsjEh6QOc377+6goJ2d4fyuLY2iITiaXE2096bXoBPLoN23bavlvESnKGHCpD9ptACz+qZA
RA1XkRjXBNtMW3FTW+oBt5Hyyv3l/UVWPWN7kiCz3onBEt0/KqZfDxNis3N1LY2e6PA6PjwLrntL
J56jf46eO4F5yjPIeQ2FuSOA9ShcOWZI7kiqxGlZUAfuHyNYb2cVinahtSIxCoP/MLoaGAdN3iFp
7G2EEO/m83YyNLydYVhcrmnC4H7pP+dCQ4+TtBDIchub1mrSKdkxcQVqFkbrJrsVjWx8I9aNf5x0
FZzDHOOi5m/OWPmv3bLrLMY2eDvxI2eM8nMuKEh2r3m6Q9h1MDIKJlZKEKzamk4FWI4UW/L7E/mA
9yvWyk97Ih6oOZSs+Sy/uarVByLn8qqsZY28kBiuMd3Sj+hs1tPYGPhu2R2BCRMcrlVs4k/51TuY
2GYl8V88t0zos8wPSbIVXXHeCKx2N/csZBQx7PGFJXU18Njptrkvszbl5R9PPsSE46waMrXAocZf
0+BgLrMrrw++xsgXk5Jo/i/NrGwjSqRaUL/gM02KtrkJttXECfss7ZvpKgAzp9IAWwDAk0KqdnWO
LGTsYbP4T8jnytNkDavStvobbZEed9PYsp076qB8Eu7D4YJ7gXfiztdUC6Nk38esLFwRjoywqg0T
sRG3KBzTyZqz8BoTNliSQDkr0R2q9Wv8DDlZDkT4pNwsOpRvBTUCLhohMmNG9gsxZ0h0zIxI5Kn8
9CFRCo5qMnfuDDq09DwZFQ36gWhACcfSA3Z9EkocxpM2ENmCKU9B64rV1lp2gMXGQLescifLpVy/
410u/h5HqLhwfNs0o9onecd5zxlPyHnta+yq3wJn4OLEZoLbGMbkkqM01oz5P4Dra/jT2+0NepCO
ghSEkWYKMRfg++1yIjh/NfA8pXzHMUCld3VuUkDI2wY+aZniMaYqJpNnoo2LQl6R7M8FQmaMVcDM
fN+wYCEHHP5AuC0lWYku8rfs5jFThb6iu14mIDceIjq8osq0YBaX+tku8KF2eTsS3Vv60Zif0g47
II0in2AkVLa3+Bs+Btg6ZqiZn6f9WmGw1xlzbyN3Kqx2GCU7DBoqcNKGCxlkDh57aryhSj86rfUz
i46q/zPzcfFcvSiqDeVk8VKSv21A9moPELIHT9MmfN74e3hxRqgXaeI3/8dORWs4BwfySvWBYFuu
DsUbi5la/+vtl1yhCIt3lyod+WWbF5hMwvAkJN8B26QLnS2AOCRX0Q/AGwyWk8SjsOs3bMQeyOYp
euaaUAvfySb92S15j9RNJU8vqF46OsQTv8y5wyCQh3uq9OvGaX4vHMHL3w/2aK26cE7EWS7qH+eM
xerUWDXJ7re3/ZSnZcJJoMbgNJqTlg5KzF+YbyA7+lXlUydLg9tcGpb0SWzD0cXWUhaVjrjybty8
2C866cZ30P1FvahVCoC31eZfgXsWzM9zX4PwO7FqMjXzOjofSOTw/86IXJ7nPVZt5oayeRgIKZpQ
y60FuxFNdOYBH3E7X/9il61xrIfitu2+2f8rmfz+qovkTw/g1HY/9BeLTsVNSA0/klVjLRlFnXJn
CEY1KNbcXALdWH/oMbBGtTut0HJBRE0d+QHqKvkckvcEBDxjCpjxXlcEWECugiK9lJkVNIBA4tbN
l8YGqYg3Igw6S+FuJzeL6vnf0ZlPrlIJ8gvqebxUetnJrEiLjFLPa1WJvG/JHGE5JlNd1uE/ySKN
eCBTUsmv3b7dbN8SgkzyJ8KNKoLv8V9xzlfLC7m/BCl87PgdFUNG62aJQQjJxvTTOnLxRTVZd8at
h5ZGgOW2yp7tMA0mqI11QfKdFkN04WU7d+9JUTfVlo+snzsm/9XN1+M/bDv2zLDLzG0sju/kXKuo
z0TQftVMrHrleQrZ6AQm3Tcjer30iHZAHYXhTfE5pTZPReJtfClZGPsNAuXYMov3LOsBqIXUfjdj
B4sgwZGmD3t9wH8Lwo+fsg7Zj/7OTNB4BiLh1ML1mpcvXygddRnguBurTpoja7W8nxWkO+hmwJyL
PhRMY6dI00+DuL394FS1f2pn4oe77u5xY8qE/zf/Jd/DfjzSt6Ib+/0WtcF4QsaKM9vWRU3pdz1+
W3dAnHLnX6hfcca4DOyeN8ybWLTumbqkgdFJvz5iNvWhjOB4KhodTuyEw2rLJIEGiuIE0R2MbmnU
c0bgv5iYVT1JnmZY5FY1YuZFTnQhoaAQdyui7fZNtlFudGrKSG/3GAKXWzDEQ6hYye/Oq9+AH4ji
bIYJ0j9wcXJBbDvjsF4U7FZQ631N4QIGl0m1HLD7KBsp9z9/1QjyYbf0izZ6rb3F5xbHfN3AOumN
O/oknVmDeg/Y7WuMnBKdgHTjB/lP9jrC9YGHcDM+xD2ZY0wP5szL2LWhFU8eAV1GPjdImag1TSvp
BiKg03BFCpJdwSVObInL32U4T13jXX/2MGYY+48COR8s5LK4VrLT91PoSX1XduVvpS9W2eHXbI/a
TwsA9Ng6fL7G+tU/1hm+YU7BHIhyC3AW0sHq9++PYjrOM7zuoba+uJf4zp+WDQ6oMXui47cQRDHy
f6vPVzAmSM0W1phJcA+A+gC/HynGNtzHDogCdw4wVsLehcDWbVrqLbkrTwqxHIEqnMZklYABjXLk
mr89mGSMyqAEudI1pFcEjaO3jWgwjAvQk68/qE9n6sHUbI7gPUNLwjuiIJnKC7/fZtn6sVgHvQuI
beg4TB6g8bj0zQGPJq6IONucBoWH3igiI/ATaZNN9y8fHbJ+sKLpIcnpJDKjXEAL66OuM8yEvNl4
YrKzx/li3E4kF/xvSkGpWM5tDnODfRuKVed7oQCm0kf65eHvoFD2JAuKnkufwxZDLlM2+WkZGnjG
oRiOL1Q2YfmAqPLZtheQdaH3AoAbefYIqMjbfND0GrOyXFQNQcG0C8nz1pM6HBo8dPImd6Q6hbw5
h1ZfZdGKoiOQvOoDQNV04M5h1qXiSm2oNQhMixa5hmEIuh1gKB+0mJmOg4byHDKb1B/V3OhhvNXa
c6qfOqA+7fyfDoVsaUY/lqAsPsreKWPvVAIZO6Kofo5rle89KmvTrjMRl58w5kdGULwvVP5N0eNZ
4nnixhlENiMpn6mrM8hvW1SrL2SXatTM0CcvNQKZSor0+Sn9Uq7dVGO6zSM8fIM4VOjnfGaKQaYW
m9EZYMGrplJbG0nwN9nQ3Kmd6PvUGNP+CCR+C2H7162Ko4OxoNXjVTZ8/WNHVIjRCQKwmxoB0xen
uBanheqZqh1ABEWmdNbm8SQCW2lKFxX79i6RAU2TtUePX1tjaTUiXVX3XzB6aD9GqP5Iv3oe2uWx
LJr++h26YBPTnt4txwfro00+ryPXjl8rS5Lef8dAVjzALtAWi17TGQouWj5DZ3b6Ue3YpG9KNDfY
Y49kWFpIfQ5lEUgj86XSTiSkcrCs9ZfTl1ancsH0UpayY54WArtppwFEuKXL8nF2x9V3UFXt9AhL
AUQOR+xzUm5lkaERUw64ij0u5SMPln4hPoxhKcZ/1TalW50CspypJF1oLQUhi8VS3HKIBmHpbnea
p4QsSLdUCKKc07JRN4hEj/zrPluixF76wyetWu092jH3GNhJkyKvHAUrlYbz5vVnjiQuxYQ2oSaw
rah//QWtbQOsnE5VMLWiU5PV5SfAWDeSca5AU7bAhZE4bEWHSr0SEexI5pjLS8q4OfSY3kQuAXx0
oPYhSCmuRdlnP35v/yCAYuGob6H/Ki4XXLYwTT94ixutSSoAI5mC+4lqFHFk5H4jDhnxc/hoZNj8
VgqIVr0+HYCMVrFLbTe5Gd0qd+IxzWS9jDzq4qJ/o7CmBctWDv5GdGb+tU+qIvO8TC4nGqk6nU8N
6m1o3iGz3zb2EJUanJMbzne7iFcNxMwGVcZYdjgcr8alFj6Jdw8cdbLq6//9f0IRl2oQ85fP3dR/
Y4XcRq7N6heBxoyVZxi3TYPsKjAmXdSFWNG9Q1wVrQG+f1xIl+5fmA0CvLNBq+WYt3Zstx9JqmY8
uSxOjUl60cEnrU3YfZzMF3YCDhCryqJ9MjXTedzc10MTpHA7tJDJXYoSyx3FqQf4KloYu+SQ9Zv9
Na/taqs+22eJOO9Yj6bliWnsyy3a2HIiNVjs1VfHpcphK/Tm2h17M4rwSkTEQvtYWNs+C3gOkdxm
xsVThIwptkVPI3CkQhWQlq0NkXwGPATL2f7b81yWuianmt2weVe+2M/A7YBqZe0PTzz2FF60F4gW
V9EXSHfTebOwFGcBTjHy+hz4aCLChFODOA8Kcv9msq33xOa2iXMz3cicuBXKRv+EQaivvwd2OSGj
wNaEIaYFubHtyDjQVeZZuRZTh8nZ01gKv5MkUpflhjys3Rqb9QDx4KejNcn/qCZPfp4AnD87IUkU
xq27CZ9kGL6LMyqEizxp9G3jMfE8R39h0ODHJZHiXwXNzMoZLLZprdgzovaJaxW+hHHalTPMBR8y
ps1XQMv+mkuP5YWqCUk4mTr2s5VcPUbtduQaMGhzFUFPcVMK0irLzP+U3IHKibuV2ZiQBJZHMNvG
TT4JksL7811BPEgaq+639HsseaTKacA940UCMCiUGSTLHjlYsVKkxlMQcHLq7q2Mvj8PJI7/D2ow
fGyKBuXUTMcEGUQfggZKLXwlm3V1gWBlKKdsdjsFFobZBZ1GL409s0lDimZ8i+XQ8aJuYrOFsCu1
MfJhGO4vVE/FkIaHm1EEHuKPjz1XhWoCUdLL6Mk7UjDxqym0Z0crEeJ67qCPmP6P4X0P1W8lbWQJ
yXt51LhgCZutnoDxCOwT8UaBkys6M9+3gfvLnSM/x3QeZlinROxBymcTfhKuXURq17dacWJ0CyVG
Tt4iT2Zzs1hEHyz935Bk/AsXQdSZzOnI6gRLj//Qaspl4uLImUjkD8ZznPJEfNSmu/SRhjZDcFjN
4VfOpmAakvVYzxihPdUzlDllkrlYMUDSvVDeOdjWFpyt10r/vdIIKxapz0Sp+nb2ymMLCp2AjhkZ
/lPL9iGVDuqySNF/TaC0vrB+qcMQjsET3o4sjMKbeteRLeDCmHcicLnXY1ga/LBP+lyUPSvTO8PC
LxhXs8C0hqNTsgAvb9Wy7M2lZlf8FYqFdpc82VcLR1xYSlOQfXAjIJ5Zjm6Vx4HRjl16IGxivS/w
460iCxtAgDBYfzumtjey0D+uBHoTDzovtZjI26i0UWYPZ74/anOYwHEwKRuzWb38cITwOZKjCuhM
7jn/ID8zcqPTpRHmSW3YPvRt3+nWNjXLcdaxwlSN/vXMLVL1MFMHWkMt5C2PFNv8tqbRTb5lb3Sh
XbO1nOQuKMizTH7/E4azehs/Wf6DaLI6SwJaE2MskpkJlN96dx939oi3FHd5xkZwzqb4SYVqGxkz
pYpm+v7dfAn9z8+YVpACUDBTLjXFC8JIPnNQdjIvuas+QY2I5PTlMqUfpr3rcMALMUwIZd3T2lXt
x696qnS0o9Y7dLQyWQSltmOF5oFbi2SXLDH3VwdftbHqqLu6UAWpNs2b4CgTLzXOkw1/zy05jP89
Q5Wbdihx4tpg8gg8PDCK2wuN9tU6leCZE8FOhl5rx7SNyLnIjLtgPhMHQYi15xF28TIOHZu1mWAn
MsUuGQ0HnjB/AVN8v+SQuG2y8vo222QAURisAX+oe/GQF7PJdu57MyFkGd6FT1G9lZywuSIr+dA/
8FSXAuBHtEiAtd/C4XxyDVlDBVSm45tCXNobwo6lV/pNwoEaLOZtY2gfFb9h/C3JBMlCx+mi+i/w
XdL1JXVaj3WsMJKMYQLSO2Iwg3dYZB6e0sdPrfgf7ok4yCLXl3T423pg9yy074+Os/PO1AthtlUR
49jUpFU7531wXzahXw3qiqgbHhKo5NxXmk70zUxiZYS1QP9exPrXJQJ9Gh5iKJ+nzfa/+KqKTeqD
R8xNTDtDX0dNwIGToeHzstYzTeAuTysHFzdQV0wr/ZmVqBbxCTdxtWRXLLsVmZvYVIdCIlVJ41N/
vC7jr9Z1g/zffXfTpULe1mm3cxhTQIYt9QBYtDlpSSxZXmu2u3T5Xaq8idSTi5sbGMX4TN9duHLb
B01xtVbnKqLrE8Khsdj5pJXaohrFcWhBHIvPF71FCGS6RsxwsxCw8pynY7eTvflPC76Jf0IXx09b
/e7KFpW73a7pcypp/RZBUWgYEMi51B9J0D+XvHFiaNZIED9frvg42KFoswI5da9rnpwqs6R3yLDq
yIc9gptYhhQ8WzWI8ohrTt6Ul4VfLZ5bDyzpYo/TfVy5c+lMbFzt2yHZKDklQH4EUlaLMv4sgXdG
BWz0VzSeyBdDi7aR0sSv81bVz2r/O6zYbKlRgcDBBIICWhVJRxJdXYC2o+18oa7lbx/6QFMVkzCt
oRx11xDETtDEx4ytvqFbQnPwGJ98ruZf8/HWrHxH5NY6O6UcV0vJc/UMr4/+JQQr+nRVHsu99RXj
TtAOmU1oxq1FXTt14Dq5jC6csJRXTHXEC3j03MPibKMVeiWPrmj3gnsNED6kdNoNkNgXtGLmcW2O
CaYxUhqw0AyVShvfEYJNrqW9ZGHn3mMhxY6cfxLj4V2cQAl0fzuDMJ/HOsfG/aVeU59krpdNMAm3
4Luj4Gc+hdEnzzTJd8OJNGNVkUM2AeajHNx4D4IaDvXW66w/WnRMdV56jgwOAEVWFwXZH4MN9l8g
qBERbNi7/Qb+y267bxIfF+Mc30tcAbtwL4nnjcZoIq7+u05ph8KbTQiQRRem13hLnMQYilbECVMF
c2VQJBrsf/SGxpUsnRV+Z2H8AyCNX58h1iY3Q9hLZEmFNnVpgrsDH1poxBmcOR/g4pMR4vmKEn/i
X6s83iPHOWgI+5FTKTEsJwDhr0Xfk1bR6WkNq6aFHeAnblvX3pZfKmHZEsLrBURWcWuqK43rrRMl
V9j3UARM588I2shRUbCjvhBtArk2NNmQmmpd4d7tv/qprF1N0YiQnmtzu7ViJ2UCrrbZTu9qzJ5g
mvzVbvui7M1T0Ac68QfGe+apCc5UpqXt1rSbVISih++qA3CUadSQxd0TqldZGf0ANhfUKVg14N3M
Icx+jmha+isxlvXUDw/TwND0tIxX87ijm2qs5FelxPTXZR3fZnNKkDFs+ZYYcIwfRm/URaIQtn+R
EKxdI5xI3KCE3BAkgMTNtS0139vx7zRVZqQulMhM+0ABpl/AXnTqoCysdXLlRzc9g0oAv5TTN5eh
y8BNS2iWexTmEdMABXPvKczBfTDtfHJLTBP+uAfYhHf5CEyqedKhQoeHXTIQkq+MQgg4d+OAxh3n
50MPqDR8Ek23uwZEBSt1oAT8L8ywRsuPAAnPw5DYGYUiTXG0+20d8F/oapGTL4yfDEIcXl3F4si5
kkkQXzFm+UrxAhWlYi5PSYh1BGg8KBNQt6bnBAUwN/3bSSbvSHwiOT3frz2TFzuLTbcfJpm6DsH9
sYxLnKVxTdT1SWRV1SfCwwAq76V1KEerhhEGfs9EzSgj1KXdLbjlGgu/KnwTIdsdrO5G9OyUp7iV
nk+z5nCkvO1BBiGtNFyDqeryQWpFvkH3eG+xxXyKvWjc9iGjh4HQXQQ/TmTOaWAOBiGpBugMMuGd
xvW5J54TF3SOALJUMIqOV2oGOjy0mWj9RZxL5InrgGaLJV4KXcMRVEYay/qhK5Cj/b5+e8MD4d0A
Bidp1ehgTgaXsr8VRwP8SEyf0BVv4EhtfiVRfn3heRTNQK4x+cZDO9YdJG1h3jpCyk88+HSMlnuI
hI4W5pizPsfpv82Kw5hhgCrAiUkUc5HCDj2jsw7EczmDQoJ270Xgx4e5ntwlPRed6bHSFXlJC6G5
fqfj9WQg6yV+9jJwsvF9y6BBf6qnvCqXUvSXbVDZ+4fun+ZcwC0wI2oQCzGciZAi49AbpkaRXLiL
XHkX0g1sOrDfnBN3GxZpFvej/IRLJ1onkyygy2ccwm0Oqp3l+38qIHFt4uOFUvASpivt8bHQw8aN
zEgDEJA7UxwsCiKx/7qObXt+dWH0ePYH91NazThwMekUp26ga5F/hmTRMByklqfis4TuQz8f6tUP
c8Wcb5bYQg1Wq9+SDYuzOJYn601MBFAcXXrJXKNotG5pDnp53fUiZhZZ3bOsfiXRUCLs7jxjXhQ8
6JQVPZXfN4m6A2ZXOFRm5NxYvVq03Bh0yXejZ8OepG8to7eWU89N7q4UM7J3j/W5jNCMt+q8+uVE
SWnct1EPSs5sly0PgkvTFFHLkTnLJpY+7jtDEU7nCPdqZNpelURoX4UXOvMN9bXxqmtPAxaqZnRW
E39xCNWrmjeSRhu+Ky79NGhcUA+/XhJBEufsgPSiFEMknc24I6ij9IxKLxArGAuy9o4jq6jVven2
fcGZtkyO3FbdmQxysWD0vWF9w0O5nCjhfTxKCTffx7AiwEaOneipZeK6hdTaA+mNkzvSAl72CWTJ
j8YJF24udGuHlZ62FGJwaWla/Y9WF9uvSWaHr5E71jZ0+mGb0yEHc5+nLwXGrSiqcUYrEtEWPJnC
TZcMaaZY5xf16C1VGnlU2eR4aLdP01RjFXcffPhG0r9ji8OQXUUjgrlOyBg8UpuTZetyhAlE6nhb
Fs/BrPuZVy2qQqcxzznEzLJqJt5RXAz8Bk70LsIk+mXStHLIt4KhV46DzD0Rc1MRdR7P9cFPAx76
3PF0Fdsbk+6MEj6t7gltO4ONdv2SZNu44mCyNp/MYC0wpCQQX5O2srAxt79yLC3xo/Tc8xg03Exy
BhdU898Ua1lellIwdlhJ9IWEE77+P7iZLYLk6eMOFgwVEVTKsFStRz3KAw5rf5A0LiyhnkRjnGgv
H1m0cyBK+JhbTxak9zjFnc/Po1H5K/xqsXazvPf8lAN1719OHbRw36VLYtBn0DI7PTkZgY1QkI/C
rf8PhnUmrLFknY5PCoiz1T0jSiDFFIHO0ZA6MoUUGN/kFj4UWC3EcDwd+uo7PfW8ajUKgSg7eHff
ddIyjWFJBMUu+D8N/2giGq2cZz2kR7iuGr/JbkKqeOevjQWdKnQSRt4+qz4ocIhemXltjDoJ6w14
CPROTNp+ZnMgmtKZoRuJPIfm0k2JcOIBF0HbWy5xHXmgs49oVQQyAfnYevdcBHwSdTv5ZW5XISoS
2yQcygoa7Ntv/odhl6Qm2Lxg+q2e9oSpoPJjQOWjhKTNpuo9SDnPR5L44BQ/Vt7+41EY5sUR8n8Z
hrcuPRWNGEvuXXePkOQcBwJP30N1XnsSxnDPu4Mzy14DIM2Ap7qYBkhnbYSBxgSvGC8WXM8hhQMA
0ELQB2mY1GxC2qQZIrqiWclinf4DGxDa9v5SJSSZnuiJ9Mkp6mVWhWpd5XeINWqcxvpqtHtZzs5i
inJllHa7Kuo+JfX595qDbONspo24v80ptwa6eI1b10NUirDgqf0tyekY/bjnr7VLV+ZnNl5mDHj3
HFvCYH3Hdv2ClyAqy6pxLOsKURhq+pfmrakbLt40Ip0R05vv/i0tucPkuEH/k6WhVCKzwyRAzdpS
CtHyFkV1bTAozK9Zc2h2GqgnQE72dibRCGmNp3SI+99gYnN16exDolqa6L0ZZ6oA65o2732R+WMv
SfAbDi4BEdi/hxzCEuzCQpUMihHD8OsMjgptw6ccGmnkNEPMqkBCH+JRq0F0ZHgII/FncXtfdQ6f
c9I5DkvKrLQci7SerlsSXfdAq4mF13ghdBpfGSbaX8bWXsGI4BhiOgncMMKqmyuAtPWI5V7h3/NW
1vgmeyFQapudqmb5Y62/dYOBexaWQ8EALuZiTSds/1BShNxsngBG20WvMlqaIVALPMryMEFiWjwp
2KAuyPPUWr/df9SNB+30NipZx1aOcqy0zKDVP40WnELRU39+5+NOThoCoh/lvhfbxRJcYDDTRKRe
wQgoj4kllg/h22QeAnLGo8F3HJCcAALzLwwBsvyIM4pyO31yvW1QeUaJJF1y3J3TQvKQiepeBjlM
vAZgEUw0nhqtSeqfApLczYlmmtbAaMgfXxKlEeYXQw7H3Dn+z82bgSysYMfUOrfZJksNr5URMT0r
mEx/FilsfBjv+5BGqYqFIcDwUt5R98LiQdMxkRe8KwlQ3Dn+FVx8TI/bpHo64pBEfG9dMNIiMUuv
JjZ9nTmODmaKEa31BVlHzYCNpnkRkDcACpR/VN8ERwaxJxwGpsTjmoegUCFlkuM9WLejg+73BPHv
sd/QUyxkHWhcl4TSck4QKGUhswWnOzW8j2+MkED4+LzXGXvtLe0au0tknZynC5GM/Wq/GQ7oTmA9
nBHb7x/RAFu6x3Kn5VysVbJjKGcBHHHE5QhFXGP+eY62jFY7E606b+L0RfB21tYe5+oLsnBfHKpx
ZRETSG/nDz+CaminFkRqYh/NVzt5kybQyS/Z6PalncE7XEC/UfT2LirSAOEuZf+WBufNlvUCKRzv
mcPXV+gaF/h6YiW0gbcWqnsxUiQEuNKNNbNG4gpaorE7hefi3c03TRAY+oLkZocSkGREFZW2rzGX
hyVmIUqnqKg77T02yv/m5UqTIXfB8emxqQ2mM4agS+o8pVyhTwXjL0CzLmpPKpWCTKubAqW8MEB5
huqtI1aFxglNUlPljlTjlazKXAsnXoiPFiA8aYR9vCRsSnl4vZr0JvdNAytetLC+WPbgT5v44O/+
XVAaakBnTcNE8Sv5NzUiuDAIuflhT2Kjhv4PpLCCqy+B2rdJomEmNQXqFMHkTRdF7FpJ/Oy6B1UP
t7AqpoMSQwS8lRbbNwQBVuUlvcUayWoZfQP3wfV8s1tTjC6hgaeKQ6WIG1HxgqI/71H3cnq8/CVQ
xRMzsIfKkXA7ogRC1itRnu+BqkeFoqDm8nQ9q1Uo4WifWu0cLFez2xmJA8o47hGrMAB0PowpFNu/
nNvafpjWov7h5CADq8H+SoNA8OFN4VNOVRqLlN5dBotfA3Fp5+cZdJTLMt8ctSWU9KOOTRyJ8wAl
A6Ei4fsZuHYnf+EpY/rXPvFVMa5i+GoKvJ0yPfJ6guOP0HJK2U3ObDU4VnKadAfZpY76YEv8ufal
VQC6M6P8Ky25agT9MSbSEnfPSxGipPouwpLIZCAmOpDSJotz9C24V/BuvRXFG7FhV3L22uo0uFIb
3wacFK9t2q81PxOILjZIOBiiEQmPaaRredVqUobdXT3tsZ3u24P0CGX5RCnrU6ZlLY5vrkdfSm9O
qFzJrlYAy2Z23QCe9GW8Q8harGSBRcL9nUN/vs8YAPcc4Yr4HbEoE/gg03uiSGhp5D2zE+obOG3E
bc21Fb+Ywgx8yplMqms5IWQ9c/dTmG12cpH7VtHiSC7gxU5uyVgNNJW6lngd6fWEi5j/9z/tYwvd
I7up7XKjJuQx6mjIKlgVlr5CUVZas70HBbMOvzqyCvJ0fXpF9HE9OwbkCJp5piwQuDeoLj5lIpvq
a2KoNY2n24GvKhypdvaCoFmsdlUC3wZjS2oY+o0i3sZX2DWcD5TppzpCdZoCTyCHnWJ5tU2J/yXG
pgUs/0SpmyeRZeItqSJcNt3RnheMQNyaF7peIKQ863KTxZqyjaA8pGoj7KozBSH5fMizpiQqCuPv
k0SWLkQTbu1DsUgFU/cwJw73w6puqnmZqeWS3dIJgNbD0wXt9OmNzUB0bbgjjGmbL4ENa4D+poj8
7URnsJV8FLghyWX+8JV4DvHzy7Ki6po9uuC6awm8bQbdaTVR1WOn9EjS0k6tITC89PioKzPj2OQ8
j2diTYhrFSzrTzHapCo5ICvunzRanC1+uKlXW4IAAyErY9SR4NwEttDFtxYgWcqEtzKi3NXWblog
Q4TIp7OB3ngTogpQUcIKun8+D9up8fUyXW+K4+OfjeAJPV+mD1cRBylmiaVesTIZffzghjscofEi
HiWDy9HXQq+NkUFvHGnxDafCXBHphUuRTdvxM9xT4iB0XjgIeed/w+cqYSip0O+mxH9DSTWT0bg1
i6L3sCi01aic/wf4SoxIOnGRAiVvTTOnU/q3HzykaOalEUkRM4hTE2i+xs1kAgnp0IVMEY+wt3pk
6ALE+BRHPkG872LOmdpRoc3SkfGkVZibxUjAOxVbyA7yvMuXsr55gXCtMxi9fSrQOR/CBhQRl7Kq
A6oRiaIVOXnRYQZCCZCCn3QlXmKz7Zol4QJEK2TDjsNuwT9yPxynv8HEWtnhP06UVDVSyIbbYOr6
xqDeN5rQZH99hVa8IKLk8KVG3xM71KVEIDcNiEYXjHHO4WNEZzDuLIx8MycJ4pFXtIcdT7HeMiIo
37h/JQypVDdB2IgjIZyPqO5HZmsVMxx52sLhVc5KGU9Js2IktSgPeJmdI4FI6UoEKGzJZ5f+7SR0
hwl8WvZnHUy4SIcsfFGVPvmRcpzhlY3NK/jlHiaVmmPtpA98oLqfnBjBksLNreIhExCoZeJarzoA
KCGIuJI5DhbDXBrWDTwRO9v9oFdpZSDaIHD2i82HVbGjHATA87f1TYHcVx5fec66GcxrMehnTZey
4zGY/W5LopnC9yhgAR8MVnq1HbU5wr4wWE/HIzqEIGDkqscoQn1fobRjGpLO22tA0VUOs2pppKjK
klD3mkbbQF9r5xOLAdP5kecqNtCS54T0gIFxNF7KdsEZWitSkmYWWLFPH+Cd4g8WxlHSB0Smttnp
dKP+GqAzCi9LQ0FjnRLubYmNLT18qi41JXV2BOOXrb+cqd02TP560B0/OECVWUKXiDvvWFRzpUn5
ufcPeDWiPLUBI0shxVUzl6vqJgYOxnHNZ4Pfqpl7iVjYe1rV3JptARL7H+dlXfVay8m6IRTvkqc8
p42hU0IsUYqSDW7/c9bjBuL2U6XCstDSaF2Ea0PFHCJ7T5tB1FnKR1d463nJyqkDDqkZiKXYnbBf
3MRVhBh6Nnwhfe/Astf0Z4fs0iK/c4P3liQy1PytWudIfIM9opGkQbXLOYDdSRi2zz2sksEhKeGJ
YsxVJR1NiE0vb+s2e4Rbob73kHl/9V/jJ4v59INNW68+e9h6PS6YDQLJrcQPYb5hxaJlRzBxO1yd
3JpO/ma82x6+fXTHUkvjQfAHfL/ohfZlUPs4ZeoRXP/4iUozhNuznlm7LC5cqAgnSr348YW3h8KN
lGh6eiLWwMDoTb6yMDI/4pUbRnWntzzf7Bugy+XQw4xu/qBOxc7lh66xztPCRV5OJVT0gEZjvjDB
rJZnPn+gdmV4wAoWIZcxuBcU/DmYB428Q/12LbCu7veLcIZ+E0RwqlpMYQ4mENfs7oOyV75XDiit
NeJECbpFE6TwkhMOmgto8vuV5dI7m007BNTWFRsRGl/KvUuvFuIcdYXUVACInL1TK1XVGgYpWqGh
l7actrZpQ6K64BW2M6SPewM8/xwA16/z5i6Pc6KgACWyyOuN7NHG6EbXZ4wTrK0CfcG6N61zwyLi
ab4Spx1L7xMA+rLtBQ8ybXKqh3ABmnJZeMwi/83d++ojRaOhX1lDejCfQGHSSRpVujDFiJCH7764
qX4Dgvd4FELc5dKRpTlHDX4/XEW2oWMPLEnANUFx827dNGOSyn4wE5pOAiMAvUWDUHU6sXnPn0G1
rxyAvRnwbSG1esKPUq2/y/v6Espe9OqtNOsr/Cb+82leQiHPeNf/dpK3rmyMfUwW11kkF/nXEALz
3cPKAG0nvqi4KkJY1H+zy4Fg2GHN9ianw+8ae+Lucp+Zx6ojFlYoMwa+5v048YN/PbGaw18II3xT
m8qRL7iraRxgYocXrWcJW3Z0VJTMwTIVXBq1rr8fN9BinLBEoomDMVTt2fpSYh17syO9khYSebDE
3Sn4RfgHxF+Yb26FLOOh7/Lbk8bgwgwff5LO4PolPXwpvwL8ROVY2UpM5vcptbwhxcnCUVKFuTZH
IFjBWVey6LOx01w881ZwsmJ5G1yjF7wo0qzr/MW87E+2ptvvy+bJsE8X8+/JVUtdkkuBm2UD0Bsz
cO5BuFTLNNWB9O8YUpTTQv0l0mmRSDd9cYwOqiqNVRj9yIqxNRpvBy6AcwTxG8kx7jNJ4XMKjBqm
IqqusYPH/t5ca7YRHn9kfU8CRuROQYIIJYJN9gnKRnWG1Ncq7MakZTxqiMnxVY5bD3KxuILjr5Pk
d5mlv+sBuNSdGpKhfb1YGwuKdym2caRPzvHjClFdhjgeq6icauBHCiXYMWSeTfYc5zbPPrbmMAe8
Fz+aNDjLj/Oq9bvPsesI9uWTdz5yfQ/nJOzJ1kDrLkoz3fMJNcau08I5rAD8IfQvv/DULPdWhr7W
q89u81Eq/n5Vt2QQu7YQ0FEeqqN2xqzLsG8ezlAUqpZScVhzRWKaAUvCul7daQUUn51KZe/3BCHs
atrKkuG/k0tSPLCa1Mv4WUlRAIO0jnZhmEjO705zr5rkoKCqb0LcXdP2/Zi3Ei7ad0IuVs2A9egL
J23nrO+32hBW+MjuO6/ESxrIj8yPTPg+0MmBd+lAHkd6MM7GCMiqdBgsjNm+/uNuDzpM9kAX52M4
Z8qv9VZve9uxljU9SJF4pe6f6/a6F7IM8Rx40tk+RV4nf+dlGQIVFIRvP5m8QoSBxzcrd5SfozDW
6xcL6ULHUAOHp1VdgovaxtFzsnBBPi6lm01oRdJuouEFiffKeCkyKBAqyrWCZGNgRgZPYHXTDN8/
7BeIDnEC2+0O+uyHtQBkTAS/3C5PtFAGXPBFLkas/S13XjpaUaask0bJfDAM/1sqn2w1lAPRuH0B
M5f/SUHFBlae6100ohynsTovu4IX9WKGMVRh5zZTGCWRYsIz1Qvqt1GU/5wCE7keIuOlPa4xQoqK
T2SBx0J9N69t0leI0k5jPoctVTRwW60haFk54Q7KXW23cLJTJ+pUXC4vDEzbnWpTp2W1Sii60tlY
EpnQ9hD9rkSpCljq5q4NUzSg960DiDfCSRYw7p4x50zItuq/HyBaKC6+LCP/e4ytFoetvxc3ODmz
OV5/KsA0BhfKIaX/9L4kLO2OzwEh17zL6NqVghDocUKsHinpYGvfA1coD42Gq2yU+AofUa9ZaC6o
RdPgVtoAYOcaki9QSv7ObICcBd1D7F8MUFkxJHvjjvYTcWL9rIYqnI6fpidst9yMq9onZfyK4G80
Koa3rxazp3PCEusY9EYbXN4bGXPVGfLKH4eDwoIQzWUh0FJJpuXwm2IFO8mEjC+iwNbjNvvfiujT
yxN23YxygJRlRQQhg3oiuwZdu+z2r0eE+8UFx0GOD+r1BfZWdz47BC08vJCqMJOvk1cSeyzqriqH
bT8Jgh4a/vR0HWnwyS203xEln3OQgZOH/evOexTyHkNB2/hVv76A4EYbBD7Lk7KJDl37xWvRJfr0
QNr/2DxOToSVERsiGLag8vHZZdrEYQtZZkFTxXzmjfu6Gk7gZHjHyvaw1srCVdB1ZBOCF+jMX1mc
01GSqWhFKWgDYL7GNB+mpCYM9Cf1aQ9ah1qUDPz+WWcUxNKXuyKEif40m4RkZc7y/7VUcICWz5+N
xAQUtqI+/Zoo97X5L0jR61V6bOKdLgE9tr7mCUo1HwTtsMQ2p1dxl+3R1d9bKTLOnnY+0qAU//Ex
MBdN8ek4jAybGbMyhku4eDGrAxRVtfSWSw74dEl1RXv6Bcp0Iq/j7YH2/OMhNLdEXCrBROlDed36
ojcxq7BFN0yOxddGxd9KqJUNgpz74o6fb2RkbAe3YO+nEVFUbs/QB2W+Z+/mu5kvLEnAVaG+KVxo
EmlRqZ2GFPBFtHpEQ55Mr7wwRzWbHOsLqR/c1AQYPKRt/zcjbu5TrKXOJI2JH2GQpfe1FHciSu+8
+pW7Ef2ybpdCQAnrjJkRMIhOJiKTzrHfgjh9cnabkTdDMg4mo5e4D+gFpSL6F1vVuNQ5LL0qY8Ti
qePgQodTPh4m0NmKv/YgMqqsbhluFx/z2eWFrEzK/gC9yu539uZDXO2wPbyugJvlvBrzsvCRnhSu
FDBVjEuOLBgYFtOyBy3nTfQl/LMGpu32u5qN798LDwrcEsgAVdsIHlvdm8Sy+qZ1tmW0IZ+gRwFB
k4ORmx/sZxsCFUJGig/P4akeshWSLFQdrZZ8en9k+JBmDxXkXGR8CLXRfmOADG4W0B16NlLrRnag
GSKJl6Ut9mmuVzyJ3Ll3IfSZtxViJJFMPVhPYCrCn6JvIaYlxC/eYlbdLlWPih9tgZPxAdKT3xUd
9H7LXeZsrF/kcdflWg7kDw8boMkCet8JDjybta9s/lQR52C9QakCKlcWjhj3sQBaWPHmbrKz9vFB
hNv/oeXT23O3UwvZNHoalcE4y9IzVqhz3NvKqKu8xotNsTXfDMYyg/lqTqZeUKw39NzvHaY7y3XC
+aGQZx2uLlVFzytvcOiMPbfhzJw2pqMybR5AF2aii1+rmKCJLJAWLQ0EePr+XocwJcvEZGq9GsrT
YvqpfRV8lq3UrtJtm/5K009kjj2dX5b8QSmchk0asXRq7VPGP6E7wpDMRYl13jZk2SD1cRkSH6f/
Xr2UliKqSHva8TEiAfyapqin8OLMh9S0YgtBZsdFYAb+Hvnpv0IHplbN+R1JtNM6Lv6AnKOdM3KE
fsxv+R2vxq4vwZUcU9k6gvtbEGSAlxBYsXL4Q1N+1J0GrPSwloe6CojRkYi+gOFP70p4Tsod0ZHI
eefS6FYYduN20TF/6Hj07tXHsitYYy4fq+Pwa4hEZYA+gcfEi/gIQbxY4pP6MxFc1UNPqgrEtIxv
sorwWiggBNu+OROOk8RGUIcdtUlsVEyojllGYC3lFWKhqEJeiWqsBbUzFN86uPdO/KbaqJJGYwoj
qseypcjg+7qJnNXUEAGA8idyVlsT8y04W5QBwJSOPNXdR3HKT+tNErPczljXZ+fbZFURtSzynL/z
4OyXpdvSevlr3oW0Yhup+0ETrSTXebAHLXZ6+2VE9NnZECunoCeE6LY1/3IQ9P99wXieLrQoz/WE
H50upSP+JuJKeWB0yNn0NIBxG1ERO77r/AP9wVcBa8Ad3556KshzC3jbIdFsp8e11ru3Mqobf0a7
JW+wh/nAvtj1m1dJd4p88MQpuMfpN5SjYjR9DaTT++5mv1egxnoqxdc0NiYOiBSLDODSxI7sAtJB
gHgoRa88wNTG5uDJ+hiRF221PWXoLQO6Wnsc7rwoL9Kq9hOaBlS0p9dnbJRN915b2+vZEVyGqcWX
Fsc6r/x6XV5Ax71Urxxg5H6pKlgdQ98ukmoOczV9unC3/K3Cthxazcu2ij/e9KPzaCSPHh6ObomW
6mrbnsqXvRuTGNvxs/q384nKEZokmfBDumd5PEklsLeC7eKXO1FrYPOCR9abjv+tyvxq35YtVbO+
Y7ED/WEUUb5pUETDhkZAnzVln6Sujz7Jy23R8Gm8rBsYvT1chNsO8g2d7NssdaV+96LoE5OdHB+5
enClNoirGjigNQU4y0lVKwk1tovz+OQhkImbg2nhalMI6OU3xjJGkrm5Kxo5qy6m+MXlhkDlySLT
PnhzDlnHJp9+aU018SFJOIWB0X2VIZdlm6MR7xbm/VUuVvsZvMzLlV77+OQH6+34dzGq9j59Yic2
C01MLcOkHWuKGhnNIFCBmmRzeuQeFIoiKxL8U8U+BF1fKH76/ioldLiAlBgF/3V3RnOz6Ht54IMp
AzRQoU33vthpdhzAHAkXYploqve5q6T3zE8zgeY1hBpHBhDrofGzy2pUD1wmcU4jyyYhgO4PVcMZ
bu9yPZjN3BzA0hsef/WpaIfiwNt1Aq6vBZ4NGrTsQOTsq4c3s+sVU8Zq7wauHNcV+rd95XLIXg2i
N3WTZ/On9LO1OmucbSu9foyJf4nH0OvZ2VqtjjI99U+jXNQQHf9+O2qiFj9DOXEtc9GlJQyt2sEq
NcvmYPm3CoKe0RaAdQlUfwzzsoX58Xn28700AOS3LDj1MI9qAdNlMxBDNekKzkym9O8T+jbePh5N
BUc84mWAKrSkaluaHzxLpSlXuPnpEzKMiY0AC9kIw1GAGOMcoRmEMZSYtzOAE+NFIMzjvJytpwdY
YwOKvIsUY165Z/ASBLB/WQ/cEKNYf3HaXXG9fxlio3490MwAekhSM7sgepF4d6To6wZVe1n1fBDv
yAZY4qD/22li8OtTdgkzOYWNyj5X1kvwAnCWB8vncqRSmeIYU3OiiDYGfdYj3JSgMzokts3Tt1Ny
DEb57Yw2bW37579TYb9E3joPJh/AK7DLhSgFvfRQ/eHgSEhEVfFwdY3GnwNYX5oQz60RODmVabay
MTWrH65qgOKsT55/Q2n2Cw5a7N4Xd8dyAbNiunY7shE1fC5wpdEsh6LMon0OMpgfc3j8HOrzzRHU
a1Va+pKydmoLkTe86HwUvY0k70epGF3V7hcEtpvPpp4/KJ2mMULkbcfAYgfj/ZAb8Ut/KSFvw7H2
nQ/Fj6RK0B8/tQyVoqhTqqCveOFUZjlZxMsD1UH5pagngoBxe5A6JE8agzgJGjwghFp51HOhhr0E
VJ550S3DQQzYedbwQNpxH8Q6qdXC8rRb526dGBEUkl4fOTNRDHbG7IJ+92kcuwbdCDUIV52dD09i
HIZ4eCVV2Ez1WHap/by3lq0SXP5l74m3ks+DNV/wcETv69QOJLylzqsK8fmdxqQSYr6MBNLUQalb
FFFzTDwclggvMQPqJ040TbXJsjjfywmKX1V5CaW9WdnhPpyW9dwzOLyKEYk1iFH7tSLLbC+7QDRY
Rc8LF1FkV6uz8zCRLxmPkuzF0TwbOMqIpyfOpnGU0xq7fZbPmPtduLoZ/PeYi5pfuMw1CCIZpcxP
ACzY7Bd1Wjtt8tFHz5UDZMHN02OF7WujLxe4+hf1jtk/abgfVyb7beMIEf55nXrvDtlRI9QFCZvj
+Qhmy7rcpAPLizV0rs65nltpfN+F13WwhIureYuw/zp/lI5ImtBKfdaMcrGJZwP0uobrekyBhnbW
TXpEfdrfxnhJiW1oI5WhtnVeduDbwfasITQVAhrFI2Kfb1IwGb0bgPcVW23zc4SjZkiStm2RyXYO
VKvQ7YHn27AflX/X8MqMif2jWUQvfWv4M63bVqc4vo1wWz2ganOf39l8LTPpdyRyl2bfAGyL2KUv
Av8ccoO6WVzBPe+63D+UlX+vTHCIBidXGrYghZ1UNe/eoDiJlESpXGUhQp4BEQxsPrLjQE1+2WUA
ijA02PQT3yyMGPszH1LkjvTHaU5XPSGkfcvAtfnqo7IcWi5cEm74VeTrUSxMEhVaniUNNCtnoTmg
EnrEjtwM28eyIBQJPHisokQLNT4uv+Zla2ci6BzpMnZHNKLbbKcqAbWE5gJSBvovnU2urEVB3UOa
lxhyOSDh2mOdAbiAX0Ru7C2QGFJIagR45oudjsm/s6If4FBCJKDMatHTK1pPPrwfPDJmqvvXRayR
AefHcPVFkZDokuqmKhotsonVN3Km08UqXNZKwinz95C972dXl1+fM4fJo4PS4eZpzFSHovi6mSyp
n3oWi0aI+fVzZJgoNM0TodRPmcdidR63MR35W0H/4GbakysVY1axvwTAmk0pp7D05ECDnUi+S0HJ
FeUKznzKkYcnuNRyMl27Wws1SlESOxG8AiyHbtswbaQbFB6KpPog25ojpPs9cp2r4ltFplBcbo0P
YqHXFMUkyFwF8ta7jQdvQ0Ym+uSqBwomRfRlq+kl2UqHioDjoUTCDUZiSK/cmjKAZ6pwvOzD+aWM
RINyBUgmuaIPLu+IN7htgVJSWrVHGzn5Usg9iCY1qZyc4G/NZWLlz+p3LDv/TeS9/nTfxwMlkdrJ
BIk6+R12uJixUNX1DMo5WZ+5Rt/DrjCkeiEprLpNJVA2sla3gdDS8WgtfvWsF4A83t9NMJfzjlYS
7sW+icIUy7Fn8qbYlU49Yu12UWnFATY4omyJ5CA2pyLLKl43ZndtDt3lLloucef56vE7GoMBbHQp
o0nqnkt9Hhzi2NLUa+C0wiokkclbwAZC+1D3+vjDO2sWIZNXm7qRldxhNuW2reqPq8qzgD1fekkU
WOGke/ZE6Qzsmddje+i5yiTsF5AnU2+NE6+Aejlt9hSAo6D/rsd+iYLdKi1daKIeELDKWYNiku+N
JEHjtVUJzY2cgRghx7dr0buszGc6E87J2+eZIFZ+KnSrdmdqOef+7b781ZaVaGhAKDGF3Ilam8eb
8feV+ygNopP1QLq8deClyGQdlCMpFSrMMP/BKYdjgK6h3SJStXXFVOsdf7JnVXlM2q1Aen/XA3ZN
8rU+4TxC6z66AWTFflRdaGJ0wHEzVZ/kB2Velj9lhpm4CmEYBdYBw/nnIraAPS8+LjsEk1fmWl5/
ID+zyIoybkkzo+plwLdbz6MHubWRKhXf4+MGF8NCdMqB2qrf4MvrAIme8xqluxuEDTjzoBk6kHcD
tNPlBGkjeECGITqhvzie64nTLmr36Hmpe7d5PpHxg8WnSn4TxbkNp0qxFbeu9JZK5J1ychKl0jPv
YEaqGx27U1cSNBl/KUffe7D6S7B/q3Y9VwfX4wjUw8Y7KODmVwDKw6xgQgE5j0kHK5e8tHXKSmrx
USzHqKQT44yNM26kQ8YqnHZSc9Eqe8K3SKCe8QeKEwmPxFFBUG0p0ZhOchHQ7ry8s/IrVTwtgDd5
zWgoEecvyiEuViSMGJig2Ke0vXz79VUDvx7RPBUaXn2sDsL8uKicKAL1BC+ABCkvFUQjhQoJlSax
XFJkWGW0Tlr1bCl0f14aXQytUtHTJ2gjvI3Wgts0BooK2hKoLjx/zC+cCKHR3DBxdEUDM2IlW5rJ
PtvgjM7F9RA1xbWJ5z4k4MbbJG75h1W42vTvvNC2JUK6iQ4X2VIBBsiIt30/SaUbtEgWU4ZnCfXv
WTQPXBi/1fWf37Lxbc6SitwY5xos2t2NhPYO0PRey5d3j3Dzxt/v9UY33gpxyP2A7BsN6ocV3Dtr
d40EGt1rQn1VjpLq+T2PQRWUc3Pbc4KfZVKMw0RxmcXNF59Y7aUetERyBRhp5mWE8KxnZhQGUzSp
HrGScN/i44n+iGDflXiHNPpjiTK80D5WIcwZLGDYD0Oguh+5/hG7OzGT1HY26cv3dxwUSS9CBEhc
fC4euM/r1LR/Nos0H+OfNXeqOLuYdeoPK8DbNHLYRTYIggMY5tRX+X9NFO26KMcrjwHelkG5OV9e
K79BrLA0hmXe0806FvbisSwkrnABY7P7/hKxsrSH2FgkeIQePFiblAb8C1Pv6tEsLqrJQ4UqH01/
yGymnC64s1xE+pfdJwzgc7IuOWIuG6BKpGpnsPLVjbrQFIHgOxBV90bGfyLosaN8pTC8PQpXYoIz
re2l8u6hK6VMLlCMbe7RYGuFt3lx/oJsMXHnS8WL9Bz+qIhc1+MFqxY7HygJ/g0OlP4PMzQx8RUA
RTVSIduZtEubhAVTAU+KR2SA2+Q/A8I2ASLhoDtpCDGio7HsMvH0OvzYLbaeIXx8WojEMpjb8zmG
RxzKbmW/StQAZnuA0XXxfSBcmItCGRDdGTpQHX3cbkra5zOWZ7/rzkAUfTGADSc+HoIw8Yi7YcZX
ug5XXU85lwkecfBs6URF1E/sxRaTzoELFLj8ZqzvHzX47tgAs34o8ATi1fOda9Ir/mU6mGz3Rysj
4B7TeRdP+65t8RB5Xe3r8bOWfseDi05x14DjG33rjO/vCS2tTZKAFeYLGlmT27yYgugOFa/EeYSY
v3+BaadKqw19Spal4ibLGqUHA6qL+uxkVZGn9cqJSdrDfjDT6gDI9dntflRKkXyIwKUepMzb6SyX
CXrz+fsPbperEX0xRZFIuWpNYlz7QjSpCIXTmiqpWYav4NGGp4kB2ffeX2KVx2dKuDDiMj1Nu003
17CihWhz6NNSFMxT4riX1H+DvDpEJunzUFXTaa07tk6VMmKCIfcCLdY75BsjUkkl2QocNcEnUw36
syVDxt8QMHSkxgesNY/6ZFB13Z0CW+5B5RyADO9F20Zri8rER5W/MkrxTmouXALbEkFlOIS+KxOs
IAEMS2miJjs8zZAxPGHE3I0Q73lGI6HRnRDa8WnxFFm6CpUw1SKojtzh2a5/oZzi0WbSlA5sOAZQ
kVYihOPDDjK4Rf+E4j8qQRB+58nBar7SCx/VpRxjadbyEKhVOMoa5HM+mKSVTzVjkd7c+bD4GqPz
A8k54GjQJstHdVXahsrTenNTE6+2jqfarVHvEgVL4koib55BkC8M6QPAMS5AY7EZuyu9HY8rAt4x
YhbIGnNadsuC4ElodOKCEeWjmLahokZe3W8+PXRvDdIITrbFLAut11wsUrNEOxdFyNXXxQSZZQ+g
BN/VlDJt9sKJTUZuHrt9kN35TmiKkw0IP9IMQCaTkXBvkJ31IlQ63BH5eq+nqATrxh7BieIOTHDU
6jvyfd7eHmZEmpNFP4saIXiE6Qr0ByLcFNuZnA7c8Lcyr+DhdCduSZUYcFLfjcQDkW2t8abfDzZy
9izC/rny8cU1J2BUZIpyRigjjj+GdcLgq6gDfoy0/V97NyvqXxrd5SKchRCWKbi6COSFQkbO2rHj
+dBJnVzxMR9o4m/gC+y80ZAlchqT02LV0MQzwm8O5k4ghlC23jzeVz7qxVefwIiKaf+B15jtJyHL
TyNox8lcwLNi4nE6/FUmB6swwi1Sdc7ufLrSy5YC66MWP2gEeX4ctLqPY+kbxsf160GqkVQD/n4u
VJhIYCUCgZYxWwhax0Az5y0+2f+g8jym5SHyvczOKUebqTux7yC7quqePZSPk5N4h2J0b5kQ6nbg
n8tyk1wSvgm1+BaMMGC5tFDBTf0WF8toS+9LkAcL7vuCmL3PTiw4NA1qwc4SwKCWQaAxx+24IPcc
51hOYQo8C9YM7v9fRmzr4d0rBUNphklybGWhjYYqQGbmD66h8Ad/Ra8MB22f3w88G9YR4NNmnUTk
yWEZ+0TFvET8Q0i5osSlpefB508nuP1sNo1l6W8N4KLi8dZlfiQ7JXYWvf56/KeW23N0qTyEDh3C
HwZ7UJRAW81w7THdYmMJ0gb6b3m6TCeDFeVVtIHeUiLoVBmqJDqEfOoDzBxVKifH0tAtsVchHhlf
OfBOFe9HAdjv7axcOC5ZW06cfIykP4jmAmvgbqtv+008aHa89oJ3NJdkWW7ItvD2VKErvpts11a7
Ly6zBxQ8AD+3O127awpPJsYfvzpQuyYq5eZ0Aj20ifVQ6poHQuh+zL5G3Jc1eZjnxXaITw8dVnNd
WjLG4qydCmzRxsqMPKlj3mWTcbCaUYAzxPRRHVHIJPLrTokzVx0jJWH3h2GVEaYa1ll8JIHeqS+R
FcTb04GHeBCzq5uLbrRzHbpzzP9xMOP1RM/5TM22KZDreylIfQJG78YSLi7sogIEJPZSmfhJ8Jq5
aWil82y5HZjgBjphgp8NUFcHfOGun19sppijWJPhpbPO4BndiZdD6YnMWOu0UndXRjqZt00O7J7J
V4WYCGzQy3pilC7ayshxNDZWy7mAuyAf+BdW7S6SJ3LXbRbFQrHZNPUn1ivfaSnCOo4D2GF9XUgA
f767O/l8nM9abpzQTPVeYm/z1SYzVX2ebdeU//rUtcSrlgtdygKQdJD6p3y2p5q2qU5n/TAW/eOZ
zIvhf02w3UHjaw4Dv8/5WnTecJyGjhngBsqIkq/HofZJum3wXL9sdBO9j3l/t4aU1ohdjhNgkRqU
2KcNlrGYFYwkzRiaWKcavBLW1NwNrrH4Ry0ZyokBe0glkdEYHAId/otl9nR4mJvLDAB/dl1uS6j+
GUHOcr98/4gMJq6flTXMMzCv7rbscO4EA2lLHoeiNT2LxEbZ6NjAMmsb3DrhrMhPnVv6KG7gJ8XJ
9NxHfTVVkIcscREg8yZJnaRd4QCXPnpgEIkDYfhA52v5UU2CJ1JFjIiSz1UvryalLO1saKNG1575
aP0cqOVFn/obi85EflD3aOqQ3x8CdZyfyOeOTJuCAEhL1iLMJSViN2zHDLdrMKK0OGRjTJ6nqIKw
1WEzXB0qCH1/3DOIXEPDBlWnICo02BVtGX4snh6lZLCrIlrA9+POW/USRLB2zOFfgJ+MQjdon+sY
Fa5R5p/coKM7y9mrmaJLSxM5i0O9EbSNnLosXZvlgyYD2z8tyg8nDIa1OXFDmCQEamknvdw4OgfE
ysIps0mf5JzOZ7o+/k1Ae+g1RVcr4qqar2Voa+4XNH7EBKGvdRBtO5R0L5DE+ufsSrUuJaEdFMtn
fl/XGCiTQDvKV3P0ssJ5jqto0ffFTZwg0+dhec3+fyQno9FL2FFTC1hPYYW1lAilYTOmzewG/0qw
fI3RqeDps4sHNLw0PmxTFW9So8r/7zHb+4O8tJeuDmn6lR3pjsdQ0HbzKKoqUKIEQbT4ZoViFmk2
ZvsVzjSx3+/wqU31x8Ct9GRNdDl/Un0c6RgLI/tHneG2irFw5wD6WJ/koRU035JumxA2Hladdar+
7ugLxWYA/I1BcqC1Wjlh+yYg2dOBAIs+RwqU1s24XTg093roKqrPAMFLaVr7mRK1xGUYwlXR8fHt
Ws44mdMoSUHmPnaJun0b9po73bvgIZnrotY33FqP/uy9qa+OkNPV8vaVa9Hq60kbo99D10P/To0K
+DT2k6+vEe6WIiXlDPxf72lX/vvcBACZ7g3IgkFkfFzNlGMXvEOjVHS8pXyceD1M7joXSRSnK3Eh
LOr5Hm8RkXYUT/eTyfl18Gid8JHgQLMSozKLqee+0qy428kVPaXaPl0jjQWvnAk+qJLBbKQfvRDG
yvXltJIhHhiuyiUTFTQqJsTOBDwf5lxrFEnSK1sUm8vtLvULZeTFfYOzDuC07fzT4NgSfyJ1TMdt
HCn11aIobHdxZf41CfWcOwipXQLMBbCk5+1mUEfn7yX5HUNsCaNGF5BakO7zDraHSn5ptPCwS+es
Vduterx3D+cVaSvOefEWhigoPkEjj04aCqESYUYZwxuVfalnz7CLNBE75s6IPUjjJpcg1voFJi+/
Yh8E2rIPHoN357KHnDMCj3lht1vojo0BKDCcHKebSpn88V4oGYOD2hYNpF2jt0Xai9R9RjucouEN
mxNw5uqttDxiKBnJ6P0zn29eoMkk9zC7mQXytIwZAoQXWlzQ4teqjQkMcXn3CJW8pZAQ/2XsUs4y
965R8xU3tZ5XqHxXX0KvkRcppg8bOHsMqit/ApUIGh8AqL95+At0C5XzMNCqYBl/ZPl8v1r1sv5s
b0bOgzrh3xm6eGD+vfXuOp1MbOdBa6Mx4vbIl6nBaOlhngrspCBGUahX+gQ5nzpc5xYva7EtZpo2
jyUqyrI9curaJgwkZ2ziwAkgWqCxWUYpuli7jHsJomutVBdu+wsyDfLMrWN+K57xf3KoXC/BzN2P
S1UtwSc9rAYFbjTOPIsclS1pL5lHvv+6HBxtpotyuFBJ6Q4fVgARfD/t0RweBxduNnM3mews0kMK
gRBLdafuqzJ4QtIFPvaAJkqfTLThxjCL/KKuUqJXY7pL/F77HYvtcmR6NLW+U4kMMlF3ZrFcx9i9
Ucm8+nztkOQIvrvoBsAUq29r8uNt3mostNvwVBUpQDBQ9xbRYaQCM9FZnoOKe26F0/yp76XLhX8T
yUA2JjdAEx0MSR8RUNJikIekb5yxaGHsI+g/MCBXxNPkbfOuDjpDVoOtXLKAu1R1sl96yWUBIeFI
FgKfkArz9XEgR5UF7kqZJCZTxYxRlLd8TB/nXt1F5AEUb+y9bZBNdzzQ6N/M/0MS/O6a55UlC7pp
iagL0Fmqzw5syAZBnK/TA3dkYVNaxaYer2u2lsZQm5PZuOOjQP1egUiw1SEW10uNM5eV3mxBSadE
NeLJD3sVfZUoh5UVp6eAp+Kq6rHO1FywCb8f0p15RItB1fVmrhSP/vYqgkS3pCs9kKpZDdoVKN64
XP/sEBZdw65c1Lgwc3yu99EC6HU2++cm5YJnSiAnTw54Sn2FRS56EygKb38rOhMQNjxRUZZDHHm+
Pg69AMw24hBhcJiN/CNZgff3jQ9kczHDqS8swBbFiI2MH14tUMAVkIb16krZ/japXy/b7PN0GhFQ
ZM9Q8eItODYecDG1R36PTweTg+L+EvR9eaVji4832Yy+3kgfVwEkGK9jmbBJ5+b9Tf0e8y7iRXUP
/SRu/tBzKps6N8Hj3RHUGwRrgSXdUxyIcgmGhfdcJXa28kKkG3NCXGyrir+uFFiQQngM7jpqrgR7
Wodn/GfyMHmItjvyApfJvO1YWPsrv6T5icRmWNO3CjfXxHPlsGucniRF0XGZ3L3ejPd99s40y+gu
4SiDInXaZpcxRVFjXB7JFnIjsrDxxnPVgW8vWcd2FD9fVNeNvGC8byZDcZlwlSroxIzC9a5ojIKv
fy/T++0NBJ8ur332euMVNNtS/+Z0Cy/bsDAf3cFTkY738Rp8HN/rcOIldKXX22XxYz7DOY40LfaQ
9OUFM6hJO02gBYliNT5cTKx76l9dzkgMv5hPQEIwYZAVf1yOz/ZArIpqDcjo3Xr4Sze2rBbaDMCq
av1RqsTiBcZfsC0QOz/fuSsIDJrtZpn7f+Tv8jvXCTk6ReOUpqAykRxMauermiWf+q8/yOelr0Xb
YPalUlOk5bXFRxWmWxXW9ZBCmFaS6SPpSbs+3q1LbVEdskXit+tB3B0pDO7tiN7DMP2UObSL6Wwn
flzwSN41jqBGJ5cwMO5/yy7fSIGxBoy7NZ6xky0bmYxj/HlrPN6aCOXWqHhxJjE9es1mYRAs188H
saaMpj5fE8u7KVSgdXvnYIewsYVTjWJkXHKRx6/UZyuiMQ+hOuBOSAOat37RxMsQVXnkWvKXD67P
TJTQ/jhuaxwd4xlzenVjCt46eQrTfXIQ+hPZGbAlc4VdkLZ6cHSJu+uxg1D78EMffk7g7TYaW8XR
tDvPO+WfZ70k1BPNSFqOf2LliiyxEP5Ai20M16WbMzdpX8nQxMYwT1CbSDw1eZt5AxMKgAETSG7/
SI/SwrdCmG2CNM1ifpz/owGF4v9Pb/rVWL5JI/Jjd6VvKuOnkkEaHnaxGdq9HS0MOoiU0wtZ8Iqa
6j0o59UjkY3JscjLaIjehAM0BwJON8sb2Gw13WtRtMy6Gv2d+PRLH+0WRkKfW0iZbObiCvNg98OI
Vm6VZSwL2xm3zAF7bbFhBRylYhQuSzQxMvry82b8hBXMV+ixSeGx1Xkwk1l/TatvhPE9S+xeEPlY
v06NbuX8FddfdSHY2nUDBxWjekSnqiCHNfrcrLc4mNJh0xz1H20UIFlZLWK1wYf8GEnfW4IfrkOr
diFfSMX3LL6SSS49FaHtuIhyeQusdnbtB5gxqm7Xlr180c+n4WIBviV4e8Au8698/oZRGxeIl2vw
TlxxhbnXdlNKoi7f605jdZvaDxtHgntGK1xcHibMbWupyekIbLyAkyvgVxksPKJt0x4N91zkyv/J
k2zt+CRRBFL/yPQoOiX3iLvPVMZnUK/8O6Bo38sCsLfbqgfdHLrxJCXz9kIM8qLS71ajnuIQecre
tGW4FYFBfbQilc8/kf+4ZN324Pahpt6MNAmsDeTs7kxNjWADXH24M3t7VIi1pZRZV6EddxMAeR0W
m4qak08yfr1APAdekroEi8GVp+uXbsXz6IQWbwhXmk3S7W8kla842/TL/SYgKcfzTsnGXPTyzyWI
Mahs8mrKFROJDAkkYSQi771ZaoQLtYcf8p51T3snmsJaDcGQrSQzdQio9kAKqSkdUx2H3KMuVBQv
ioZFyr1POIpf/jy7lrhTVw8b9hXhCdFMXYZHWxftY/YmAUBy/UWyKyeLVwG4/1cCsQfhxHVf07W/
lsAfDq0zPjZ+ABC3QmN1KErlGBS1GhDx5CzpdXOd9jQfvIM55uliwYMYPwHCPahvLd1kRVYngRfY
2Ag+bxWfD5XfRUlQeQmLsa2iE80inKPRS81e0vJF3lOMtFD9GjRcBDqp3K5H67ziFG94iSb5hgdt
ptJRmnFMbTzjC6BoP57GoL90D4sQldYRisT0h2br8Z2QuSlZaw+Y2IGHo0MgKmmB0vez74HLhRtQ
A5uDIhHUuMKaQlJGyFy08E5Y9FE/SdkxOXdk/3BmFkdGhNcQF2bUBzf0IHNX+ekCEyzAWQVy5PhS
Wv5FMih9+wb3p+MiGGTWW0T7DFHhWYge/V9fkAvfnHVqfrE/9Z5tfpBAAqu3PkITgoPZ4eEOWKTz
rUZVxven9pMzilX+7ea0CUBojlKMz8M4mB+bxXEBtY6vcxiWzjLswH1fpi/66RcP2gDtNR5egd+u
OUMjijrjUSwIKqB3A1YgnGniZRjBxMLSLbZ1rR+xQkUmmySaJX0EbPeyri8NDHTctyS8Qqt3slBm
F3r40lyKiHq+7Xdu7C5+syOCWC19/PL2eFMlR8k4MbL/7dij+q115l4tnUocEtoBEGu7sFaBClHi
NlZtm+1NzgxZnHsCFvUgvWV62VxhJx5N/7cVl2JerJ1OYNlZ6KkQVbGfqq5CFU2R18iin12UOJR9
j/Lxxc8VbatnfQBi+ETi85uHPP1aEqsFHnQrpd2AoCgHCA027fYzMrASlIfSgvpZ0GGRXvcKWy5b
/HLE9IslqiQ40JR+7nSPG4vFfVMfLvs8w40HItopGnABPcFeqrz/m7X33pZOTq8W0vVb3v2FiWMe
CQfmQQ3JKZz/ElaAplbBTbYMR9/GMjdquvxPknc9fuUHoaGACeEc2fRV3O5zUTSm/aR88jRuxugC
b9ePNYzFDGWOlEfsC0y7o7Hl+u6DCX3MjzIOFIcOWskccUM3oCgXwj1j0Hq4Pzjrb0OsS+cmzRQx
L+sFUAhUvVES70XwgZQPqsOmb/yuJJwBBQngJGIEzkHm2g/0ChiGIYpQkN+3EM1rfvwzJJvdLUw6
A2IQfbJsGWdUDw4QCujmofkKKcdcwlYr8KuBbvRQRMQUM41cNO5RZUoZIBqYy/HRrXX0uHUOj+zg
o8VGjmkOEpbS1BxjjD1OifmtFXiitWWrYct8qiU1u7gjdMxTbr5Zxx7FecvV7trLbnEzIO8Dq1hm
AdYDs+R+QOEpzWoqKCti5Hz4cymOd8Sy9yLWV6EkzqcN3KlPAHZLyfna+vBDq+QQm/21IXFgcDGN
Lgp+LBx3DvjPsaE7LeE0YwOBYk/vi4/dj+P9CVgfB57StY3BiiqYdq/oTwcltPaZoKEeA6Ip5gpJ
YX4P45gvgWmTWgupMhzVMxa3Dn8Jb28MM4sXG9f+/yY3CEWy4VAlpyVlCWrPRPCcoSMuzaubUAfs
/S5yvOfNEJKZVff9+6orFQLbkU2pMCcZhjFTyTAT0j+dXC5S3ta0OgCYRjy9KkRFEpH86LgVGbvP
yMkqWphKRqUfKSrpBWpNw3wXzmyPNJ40JQdQ9gnzDsC0r/lsp1DGYhzg3R9gnYoF/2AVSFnl7Vwe
p/8op+A7Kxhr6P0FJPQ368hON3VHaQKSz0IV52OiI8O96EdapyVhkOu0uOc0Ovt7DXSMzCQVH5kN
hjB4qgwMgO1aFe8lPmgVAkfNnYlI7dl/tWL2F06NzmXjDsc5WEVq5q1wmbgpPCtb5tj8pLwCz1uN
9++j5fHA2xLs8oYmNO5lChXQxo/HnBy9ZdVUVJ7rvSO7vIcj5uAsIL6+SmXONfaEV7lTxTFwD618
frBapYWkf2n5lnyPAQcYVQlbO1BD8nFot4P0rLfXUo9sAuPsqoRAiS0vJpeOFK3Q0ItqCKq+UM6r
k8DlwsyEoJeCr+1vxpry5VlqzxM/E2bPEAv+oe5WbYUXZszjWT3SUdap8F7Kl+VbIZ4TTgPAxDq1
KsUK8sj4ARaw9xGNdPIjqE8SJzTChvPTKXBUsTL7NuHoYW6lgK1X8LjxUhOEplCiX38f/VEOh67g
sDwrzZb0RDJVSSgzyQk5QzhnzRJA3tJrNGPx8H1HA/pre3I0JIMFXm0g37bHX0FKMnJWrGt0z2N4
4Gp3q3Nvq0eYn2L6pCPdgVvUXs7DzjxOPJuURRyJLCVBFDDnVaRtJ/rRwhLt/1MhMN+sA7wXiDN+
nWK+r8d6gXUStGtAe64Ah/zHn9WbtyzZnuB5IGtWVIg4+upTjy30jPf9bkbHtkffSOAlf464d+J3
gIdbF8xdVUcUVMnU+ZcZcUNMzpv3o0BwNM1KoDaxFqyeKrcWxxRIWXJdBGbHOP8KsGwoVxhsWFKR
egbonvA+3RGmF9rKCujH8MShvCz5eAxxpLE6cfOPWoPCxhcEcFHif4mu9sNq6PcMoKjplMlZTMoL
BJgeJqMo0q76AGGXhHqf8cQFuZbVlsAFRx/m20+gbt6Di1bF4zVp7FPQcdVRqrv/YYRJ/iqWIRTi
Xq3/65LAAHGwnQrM8phR2U3GuUMt0Dvbdz2Xx2rgxLsjqvlGzGI3pI2BD5uOaNlOyMbWFBwx1qLn
sbmarfToH1tyGtNc/Ns+G1SSHV3NXGtkGJfnI0LFErURcOOT5WTr73fTJ+Rp6ne0CyHu7GlGIaUm
ur1TT5xEloFyPx22+X2k/PBF1XhnOMtzMh91fYS8tva+jRCiKb0QetDtqVqjdwy5Dy9sNrW3xqEi
6zrBI2ax2tmbpRSp5n6Ve2F6dMN3iCB+gjU8K5f6+vSWKnpOYg0bkzcTJsurtC45mt0/iidqOcJU
NvcUdzCpzVnvsrS7mIu5lJJ7QTnJWYCLLqLuixGIHhBDeQdfNQ/0/Yb2uAiuOdVuzxpk3aEaBZ7P
hs4/6tVvZVe8FkL2Wb7KGYpmLZ5A0IaQoOZiNuiCCP6HVEV4BOHPbjL8qg5ht/sPrcZYmpYAk11T
cVVYuW1hUx4oBwwcLUE7fNwy5vRysCUb6HGEyMx/Lj4/T9LEx/NXTQUFUgUQSW0vCl6uweoPl96O
6flL3L7+uhe4/aZWCV7VxhoykVX8z40bCBIYEf1MrBqXNyTAdh/6h0ROquTX5q1MwdrMsvLtulev
d7GbZwODoaCpnRYlRfmrLVenZo9lNcb2fPivumJQyLwxTZBIP5wFzu5Bzll8wcZMI8BulLkgne0k
/SyaUhfjGgX7UMa7KUR99QWEd8knPt1sEEe++83pmApwmmFMJ5l594aApwyv6kOwAOQ6nlKqq9bD
5ZzsMW2YH+bCZUIR6bR8JRwnwZWAvrW0BXdvv4lgYbhahuk2mHisk+BbwryLZddvp2RHWCKD7KPB
reTa4qifs627aohL68iQ7KsXSDgt5+3HHVM896XdoKqCfC6ZWASfK/yPtqUr/mIAnNusD7RmNdmV
8270cRUs93Lb7ht88n7tuFJuFPQ0C1aDNOgHkgm+qPlg5hDd2CoLxh+OOdUHX2joeH0JtIke6nRD
acANfEFN9TaK9pLvABwihbNpqvuVYjofsuGYTNAsKACs8G/Un4ilVjcANlAWAivezQTmlpnYs6hD
JUzY0CfySyeYcXlzpYBkaHQGGxVQQCqM0JsazOA4i3GoH7onUJkypOfQkqZzuZVNQyj+i0DRFu13
Elo23+dMI+LL73KAGaa9qCFP15/Qp240FMsdS3kZzmGk+vP27rTQyqzMIUeIDyrAIUHcVJuTBSFr
SpPqOwtdJJ2NtG/ErN13rfQzzEGtGy4+vLz5/SYSG+xZKR0713o+TlOIXU/rsKZBFVp+kHaU5+eY
/jr99yfVfaf/ukPPIdvJqeYTQE5BC53hGMhoNdNQfhDw54eAtAjFOATMIdCd3UeYDPjOoCNosMdT
e2NdqFOga4yhB1Hfs0TDmAKHfOV2Zbwj/1nZRtX2vlfvuRjri511ff27L/LMC7bcBSsuobWMzDru
hqngUNYdI38ZWCzIOirEUF/5pLkUeFv11ms80wW+usOkLj6iYZ9ZJ94PtvN5JevoafDZrwLBdqZW
67qL9zBwoBxbXtHUByf8F+pxWowr/vXf1sn/H4lVTcbDmzyvwbyt75eUgVUABL8tJu/SF02/WzaT
41y82KUd9waH775C9l0a54Eqnz2Fr5K7Pu0A19RyLaBWK7cbRfzKlqD3p1KKYc7wH5rc4UyCtqya
bHzbsOr/fPRK5xBVYPyYvhqyrhHluyX+QZqafKIDR7fBT6rz5e8t0J8pa5B3iob1BSOWg4yv3Ufs
Sn/xWD2S2IUTMA4r/vIRzU+A63meXuXPusBZprll+rBrSy1/4sx9sJ4AhF7eljybrPCahFw/vUy/
dVpI8QYMRjGYBXTPLwKbtjXIE3nGZF5Oxuotco9k7yuwr4bijgaFbz6MdXy47PVr2NFHTMfTcnwE
wEeX5RcMavUwlzcroPSRh1mADym2wJZqYnWvb2aRcvTYEouYupPngzFTmo77LaWeELlhq1aTauvm
h5+Mea7NSwRxjHZ6Zxpug0Mif0c25HZMUDhCWF4zNLvA+dl6yykzCEPMuG8qBVe0KxHfGs8/u6D6
bZ5nuUjgzS9p7QWLEaakfCZqJLitnz2mF/YPtA7J5sH2x97/DRw1cbvV0nR+z/i08lZhdCdPATtT
pSUsOmvhn758NRYE086nldAWc20nBlrxt8Sujk0CH8ZJRgP/UScdtkJ2G5rY26gJ1o54pI7dgLkA
CIPg3DUv2vNRuum/8DuSwny5igoBgNBBKeFfo/BjJ83DViP2pbcNkSff/FrtH3tNVJip0HyIiJTq
KIrser7p99tcTAmsFhZ7pi7gn+IG/xZywLwTx6dtIZAdQih7UYOYyxtrWjEIOXGfaoDQDvRuPIxa
vmDCGrXpVHkYvkZC6DJbF+sVam11fPBahK4IP89VFbUjpvjAsROdtZHgre8olBpv6J1f0JxSPLgD
/r3YMm7hk6i4Eox/7+5BI93RzABVy/TwIDFjISdQrZ2y0zkOww5Ex9AdqSURtEBp4gvp8XHJjfzJ
fDGeh7Ezfgaw77O9ytRU5Nyn9fzhT0Rw5cvOFuzfMSkhSgUmUV+6zXn23JYbmwFt1VDPt7EozkUt
2GUY9E7CfOpS5S+/8itrmM/0RIUyHxMla1kV0fxYk0ByXcwV2woZ/5JBOVfD5HpnIpHChp0icWp4
DAEHBOi9ArOgqpn/k/gTjIh3eeh1iCCQMxmEyxUr0639eqzF+HT83gK0RQhZb9gZlYe0IALmgytC
HpOLRqqhERnOMcN8S80TR9BA9EUCloE+/xv9NWgHgOFhGtKYqfp5n3JgHZj4nBcUajzYntLky7fD
jci60zbRpm4XZN2vxMFacswntU6cqsY6Wy1ypulwDlsM56zWvmme9nCCXPpS2NY/qjPdc/XenfAY
R1mPBKONzwyh0W11+3cAgwk+G656xPw4zcF5G9qs+xdIwZUSLUcKJfTiEpQk14aDvLs7TjQm7rCa
XHI2L67O85jXxfNdTVU1Vo3KXBo6uaGPOz6rzQHT+4rDfzvqsuqSe1jINqwZcyyz4k2PrxXSI6Ty
6Iltapaf3InSfo7EtuEElYte03mD+quW9BILYk6vO3Th4EebR8d0hRTqkRpy9lmDPr8UYL/G74iQ
4aulfcb4Z5N0FgnqP+M4sefpoxS9be4L3LZb4/YbFNEn1TK+y7S3ssXtLSPOyiCRz9d6wAoG9ozB
4GQVeJfJIwkwnr6vwu1MVZrHk59lW4esOsvSz7WjHNaXsvJT4KVTy4wgldziyfqqzXzojHzzlNPg
vsV3f3mG9uY4ln+9Rhs12H65lgFJfNCwSepn9JrRwRTIIsvFGAhuY83jXvCEoCxNSmiUs+E5bBW1
lbJgTfBo6drfvJgQ6oITdhVbTK5n/VNW8F2Zh0edQ0pALVxJhqoq2momB36T4wofWg1DO693LxAz
EeqXpqyIblpI7jsaqMPh9JvLQWwasl2QR9PXWuE0KqR4TW0uVQFLCb1ysqhhycbhA3Coc322GWum
Asphm/p8DjJQkrtXO538jHMtW3OTubCD5w6eVmq6B/yndOQ5kMotPlCqgUCnuWsRor/z8uwcsgSH
sUHZnykBRIf6iaKIcz/s/sK4SuN78Gar1W9Tu6ZjCfWXw4/1DT3sZWhcyC6fEG4gw4P6Rj4x2zxE
D6TjFRsqx9RKLyK1j8Lw06yqnHSKa+ajGD4gwmWr5fsJkA0vJ9w2edmmlMEi52ByqQFwBOkkqzTj
01kubEA2/UfViq8UjU+YTkZ26oDxFfALjjDjhskdPfEx/PbbBeETNEHsiPxbxyN8z9wzmUr1tACa
9nwf/g/puwodsGHROi1NM0GUjp5I8NAbDDm8GiqWq3z/C+/NEij1JCLrpcJ3HGE07jc4eLhR0e8S
HAN8n+3SK84RsKpUweOsN7p9SuM+U6HZWWRqT0KIRBAnl4OPNJFb33BEvv8Rzkp90cGU30+yuBd7
IpPFIMVf7Cd36zrbuh2sV2Jqv1OYmiymFB9qxDTVUI4MlKpCovx4iToIwAjPSL9nMqfWB3eLqfT5
QycDNsRl9iMZAX14wJJqKwvpqnO7hO5L2tvVIaSOqtpYjVIQL0ckBhBB3qDI10Iws0NRK3aoJgl4
GGpQtE0lFDwRtbom0WpFhtJlDAq7/f3yVxH3pUqzSI+H8FagEwMpdXJfmWLJRaY7rSb4dYdgdrOv
t4gI6JtzLHqLJVEaon0KY6BK1FaecdAKQkgMTkBq1sGRqQRDqNbYy4YZP9MbhCtQr5VXcj6yu3CM
XGKVQ4grZ4YGbco1xtthLAZxiisgVhnqRO2YcHDeBXG96l3PftO0OVEZwEF0KeqbMNHPtM5vHKpd
oN5lePcaRLxSLvrPcefIZIEaf+jG2mSAvZx4dznTmWlBPuMG1oRv427bBzPkOx+sJfwme/DgOX0N
m+bTc+tyyuDuSZ9+Jy0voq11fISTusEOaFu0ulWLZfoXq7Vs4w4AxdYL06m9lIAfP697UVQbHWTF
RCbh6pp6wtUA4sW1YoYUaUKWHDRT0EdDrrJFpJakHNpI5eYeU3CPNzrWTt6S3hd6jHWmbPHj1f+R
FzuRypswW+zBrCtoYVfhFwCrzxPE2+mZM//oK/7CFHcrK+oPoAyrLQvBaRNax8aUG5ws5Cxespcx
iJJImDDE81BW0gU+nKbC4yizWWMIFWqpXhIL3WrE38iJmKICY3+tToVsGFOwMIScDfikZeYmctg7
xTXe1xRISkOLYgmXYAtnHZXzvtmpt60Hf3tNVpW7zvwv54BOuGAfBA9ht6om29f45vjxfCdrJ/bT
bjG52lLSl8yVRcMSYpB9nR9D4nLAMyecSG4iFM83hjKhWGa7VLO9GCFNbwSkY64lA5/ksn5JNfQp
Ohb9tngRwBJbLMFyHjIidHbP/0BlFHsM52Y9OG3HLKGqUVEsn5mwDdl+FA5x9u7Y4w6QDwW5ceS6
N7glkksD+X4BK6Q/lWbUG9eXqdc2BIVXoGW7O4XErxhToNkLJK+spnsyHE26IIMSOYiU0ClIjKTi
cFoXZeAwIgLW4xeJeQVUPAWIhl9+G3+32StkZ8FfoROsrXUg5GgVtk6jw/qwXDFiXlkfA7sYxERD
VRL5QKCSWYgKo9Plv0OSGlx6o/QeLicZGnO1yo9ohUW29I4yHisf/ClC540R2yH1JNL7ZSbtOEEu
W6Yg+XiYQUxNZJdxCtYIqB//GG3VzAfuZ4gih+WXXnXYSRM2PWH0SFAA+EBUxcbGV69qwsKCevvD
Vk71ZIfjgJ6o1ecsSao0tO3uxjq5ewfrgcdOX2hL9tWFJ+NbdoJmx66WZTds15PH85hdRgReVwb3
EBI1iAZc9BbtpPfaxCQ//ryKT/y3P77Ttj8vnEPeECEMeDbalA6fX03u+36ZJZUy+X/jB79m+AxR
iM6MI/UvtSDcC/fMN7IuAIH6kwyFrcXxUPeyZTTFrKkgjGCiJphbCX0Gy0KaSBAv1nd3gzjvAVsZ
f0fsN1x/PEmAdxF7G6dEKxWWEtmDpf0WAzHsfIhzJ9UcX5HrBhj7Nkl5iys3aXoR1oVwy3x8LGZc
P31YNMXnAfHNdzgryJWHNIBjuabXKgjKGJUCIlaU0ckEZHrnte056tOAwLXiVCYghpumfJP10LbZ
m6+OCzm1Cthmvecq+A1lTWpDL03lV1LHn9OOycqFNvarFcTdHHw7OU2f4ctlb2Jy74WnxzvVXrx2
kyIQqnV6ceHccW8FsuSo6sCo4zLA4oxkW0eFx9h6VWp3MW5EDIu6P+cGtFRYApExqGcdO+NOLhMU
jf+7EO/n+FafuM9KySpIVshzBLnrOWCpz0Ldm/CYUwxWTvosXXUONuWbLYroL3MtfU4mQ93xQwyK
gdpYOxe9uLH4Knp6pl3767pvq5ojSaIjO7JTqZlx4uGt/HdLiNcomqZ0D2S4Eb/abeyIKHN8yfPf
xqR9CfyE+h/aodDdMPq0ibOEvkAeHfXyR1IgJO5NhbOBx9VnmX9QRYTvLnw7ENF96hvQ/wiBgWyi
5Gf6/YLZMlMYJXxSFq/NGNCstYYgZAxOgwigTcNP/JiKGQYlLNphZ1snLhPGP/ayny/0xa1Q3BE8
+OutoXVi1q2HhBDrezvZyNv7wVjTzIJdQGDy95D0aMIt9KIVOGJvsxfmbPy141hQxUF8VVgrG/cc
LFZ8JqqWDxbHho3dxZ91V4vHlZdVspAiTkftp/q9sblU3M/+7v5/DiH9LZgeQqaS+SrDWimDre6N
34XBJ7ggxngMnfAQARqfolVkPT2fX09CGuw+tk8MNfgHPBBVILreP89dJh73VOu7+ImNCCw3QHen
VpXMKe9p/f2YKszcCkC0B1YhK9Fcal4wr5bwPRIpdJnUth6/XKGUlg+V+yY43qaZPbMkfGqNUWH2
3O15z3AXZbapmXEFh3MPookHuAGzet2szsxh8oh8p615LtfYgIi8h/mF0fbEhS7BMZNIRPoc0iRO
L8xmFzXG7pdeTvuze5CaQyc2LU7EjJx0KJqLO3ST3muweNLDiGvM0ckuqpSHm6VOCZlZpjKVoXoS
8FgPtfqkxnW9Y24CuyJwLNnFOw/R0t5VJNV1tuF0ssDiBV8Nsu2mK5czSlnyNF2Z3BygO8WvpwNj
nkBYrMhM1qAmqoZ2cxMrYR/oRiFiyiaUxTvypu93uI9fmt18BijrIDH+Y8g0nN2zl1vYK9a0eBfn
h5dC7p8Z5xSuE0vYJEHEmP801qAfJLIGexzBgKgTOg/zD1QLImH0+iXkuwwu6NcyjpgUh9nNTd7a
Ah6zzxA6ouPRTjwwZ1SM6KypDSFexxSUNHJ2gKG70V+Ma8cMHx/nhb5sKakrXgtO9rEZ8hVC/3+x
MA+UZqPCrL9lPcp+2xTW/K8V6o/Hw26OXv9jrNRdAoO3+G7VbIt7ZLLh9qQMVBGpn2kvN4Qzyh8z
vjbLDB4dla4HRm02odauzBa2RDooZHdPCRu0jZ4l4GuxjlYVkEsfHDbYyy1iTxxz02+bla2ffoDk
CXZwbnQbFNpSWH7vbmnTj6OQX1LsYr2K1xjLu2V32QGxBtZ7zWWtYifx3jiHcwtdJF/f4PfVDt8Y
w2v/DIYaVklfMmc8o4mpVidk3zJxk9bAQc8ssawtXLTS6LPWlsDvcCNufbb0Mnq8Hq48V2o1u2MG
AP+2M7Pi7v7Yjt5ROzD4fBK4qhcEzqh+IdygwLLS/PEmX3I1uplJlGTipaqVe9HciiJc+eq05xfh
oFW/uwEtuAWKTL03P1Z4MgzphaghxjoHA8TCLm7Zy9+SBZOWAjS5w24aDnVHwXlRjm10vkhWeTxQ
X6fEwTk88pTGSNeQ1W43JjgklMlIO55eFAL5QLx6FxqwYNzh5x7avs9MsLe9N01SWNai3NdEi2u/
Pcy68KUf5zwlBCGJ0+8cYXaQet0R6bGXDfxLzWzRv4Lt+G+Zl8o+s5tQvaU0wYo1SKYqkxg2l1M5
m9/JFgFY4+/ua+5CWXOq+Plu3piu3JqeNnMzS1OYf1SP8xuHKorvcwK1XHGsijMZbjfHiHm1IaGU
ORWiJDJZu2Kz+g/rHtkSggc3E/Y2LZL+5LvnYrdeShxMftA8s3E5hjxWisWLwIY3m2HXL0rxBVpJ
dsz6T5qLUosf5JgKA0aN8J1LDXTmfSI6lVRVGIfq8yx7YXvB5E1dP1J1za/VkBDfxcUEYZ+uonVA
3GD5rpjn8znNj5NSgqTw786BcJgZncYJ2DgQ6L3YEashZwOMyMNBicUSzcgPzK+Hx0RM0hxyFs2F
E72AeF3ezjTrTiZru1yiuMbe9bvlz2+AwZMV4Sc+lnnUrJEG4sPTxPtBkil7hZogwyslVxwjPuHc
3x0D2MLvN8sA11IBX//4Pj0LTviZNToAvE5cjMzPO8LVRq6GbJOtijbibICGqIZDr928H7IDvhZZ
0OTV4tu657/POb5MT6PPhT4SxgezOwqecXhMRR/OBJUDEGrVTABoVH6F2VU1ENIsKRw9z6Vqchy1
rHSkTG1RP8AKakYLeoIFR6AZaqmXuEjoSD2v5lsvVRch+eEbRVnxcbKnIt8iVpCfE5A6Y+PScc7b
dUGIRiREAois3mTE5II5df8LNpDfaRxADTk8Vm8yRw0/I2ML7Mw3QqWU1/yL+4Na3Ciyba2TfF08
iUsuPQZM+iaYsaHLVdFaFpmx5ziwFJOdLBIcTzz4BoPMZdbgRgW19KNU4fiWXaYeseBzfpLXn2s3
58Oa/MdKfN4KGPH3AoXRsau9K6ud3wHNFXBMcuOd9cORJejWRUzhm+BV4mczhUW4lj6VpUWUAjm6
aOU+1HOjHSsqTIQBvWRSueK2mX+Q+fXVvxFiVcuRwcS9uimmMKJTOSvqtkxi9jDZLSIQZGVIKxDc
/cxQNqCoUFqFJlUQpwsl76fiYoSPrxoiS0errg3/yWqPV5l4lY6ao13xQ3/gTWP6se75G4zHOJ0V
vdNWE+vWF361lZsNApmOEaYqHpqHGpz1Mf5TCaIRSnD7onOzNd6GVW4NoSwUWTefbftPeQX3UuGU
iy7r6TRumjqu0QO4LIjOjPKGkkc/63C4k6PzuiQ54yXn153Fk5pVfT+35y54fbFfeAje4vuBltYH
U6P8J4AOgx74PrVqH2a7EGsC3qrBVdvPWh9d3GATgMfHEVt6DHce1QRYsLYKXyMXrbQPu77f87Qh
ShPRSzEnHwofwzZWXU47rl2NjhEL5Wm/2p4ELC3281Fm/33LhdF0H6jW/jNbGzxUjpZWvb+cO6kB
LE/ayDCnC1a7v7zsYxNr4JBEYgw6mGa2U8zfTRc4xvSpcSn8fHcJyWtK+kQkZ+5MLQTs0R8L5Fb7
PEOie3vBfvyvHufdtEVNdajrIUMdLK8gFhKezuGIOuSRcUiQzSfgRWM+qenwZARYTBMGol7qilI6
t+95/ImvMh65G8smr7KYOTo/rFyhQMrS/OxAN7BQqndGcVWF+Ziq/VcbGGNJRdE54Rw7LX2H1qWb
54nrTWfPkQ50Eu1P2JJSDIsJ5X01kedBv69ooyIgA/D4GZxCgFqhEf2gbdz0qDXLvLa2koGKh+E1
IsiJ5PFxMjImWBgjSzP4OUhj44tJoLFyoWN9FC2a79jg0S7KSJx7Cy+0fXS3JNDIcFX8ZYxnPrdz
0Jzgf1jAGPpGVSUrO9G7IhptqQVbwmwbXt19fcE6eFrHeTdR1JjK1EtayRKdN0Xd988lD50MLyBI
K5qYFuNYVX4H/pHdfc1cEjwilyl63TIcvRc+5eXPkgrQ2E5+ZYtjkgpcqIa14BNMLwrDoy4o1sEk
ywn8rAho+Esqmd1k1Fc6F0TXokLutOiR2popLDhVLqvzPe1jqZNi5ASl4N15SppTbi+GpBS+uyh3
dWFh+2vRrE2I4yEU5jchq6yAGRahROWVRH7NJB9tUvIhyb+6DLi6/OxCN11yIx52gOlIq77cSPM0
L0e0duMgBJrR3OZPxqeWaUYyrGSdKwo4jt08sxWe8of72wcz5cAZdGYdhVEvIQipeke90GtBvMYO
xJGiEkzXvBAfvq+Zf52EA9aMibLdB9wpuiEXJdEOG195fH3SQ+7ARQ52lyPTYeLKfftJr+Q6gmQJ
eRK3ARnAX/+ZyRDblekTowEqI6QGjO76WzFD1vf5/5eFee5lWzgd4IqZSCvzx7ha+sIiLPU5UhuT
QG2BMMv+SPiG5y4XNRTai78u7gTU/hctQffrZhN8OPVYrf2+rc7/VvBuhyYegPyIvwDPlLwrxTfA
WXk/mqG/0AT2gafrawPO6KAx6ZMyW6Y9U6M2Haec5xkH7b3/a9vS26WC3080bOnCmrmiT2WNyqJR
WqB/Wp7YUTDm7LBYQqwIdilNznbe6XTvYmOeMPJlC2CvimP9yCXELCpwaOYclTDrH6tlybTcAo9W
yHdSaGx6QSXMI42wIJASqaFds6nKA/RTn0v5an65IaILI0H/fV4LylBMlm7AkCzV466wNUPEgSaa
Nxf22qtocdaXLuPabz2IOu5dND3OC8TvQ9RHPPhD4EOQSfWukoNFMEU6B7H79ya7MZndyxra6y3D
D5xK2geyD3VaW7nFLi0FzBBtdJX3gFb5cFrJJ7hLWyegD3C+WQhuvc26VxRi7t1yRZMVHHsTKV65
gr7e0Q7Ze25wIJJVsQFgRkdkuVNrmeCmrabxtPp9Xn2lzguePsrh37vlalMqLdUiJ1hdj2ZyX91F
J0fxaIZ/OfkzrOcl/n8DW5ZgHSUzYF1/ALhcbuIcQuSbch6pxmez1xqQ0AR3szSOtaoH+2AyUtms
BoXSnNv49kxlQxexBZbkmUST29DFmE2QnGs4rNgAx2do2fdhQE0ClCd50DhtbqCuNfxBHRLNaKfY
f0sThulB7R3PUnX1fXqfLCcGOS+hksOF76iUNYiVIX2C0FHHEDuRd4d+lonf2TCmSZi+MQbJQZb/
QMkBfph9SrKWDWti0qz/CpjoOY7FIcbtCMnpW/IAjczM+VpH4AsfBWRwROugJj1eZj7eVs8z2azi
IdU0FOHe2Enp9498vZxqEPhgz48sEcfkuoZACFsSVSID5AgpLTKtatmVsassssvwpunUqvInLwrK
YI5hOlLXmjxCtFFkXzUeBtz0DtyKsI4vSTBxXCRoNIbve0nzF1aZ08vMRkfsvHpdW5DxxAwC24CE
+jtZ1ji62egTfguPnDlnIIbf/2R4Wzi1yXzKWHXoK7JIPBA1L1vIF0r48PORmdT3HssOYTaoZMKy
QKHVu6ClGOt0xe7vZ8dYaUm/0nSUrxYow1Cgx9Pnoh+fhbuKQr4NKDe7CEqBcoUZISN0dLPU+xf3
RWtf6BcmwGwG/6RtotWPiekaZc/7V3LOxnKLAawd3r26Uho+zmXmSpUYzm4148PIoPAHBREedUHr
TqLLqbbTasO2F4fzi9yo60OfrW+TTI5zuXNMastt2qzNMNhzVsIThRSzy0zlJrTdZ6fU0YHYJQX/
iAbuFtJYDG07SXkrXNKJLHIKF8lURakUPfhLQZJXMzqOtLfF1UImx0RDtZx3zS6AEaRsu3NMdTED
4OekiysEopDK/WGnCLVKM8zsFicke4STqa6FMYb+aYkMugkb/N/0RA5Zyv1L+8qWbJf8BWluL4vR
CByNNpXIdxW3oPo7tMCsFZErbQkEbq8YIn4mqI7r/5x00YIZpKI7mfAjWiKWLa33EzzyZ3kGhqTj
0qTY0f0GYmQEYd0jhc1FNITmyBkAiPfFWLa5Br4h2qUoRTk3hbixwVPvPzxYNilYhkUWi4sJyPS0
Hczkxn2C4iYSHX5x+sc6aSGQ4tjsBdOx+bFx7AZj42CYde96SqM+60x0puz8XB1lbebohBtIQiou
SkQ3bJXx9jlH0s/wDkUvJylqR+V+vf3q6Mzf6Zu3nssPZEtHECbUSD9WTRf/il/Kh4LPl69Y5dEf
jSoDaEfruMz32foh3Q38u4wfdux73rw8H5RdFYARJgeyqK8RcbRGDuXSlmCeAPYNOHVcUET0hfqW
zxNwDRfEvsY5CD0cBGFogRWSc1ht9501Rj75O6TVmNFgwfNwl6ts8PCCDz+j9YzzqFTc71zUoSi3
RzkHaao7beGW7ThCtvqav2lJgkWBrF3QLQn1nwdnaMtDZpkmYT7F16tU4/by1J+fryA60S/Jwv5K
4bDD4EhyYtCipeWKHlBEELMa50PvHFVopUe7eZQdcEnWRab8FhO+VqCdxoFcHRMADS2ClFKYVkGy
kZq5uT3dEURWzD93iQdPVf/QVTMpcTsvsWFq/derZ4PMk0/qGJ5wGgIU5tRNcFca/rVZsiM0AxPw
+z/h7UdMgv2/EQpGjz4Yh/DybE6hG83AxIfCfe2YzSGVJGTozu1H1oAjGdHDeOgAiU5xucHb1nwi
LlpNJSjcGj2NvQ3KhmuK9uMQzWbM9JsBL9292TQ4tj4yyexjqb7ZtVTHCgHqWStc8IYsgGiEVibg
5PaHqr6C2TB+BEgu/Iwm/tElwPRT/Fy7LzJCdJSPu1wi82MnuaOG/ziSi6aeerN2fkGYQq7XaYKG
0oug6quuTeWaoHpf9LfevOtEzMS1KGAxgfzvL1nQLvmR4Jjs/NvFLfG79nctRxGlJh2XjdKisIik
rCeHbEGvBxEhLH1IhYEEbJCws0P328wLOEXB4FDpnkVGpRuxnCs8wU2baCEyb9vlc7R86y84OdO2
yawJkeVcI1rAnnHMEBohKDQLnUTW5QCpr4PjPoZAez9sWQ83Po0YO/utedQIjwklytLuk+qGkYkV
mgv2IME4VKP97IanEsYf7IWP2I5QhIhpbda2OSqnw9K0RgVzyHI6JlCcqPwke3iqaV30Bj3nnMeV
e0Ho6/deoBXxF4q5unrAaSzFEiGqrWGaO+U/lz7Cosf3lzsER8q4mPkZ/axG3sycZ25GMrw/5B8f
dfVDCmpF27YkGMdtC++PA3xlrZYqlga4RVcnAQAvGNyN7OgGpEkjFb8irtbrwd9dsQAIrl0dwvsv
gTe0R7Cr7/dm3wum5egUK10tvxAntF0KVUUYwXWZu869f2PtzrDBfpmU6O5ASNrveweCQR2bUMPK
Y8KcXUEiwVFIpmx88wf/LJSP5PrDzUNSFugA+ISy2IlLsF71wfMMgdvGwo+Bnbx7Xjn+K1G1OXsQ
jSQwNKV1jSk9JMvMYvAAbmGNVx1O0gLfvML7a8sTp7W/Ud7FqZk6vEMBiH8+Aa+EGpRqRj3YP1ZY
NM3gDZARlv6VvXvKY1Xd5shOb75tdXAiUIDiTgjwSzdh7Ln4bFBGAm2tVKvaexlA9YZ6ErFhTRUv
F4rJv7ITqkyG9KVjE82KFGNBtUIpHO5ngbPHcy66PLvtn0p8pywJ90K1fuvEqmiGva9iV0uRrV3E
3zNHBojOIo7ltswag3l78j1ArbGWPDMWUHw9WsPPwgRaABgUXIyCSOy4CeOWVL8VgDIEc1MrdRfD
pP0mX6lJYtHqv18hHIX12mVt7s1qenMa2o7yL53sPkSaWQZz/Q669/LE61065iJc4tHD2IdBD9xi
fnTwWfcAxayPYXhqehx70usQJ7QFlSyggWjqxac62aLYolFjcmiYQeF7FOCyUUgJpmHYQSgPHrr7
MB3F9oa3QHJ3QcMDAAYPW90EINqN/3dl3WF53t7MPeLzzGLYFnLtccdZlCh7+80by/NgsIutgMJL
ndXWkWzd6OXC6uQXLXgeAvbU6+OqXqtiVIgUdDyaZHHCz87s4JefXQ4PjdTyeST6+EWzfa3JOVzw
IsG8n/niLqOQv0XaGO+l/zCEv8MYFxUWG7C+JsRzn4zT8DtZ4TMc0P1mw2bOFRMuv0OK+pC0Wvz2
1ztpBmybymOAOg49o3Gx9A9YH4Ps5L8/UdVUU07oN7N19lRzrj0aen9lcwLRMwIwewwHk/D1p+io
K8FhYktApoCSnU4YX+h9RVsk58eKyChVTJvQvCypindtnjFls8tK25MaPX/DL2V6cHbdLnlFiWKW
Nmn9JsPLXtsPHM0OKDGdTwUKamHEmWviBEWQZ9okIGUM/YrBq+P13Aqsq1jRZO+Gn8LkH1oMRXvO
/mLfzLongzgFkbb+werlBJ4eHjkegEz09BNOY8t3uqgeVP1M2IMNc1qZRkr1fwCkb6VQWpKf4H54
u2kyYv5cUx5F+A/8NaWO8gmp4TNDgqWO4i1rUvjGCKqMIaDVG1EO2J4o+i9GOnTWcN8X7YkfwVGp
1V/bP1w6+4J5gBCae8nub+MIWKQZQXnsWXDI5vUcvi/EeLC2JId39sK/37J8NrqGaWUzqhQ4naRg
NzYuRv5Xj7pJltM/KjXLtlZAOfCU0wU0mlHhxuFyhCBL1biNtPbs4zhcdDOSkgOzRBsnh40lDYMx
JM06/jqp/r7zaGTMA8H62ruaqK+FmfaI1abf70qNWnn++6FoWPDyLeuzB5sQcA4gb9dgh25DtxZa
V0+kTt+xKh4g551VJ/9BFhWvc/HqSc++ERLeHk95/ctbn2eWm/vGgjgg3epw1p8FTRq2PlRkml5z
k+Tc+d6GQRsRThYmHm9+CGRGMAj2HKA33a9keuTOAGJLRlgooHPf8BpFsN6VtE0+eP1tMyz8ENEh
nh05/7DpK9uXkCSexribrZidU2sqECwrUNe2b8hCcAX4aa5q7zk5CVhxbI0tKQlUuC+PYENDZI+Q
6WdEcisF4AErCDMeWuIlUWtfkn1CF42r6zYhyQtyZIUZmlVRY2O3lc1CcfEBtFfdkSfYmDIrfG49
TRtfioYVPgBCQNKbFpyfsHxc1LcIcuXSi7UEU9y5RErHBQRMsabLiQtDj/vcjzKS1po1XF6yOoBk
c/pEmLPncDhZxTvskUbFggizkDD/9q3jje1sWjSbnCQHZbeucox73+H1wayax7J3QXLlUQXXFxO+
yDgw5MESt76G2+uM2RGJ8d+MDKBzfeTsxuQPKvZmX+MJCM+UWgGcewNjIG+G2EeckCiEOi/AbMPx
1KnAwNv9IM1m2eMPwywfkka4vWQElxwjvOoSCfSLFMNFDAWpCOhCynGAO1wI9+VMu517/DEtuy3g
XXXE84d7hqpgtQ6ifFW7EWUt1du4oDK7SKvxqKv8vqv+Gy1G+/D660GkEF7Xcv6lF07d+UmpZYMv
mM2AuO5+YGBETfx8j16cVjPKzgNnT7wegLCmkUDGCzHlARpkjiHctXSNO2OBjyhsVx97AOpjw5fy
FteClO719TK77om87CE8K4tgxZoA8yoJVI1k0oD16zcoke46Fe90v0u2BQOkkd0cHeeMtQqSFTKj
H3GmvrzmXeUfjxBvRuC8LDsCi1W1rARQaGEDoSy8zJjQlgHyP7Q0NP4jepXtdojPt70uIuHvxezm
r+KkBK2pLLBsBXWBrG2qP78tfcs0Akjd+ZtwHdoDpryj+4PggzwI0bcQt4dGuLtOcCieRD5kF062
mfRCHA7fYqYLeliW/KnlyKiW77vCqZHuo9r3ogm+lj6dQDF+tQqOOG1oBsVwaGxCmz3mfDPGoEFo
zU1CqR0yJtK3CgGiejJgDx7MEO93JSN678t8H+sjw1rWTOHLuaybOOd2JGcDeAuic8eAXQJo3adO
b4r8jQrbFzTe2vvUNnQ8cP3u+2M3dJJKLdnOkuV1UM55eOOtX01bbBEJro5EF2WKf5yFsCa6xcLK
Zc+dDyBEXme7RC30dRUjiWC/Ju/h8oeh547sHmC93ou2aqYjmKUVY0tiGfxb0xFLsUoj+mDIX0Nz
G7hm2aPZoSwTCJWXhSY1jNkgJ1ZD9L3gvnGhWpMDi63j0HLHweGt9xZOeWpkZBXZgpuoHJ85d6X3
IDZzL6vZeQdE5175UQEJmjIo582oj7n9OhiwkI0607KiUNnHsm7Rh+2qpGyW7tNwyM6k5djAzQqJ
5bXgUsnWQN2VGlhu5FwPTfKr0bk+EAnFA7N+mlw3z4XpMb73xvbPqzKMWA7AtcQflbdipFriDgAn
sxuzOdAKMgGsVd78jUArka4WUriI6Pi/atNVCTDlFz/04KsraRIkwEji+PhfMvSN2GVj8/yM3zLA
DphRlfQP0P8YdeJ1er40ohssuHPWexJKCsNcS1QTXW3dUG5v7NA8Mq796Z0Y0ISAsJUIxNB8r84G
uqBt3FJ234FclZW1ltgKPxECsZCAF3V9rBeLgBhgRlDABUJ8hOW6DATRPmbOH/QgP4LSRaf1Nxz/
ZoxrH7o8c8S+/riZSbyBI6p9FgWzsZXD34egPwxr0tU2k3tYEbB2TDUzSQI4d109O0p+UHZiWqBa
Y639uaQWvnkY0/hIN4UwkI1blPdse27w24JKD0k3s2uRm+R3D3bLZC7MeDo88sBZzTfPKHCWoG2s
sEfdJVxPuTOC0CqzTNBSYr1KfT+fl7XipqfbP9IDnANt3gnR+HTGe7iQPAD8xr528fh0iBZEIEJk
31xSsiyjp/ZEUcV9oPU9ZnAKKWlGUN1DqZxun9LvO3nZ4+yXMKXUThiS/xx/D925MeJzMC7pjdVR
k+umHqIMwI2guF1QSG256YfiHpRJoD7Mvfyu2fqIdwf3bC7MKlXLW98eiessNYEUamHvS1omlUp8
asKY/FORP8iSmDkWKiW6xDm7tvhjtoK1bGbZM02RC9I3bmWJaiTrJ9v20ud3Q0yA+PQb6RczPd4k
WxRoVGzRzStNI15Er7eF9os/Ny7bl6NwTTZwmMDjXFUwTlT9LsudWU7cZEPTBuXXPrfjKAh6l/TL
8xPQz7MkTykYiKdho6lSCiy+rbuS6rynx9j0cb2e+5J86vaDTZa66eko11IGyE10WPBcKfvfF75A
t0LmhYZCWDNJM1CM9+cq27AhCkrldLer6gCbUn/m2T/sTEfdmYx3XryjF3B8XrPQgD5aypOPTpU4
tlp9wPnvPkMG7ctW3T/ihqySS6Sn3GbaTKd//mUtMUpkcUilmfkHu0nj8+rI/Fmn4rQvefwnp4x5
LOC3Dtp82cvjSlnbYcO0ATNSade3cUiXDvHWOTB4OfJGHEc6Gt7uEfz+SwFdmt9LCCZMrL0WJiem
pMqI3xLrd4DjglnVGZ7bhQPKrZEjP79yUJwIYVnWEBA1zwYg1TJqObgOv6Zn04f55Q0b5RARr6T/
aHNKwsc9ZJ0koEHENSJAyb96boAG9K6sblUdIn3Z0yEOHSJBFGYGDGdwZa9y9PVT6r9AZ6IFPwrC
yxtg4nGvNgV4YWP3vfZ+3FKCzex3ZTPDPe+pWb1+VxKbtvlT65dI8zU4dL0oUTlZEo7G30EZufNR
utgvVUXPjCb7/2koLyhwxA+zQ1qRPOIKRxk9r7RV0KPZ3eIXqgSUxKVmv6lTqpXc3ofzcbxB7s5S
Mm2csAS63jWv7tAR69x6J6PC5APeYtFJUnuacVih0uSBCtjKg++xKR9KItVJ5FsS4tujh5wj5xni
YR0p+0Fp6AwHqAx8ouOCe4vuZKvqdzVO1yFMv+USJDzSc3zl24ZG018iU3Tmr1VvfkvpbJ8x1SDf
Xtr1/CMC3RWMJ84J7Hj+4LOOJJeL4yMDJZKwulJ3tlD59S08HYUAGUbVxCQSJ75Y2SWkJYiLj6yM
hodyQ5/82qZ16hXXH+ASg9nS/DascI7gH2YJWMGeD7Rhe0domM1/OzvGUfxw0XA0Dx47lyr0HFcL
5DrQoUQwVw3A2Gju2Y962/XFCuhMt6A4nnr4GBJLM/hFgWk39MIfXMzQ8USoGgebvl4nJgpMezwh
PmhAW4teaQNKsG/n3W/0Q4yYO6+BGhm1fhgIUHE3ag/tK2jPAvlSrNm10fYUGU8IqP78ss1ffBKt
EzjdRJ8fQvhgZZEOTopeiJpZ7t0AqHCihFUY0Ab43vZnnpXIxlWkjJQcLw2MltaNvqeJQab0X08e
Aae2LHxaT6GiPiAKbNDEafPRrAyQgyau9+re2bqiTSw6uwHLbSYFZ+2fK7Nqwa4UgLYJx8E3BE41
dpYb/xPDyjmO6mogiIsr8qcTohESd2KIGRc9HeNy9N9JqG7O8ZVYEyulbKlqndiHn+17OyeaaxMN
Z9IjOoclV5PcVbhJjM8B7lbI5ohClFcxnrWWuJUYOmaS6RHzHCIcT+4YEysKU5UBEhTxXVw4DBWw
SFjZo6n5090EqyIbI3nMLOtm5y3KFVRAllqrpxSSpsUmCihOL6PsuUtUfd+h0umJAx78zPVWkLW7
pgd7CCuHc5H27arRt85tFy7xtO0BUZkxHcTQGas81qv3rX/pG/5CkIv8WeMCV5EjcxKgoIVlcVI5
w7sKtOOUKFwrVXktWmXxY3kfzPkfOQlv4xdGyfJ3C3jkDfxgPPFzmvmO7SZCXMpoJb2PPD4ebx6d
WP1/V6Ds6nNuwo+p0AIGQ+r1qmcrhQ/KSXTiZQXozRc0oae7Hux/M6JbcV8ZN15yVLFD/EQwAE0L
ugqo3dj2v4B/6tyErVJjU+Pp3rvuDT3IX1eGOpPJrfiPKIBIWCFVE0FXX31VeoO0nkeAeDIM31av
Vi59Cu2qUM48x9ACSiZR09z3lL4uGgPZPCisJYGa7oy6Ad9Y/HVWUDVvVJ7bqU07o1e8NaiZGusy
gUSWoqptYQD+GKUmNen2uVkUfkLMwR5lvKk5UjHxmHqiIj6ODCRAIElYNigYwHk6YyZ3NdGYyb5a
SEqFsEPrfr3KgJt32qzlloAbTGoHxIOMohk7zuKmgXVCviZZ2DbrEBvUKO+VsGYGFO6bJucNooZA
W3ukDaOzDRm+iJ4ecdNTjBlB7tLQygFjKIDnDGXoxf6VLO5K4DOZpzMk6mRxImK+v7i7L9QGjIZm
mL/SrMJC9xU/D7kV7bjz2rOEtjMZ37KY3CEQZaL4DBweDaybOFWbWt6Einnw05LTSbZS1jmI2AcX
LokqNjtS2jTxf3PmoTRBABrSy4Fpod+T6vIEOhhMqd9QOBwE5fbVWpRhdSEDWHnzHKx4sJ41QMF1
Z+flWWbqFXhPXS/hovCo0iZc0x+iPJHiP/Hiibm7T0wX2wFUqQxAeea0mBri2PAaqV2bT3N6oJ3O
vrWHFyQyXLQO5rpCOwf23zrFlwsJdMCC7z/ux1sWvOgvuBImHsA4SVZncTdrZje/1VRoRR3m7NWt
WTP4N3MCpzxxbEqn2V9QSay7Ay0gKVzBo+YoaRSPnRMMc/b0VW8Kwxq9nTyw187qzwGEEn6gtjnO
0/VVr3rWKYGGbDWdHTGbxgOF/ApqpGD3hpIoTpO2Pw30JzxjZwpRIS4JNLDIoDj0IoXeKzWDNYo9
t6WWRHBVu2Q6HqWryjdeEK6mlphgXP/TBWs8CBIR+ZqQbxSa/ZRn6RmvrHIilXDD8ZqvcssUzUn6
IzEgTjW9mBoOd/1Qc+JKW3Nvqm1SYh2lEFWjySwr4jq2es4iBi3txfsricGjl8U8BMr/Q3AtJDdP
BJPa27UUVFXzgeEih0v1aRkWcC3pdjIGuBVU/NYQuya6HuTVmUmUjiobbbfkUwRfrEpnp4YiB+WP
SHogWeSox7dAM7SQbaUI7L/OmhZzWH+B5TIX7HNY0yUqFtMtzf9AsUW7hYnXZ5rcfLRYOXUHgJ9P
RyIoYU23FEno0fKeAMt9tujr9fPyyoP9buqRYzP4UGwgQ3F/5hDXxmMZ70tQWSkaET14swBQNt/e
n3m3E97+ywGxGxQGyo6feRenUF/cP+MdqLaABo32yuWihNgg5DzdRY/jO6Agtw4+qibMwebMVKlF
CETTYGdDaQeUxGUuGLcS4cqBET03aaKuDJqQegXBFbXSQprlpdYrDvwWr/HRWq2dZQIG0fJ77oU7
22Cg/a7FdxK/LWK0fIbylOXO5BL8OUwkHiaHVChzQ46PrpN/GGMkwi29hAF098CODbEaz8+861y1
omc95hhQFeYSD9xxmBJOR4cwMQi5KLgezpsaEwNAvaN0AKAhTrIw+L7kab41OVwUpLKlX94XDsQ5
XztY6QbjXKaAlcxDWCqxU4DlN+fE4NfePgNou4eOniaiX7oEdgJx0EdvvXf8835kiDWFVY7Elz/5
fNZth9E3SgdUTHwvTbJTtdxwq3GUsGXew5Vv+04+FRdTPbbejgc7Fs/KC8zFQ/xdm2kyH8yE+uZZ
2QKrE5ozfiWJuB82tOCza15BPQC04b4XC77pbcph0H71zY3jCa42CICTvFTFGwIuipxBsW0NvbQb
uHKdXPGfxysS7dM6s9dcnsFGv1RE13+YY8A5wioaFD4Js43CVkxdTjrKWBI6ZFAmzcnikk7e3H+5
Ic8hWGLYL2hPsFPRJbZCGSfSRPZp+EKFIcn28N86gkTX8PSizU1zs4iZUri+Z3uH7XE50DGKQob6
NsqOUSwT6HwwrZ1J7PB4k7NQyyn7EFaQEI9MaQH+K4R3HoQbDFeCxa/DTPmS9TZ2/JgyQeiRih8/
uCJCA0D5ZdPdHMQfLfoWbJaqX8JqlQlMucSHe8p1/oZA8wp2NUXJUJJ4YVj8RPWuxn/bOEv4ebUq
ewZALbVVTJ1C4/ubB8jbzbuPqcPIgJyccvRGblksdsmd7OC3n0KLF/GuhTpy6Ej6WhEuEWz3ue2I
ZtZfmPIfDUTUX9TyyehkbJ/amjT9DMo5Y/MhrXtN91FQxFMPZoB/yQLG24vFJ3KnNNppLDfZkUdE
A+2fAaCKnsAdKvraX7R0psdtQGmBVpfi9EqHxfSD15gnJTCFGivZy8JlezWdOYgjzFwBdsvv6UwH
s2vSn2LDs1Owf0Dn7JSbu4zgkn+sc2WNElF2IhuqiQCJ9RhPyf5qDh0Hvm56l0p0LDY27NbZNPo5
deuFtUG0SD3L2t/f90wa5Wo2QQgL7H6Y7CzUtrX5RZCCioMsu/rRl47Kt9KPvnUMPRzsPjhmw+nL
x7DAn+q+NWmTu7K/G2bEqH8UTNsXUxJ2/+nOCbM4pYK6UC24Vq+4lmXvqnaJ2AO78EitlSvydI+s
EAr5agrMENNJEwMHxe8ThSedq7CVfhDeSZT+0tXN9Sltcx+QQTO+YQ9FGPRg2xfboClw/TpqUMP8
LY+HiKy1d5oudiGgqWsNohMC4ZJdXgHkboF0Dc6+VVsXmYDoJJAZuzkrt32W42+xz/97h9E0wH1l
eyqpgAkYG/UiRyU/FRbOw9Vszwk2QwSt1OgUQYQ+aVXtIlHvlgaRbV19WftIa+kmQ6J5BZZLGZmh
HYA3ixvklEQK3z21MJWv3cBwNGzdNxO4JhvCfe+4mI8AN+/7OtfeH0Fbr/IvDlR/Tck8UHpL657I
OZCj0o1F37Wuqujj8iqvKu505S5KOwVQN9LiG1FJmmiLFoxF6VwbDRcXO06v+XuGAgPQm6bvnu0X
x1cUx1Ge3cQvSEglNBll/DQXDSHYNEEQFmD71ZMu0B0rFHHySY4PEOYkL+M1lDZz4wFe5Lig85JZ
UaahSe96kJntrJioioegt9QWGu2T+5sTNv/TP8ntlZmirx5slgnFhn8DjxinjRvRCLcYAOsTS4+n
H4J1h+RvIpTaHNPxJFjepRKQArjPuSGdIWUo1kOC3EIn+jeK5Askw9locQbWk5Cv/cDZNprswLbK
xugk/Fm8F2SGcqLAkSLLZ1y5dGw4esTb+T+LfaYDbiyOfWaoxuc3OJEGr0odOU3s15UlGr9LZASm
vrfc+SnLIu1PNoI4eOoRvQSsOOBLsjhevu/wj1v6YMEmB3cEOA55bkRpCc5X/RELjNBbE3/T6x6b
6Cx6dTePSG9s7waiuwqFsd1QZ4/lGAV51gLzpeTqZEgohcSL/VdQUlrc1dAh/a1/5E/cXirPGj+l
pC/+nJOBmf8T/Es8SaF85L3D8kuzdVJebMTgPRBIA3SekIubTHTWfHp+4mc2T1+3xuGDee0ZyC0/
SlAmQ954xsX+UeAu2jCCBaP+5lyvXBlMqjdMCrd3x0bRUoNhKfmH6z26jaGaO+j6qBeXNjNoQczs
GJlKHy8CgGYofJDFNi1qzeuCYAJbSZyeBZbhA3WyInn0l8IGkCra4QlJM3squS+vUwmTP47b/00W
Pt0wErQ46DOlDHvxDVnhI91XCl8MfiN3IhsKUveIzCmmDH+kNtnEQr3x0CTavtcvNFcQh406Dt59
5rW879MWDon7T9lMCgm9siCVNSF5peilOtgiNh6MW5KLojd1Mgm2UEyFniEjI8KJs+4hu95XjeSP
t29k5pw3XUx+phwNO/T4fK8i8SFZITsrDiq2HfWURzVY5hJpOZHXdWgNbXbQY5k6h+tRc0QpJCbQ
lBDXfAq+vD67koQ2xQc14kYcFssxaL6zma4FIzARQV3s2A/K9lG3J/mbtDL2iUlJND6TkyoxlSsK
JnFF3qn6zWeqRmIAnqIF25bLD8Ys5IBKnozarXKEQAz1EwpyOGFqLYMTCK96mrGBrrpekuAUaG9Y
hym0oZcq6g2aglYNpeKGAFRpQRcoTqFFnZ9kotQP0GxqkroTKyV8LixUemeS1sRmjy8AJSrp2p7S
VVKCjDKaQXqoSu11pCze9I4gDQ2YeySmUguh7XI43cSsO+COY09OHgsPoANVsUlWmmi059BIhclT
wGUZvhpE1smqY5xyVq8CyfTKX9dIXNyhQ2nmFnOOisKWRUmD/Lf5j50O7cjLRW0NQ6dfO0f98g6p
ATc8gw2OG28WFq8dr5CCz6lT5GKQTl93IdYwWwgoHhtH6/XisaxZ2wuqdH2k+bNz21Nh6motvd5Y
GySGtL4A4VFtreaKG7Kw9i1iOs071fw65ZjphUxSZImj2SGKQ4V6OLNzNbCjDphct/1+cs6pdLvt
nxik+EYG/PMRiwJtFh9grFpry2AAhL+7ccJEM/BNAUjriuswzw/zW8onJXhJPHAa6da/GrMSSM1X
2YN+Rc3rt8R37/s90WQnEseR8xXrWA2GMsMLSYNsLwGAwL6iazti4ECjTTFN9yjVmpEYDF41IPIC
bufp3Om5X9d8e6XURP00/W/J50+1qZ1YtfYDlGMLrIhELhLPfxqFIgrTnl7r5QTF8Wtox4vfKTP3
+YfEHWJftA5FQIwSqAh1pssgWJRFQj9OVkObFNsU3n64yJyBJQMAJUY67TAn2bNGw/F3I7Ir5u2d
CoI1SX2cvGFS7IhBhMGX063kuzYLlc1E5CtyUjrMVaURMmd+hXs+K2Om1kC5vBLZ3Tx8XQDIsrKa
hEgnPhVg/IKsVJ82YyU9d/STKr5zzUpaFn/Tk7HlE0NgmKeuq28LrBAukAmA8bdqTxMKB5CX8oT9
Wy8JRZW6newkDwO2hnd0zkhNWP5eAei349fM+uDOhKS0hAOV1vW1umOLXgEtj/b4PR3DkUmVRPGf
k447bnxZZEzS6+mJ8tm6b86xe2huwzc78Jivjc1gC5nE/OG6Wrgk5S+uc2DAf6PVjZLMenBuyH6f
pTRwchiM5HpqDkn+Buf2KcXr/XcMulL/+YoMjQ8VeWvu/NImB88paMHDcGIkV/XkBZ3nIDAksEFo
kwDg/0cK7ZkBSEIjQzgzP6Z8F/F8PTDNspGu/RBtt0nSPuuxr6j8FB6O3dJsjmzi4EGOr/JgNJD4
OP/4xguw6aunrVXB1tXBmnn/R0EMjaYYSlOzjVJmJEigdgzXZhiexkuP5HQEqNZG5VbOIWn2FLX8
O7Dl4Nv6AC+ro2Z5xkiU8Ld6N0gYSuWN9UU9hZXchqo2BrqJnOyysiAOl4P+OK7fiE3vj7V/ACMY
H4MNCUuhShfE97jkCvlb/dtVRXKM3bi0jzQ3hzWTD6JgiSCmYPknNuamYty0qZnSER3IPUD6zxHr
prOZDfEqEvUzxW8wfn/iAumI5A7TESg9RdMN8BzqOzHBCWtf54TfYv+gopP9Ap8TMqbPRpOZsf/I
Ch1XpUqdXU+eCxsHsQv28s6Imtbo4qPm3LeZf9Gz9xOKQtAuhEIvjHpnSUOz0GcabStcC0PJcEx3
NvE2uo0nEMqeJKhkQFNbid2T/7VSmw/3RNyB1NmwaE/+T+PYh2O4gyiDrduzgjRM1oPONn0lV1P5
We8ph5aTcZy/fBTnO6FxTcCa6wuKIhc8fTiGUc//Ch2cMp7b3NbUpG5cFz6uLv2XH/NdxOtnBl9E
7AwhtnOv9tdQa6Mbx0mMOy8J0RYho/sriw1TaHoT2WEsvpLTIlUt3ujHwain27fKwCobthMepzmW
roMthDDM5Bpa2XVv8xhL4Yc5OPLCK0rqW01mjQwpIosOk+RQwcG0JuEHSG5oS8pSExGywyB8ky3O
DUqSq5OSbZK2lts94aPpQCJrsawsbUy92Q7ComuoJQ3Pr6yJVfHw+fb5r8SKROMZ/o0+x2fH/dw9
AjIm9lW14IyJ37eIBZfTPhHFzksD5kJHVtKVPxnyVuQ3jeT3ikAXyMgykpJFr5AOAhjBnHRkE5/7
uuk0LJUrS1kZ4JuxONPYex2gIEa5y54HZCZm+j9OIzgVJiw1p8ge1S7xsFR0KGz3QLjc7eoDfvDv
hOOVGH4x0B1u6OO6jS6NKYI372Hm5X2H53i95XZeV7g2O5y+0BJ+/aICC54Qb3B8KTvTmlSfvXEt
hS9yr8KWHpGsJlsfjTdHGP+b5A7w47zyPNuDTSCHsFMvVvq5h7l8gz+j3ShrIe76RggdVN5MqUZE
VCwPVAW5aCe7MDfhWLborkVLz8pj7gbZjlS9sGJuM/qoEfqF/yF/S36hzbx0FxdJYBv0q3hgdg67
hqnz+Xy0vA/xYij8wZyx+p4CYIuX9pMle8FZa/RIcML4qUqXw9Xxul0RhUUcN2R/4D72Bqzsapg5
JVuLTYugkdia8OP7wTBhj+0Lo6eu+SfFL0E6+3zlIDZk1HYVmRwZAb/Donlnj155pMNmp2z7H6yT
1DzJ07oczxEDiKSUMUyJPuCRCsPgFu8VWjwncsDacPoIcuFia7Rriwgc9/UTYZW0lQ7N1w37bbOQ
9XgE0grebmi+Ji/uosV0z+EdCjs3gbA4KHfW8Jy9zIjBGSFKP6gVxKoflmM+xDOAj6Fi6PEv5vQF
jqbbhfbQAnrhDfSFEV5fLpbRf7T67nifBiQk4FcmijpomOj74LhJN7ct8TM4jE6Gwhm5o8afZ/EF
IbP8dLzY7mCP2lPBJahgR1mv0OBqj1BCPnT0sjN0BgkK02Paw6iKjmvgMo8dR04dIxvZsUMroqrv
BycD8W8HMwmog/+DxAr+1e1cu11zJsMjvMacf5lOzLxXDJ0s0ATxjSg2SvBRAwgnOPbDLTFGG6Zx
MTbdcQCw+CuUB3zhi+SPhr7TAF/T41GZisXyYTxBT8HLDx81idpYll7h4u5IPjn7MzwyzGDPB4sS
s55XmBkE4+N+7nzH/hOJZYTyxLckR1SSYACwTeCzK2EAO8dOBVlHkGOgW+2G72EYZt0w7+IIclrZ
uFF3KXyid8QGzQyDO8PS644k1rsEm6hUieBnL40DyQouW0d0zX5EPRbuAjOYeHojR/rud/Oac6wT
DZ8Xe8Q3teGIUoKojRTgt6UoDKI6k/RPYq6rbZ4Hej10x8oJJspZB869J2Q6nagIM8p+84SSwi2g
jLGt9lKPmLCO8HlrDiN0oPgnXn+jheSn1YaGq0pMoKi3Pnv3mKmq9IZfAFsxZIX8LTiqV0RroSzp
tsA12Hhp1HDFduTuYZxFuQEJl9GA5U0ZzMufA+F411//3wuemUPwDdgiBfnHuDjwU9e5vSwlgQXv
V1OkHIPih7QNuQQ1nTV0FiIJCHlh9KQd0/L+af2TmYwKv31EszkdLc39VgnUBsnprR8CnuCDaugK
HaGp0ZZt6ddkFZ0AtzehXUQlkDOuEKKypdH9vxA7H2LB3FO3Q8uJPGV9NmOA/NhCVnVj0DrjvQx5
4rQoS9z02KoWVv006oNwsIoenSY9fDU7wY+G5KS6DZe0v3IOq2JtTtjP+kfHacE2FgN001i7gK7i
uNQ4yfce8LOxpcjN8NZ4kT5fMkaC9veaMRDqvrQBXH913nB3M75r/xbGquzsek7BAnqIN9j9P9zU
NjbqFfW2gorFj1/pCy7cVm6KuY0Dx51mhkG5ULWs9wtR726BMFBWWZ3Ymj1TbrQJPyOkWMskew2/
QLeUjBAxoiLzUUp1OxukBMJ4+n7kWt5XYcSRHOfySfBDK7jRhWXR0sL/mU7i9XZc+8LdlrLcMxm/
rbNawgb5X38GxYUfhmWcZE46LEdyY8VzH6mppIpz/mgokY5UXx8Zya+mQBY0zxBk59JkJK2d4o/4
QqdtkMlvRnRj9dMDiGvK1Hamxn7AlSgE2IxF4PBztBUEnnjDOFA8INv7bNPXCKf+Iht0dV9cvn/e
Lpj3b/PJTsxHRtJ6EPp9jjxvVTyracPLp7gCN26QR3upexZw1MWLGGP594i42I5qHv7CkINEIqfI
9VH1X/EGwALCa+jST7yymFDPbak6q1H6C/YuLFpHtRhnoWIC0mPyIqGPs/3MF0G4XbVMlUvZB1cE
VyD9aLvYoZqdNVcIm+/NQ6bL6/sBhZf8HQp7c13naG9fU4uGSVP/ILt+2BtPgiesG1dBWU0t1bCY
RAhkZnHE4XNydkzVOyNGYuaXkOMuPqepNloFG52xmFApM9LrjeufYaB6xoNUcdgKGE7+U5MnaNZb
otpd0RTmueNElbcpSbXJz7mfyzEMHFBdc+WpM1GrDeveNxgk0XBLeSnqqk4vKXVIM55yDunrGfxg
IsiuR3dVbvcozWEn9GadsJ7EiKRUMzLkrtg+ed35pnfb3xfAgQeCYlIegbPNwIDr8XA1OC5qduiu
FNPEkYV4Nnc5G1XmJ96HUg0I9u9ou9sN4q6LwjJZnlwMRXZMvZa/iTolY+7Zgsl6Z74S5QPlHMWV
HXH1MHuGy0tnoW0SVnZPwh9eILEeo1NIwQcKzyQS30NRuKbM0akU5BFHov99WRT2XXN5gPRy/kuV
d3NGLrCW3jBOSGKNAf8Hv9V/+pozlAs56Gn7FlvqhlcuAWvutqwvMG0+aOijJGWz4gzJgBaEHOAP
BPnMJK/CmYPwqVC/fBxZjYNiMEIM3hX5IVAjTcMZqZSQHcqHSmB7dpv/gEDwv6pp2IlpFZuEC1ht
pJCqVCXKPJ1WaOgTGgHsws8JoK9DCYdtOsbpx3Wc8P5ci8BDwO6HGRhfON1VjsXtcPde0V0As5OU
XsYdPkJoyV9l/R/hpesEM4wOGXZFZ4z6Rya90twYFfCV5MkiE7n4nbE3t/9sq4b/Ttoan9EX0kJ0
3B6CaTxS5elLXL4n/expBl2LgeGcDmPDVcWRclM0wroRXyPkXfMgsz0C910lOhBXx19jSo5jnf70
z5UF27d5BZ438PS1xPokcK9Y6PGDhvccN/tRYl1/r6EO8ESnqjN7MF2ueZVFM2QQ7SKyICSaa3H3
hqgJEkkS1OLVy2Xd5fayI0ockRQp1QN8zcuVnDfft/fs0gNGI5AMR0AsDKkK/4np/uPNfjlDCRwF
u28i53hHOa+X5YyfQjQP+/+QxKsGF5PBk1IQQaVes74S7u4zPRPcF90JUWQZLqHLZp7xQytOLEXf
hM/7rDKCURFKZueCirudVM7YHh2VANW9L3Q8tRqCgpn20acummKJaVzRnyxfpkNxwWEl7tmtIGkX
Sentu+42iA/jq48wkXetT71hjLm2flGayKQGM7KmZ0HLOTcnoQ87PaIqMmnVcocKrXNO7dQxSB3B
fYHzrNHz8E3oQT4/eZ8m4QEX+SPuVtx7UoHlbbkVn9MbdTROD8TOE/HGzYfX/Eeo9qDTFzo0BZF0
thJB2rsUHMSFumLFgen7CmVyPhWYA5Ah6GR3BcyoVb7dVfEKe+1nSm9+2Ecp9Z/c7WDdeNyLuFyz
BcNVxgV4Nb9QXvReufYiAYRPhrcsfDF5m6ch08MvxmovPtBq5GOqQCXq7xnccELNfuOFlMHSZSJB
UadQAnqW1PZi8z3d2evKl+z9ni2g06KlGj+ia3veK5KFgCmJqA+njiPzaX1WjgYi9sS1RGlm0OOY
0UO/8fXZyFi09ySpCwkl1wA2mNLqRBv8oGgJeemzNPWxF6O85ESUxgACa+zTjFnC4Aq48h78y11z
p8wHFCVBmCIWvvBBKi42XKJjlvVOSxl4zDWL3oHT3nuhIe0ZZ/RKuz1HU125n1Us8zNnaOegHBYI
Snk+aWRKbhQpFEZaPzE1Upmu18On569rtH2YNfAwG6N483JXpEuc2xbvil7SU3T0etBb84xBsG0P
eFRLKSsdp4Ty3z/x38KrIowE8mvWmJsMOhy3TbPAW2pgl5ilHAh8Nh5Fhhsk2nTRPZxZA2fZ10j6
i6pEqJwgeOGAJYZXEQJK69MrxumglQB1bhhMH7jdTBeMW6J98fwwpgeEamBvgM39jWTZXhVMW3K+
FOdVE0mzJmBdR/hb/6grach7+iQfvaq52O+SQGXl20PRB5whp1E/GRKd7o/A/2TY9GtVtC2xppZf
hiO4GlS3uydBuYlonrGYj8Uk8Fi0mfgAwkDk1Bg7D715GoBIxI3BaCKKp//b+WaVUDhlfgHiJMvh
D0wFMgi5miwevPyW4aiIRa08Muer8Mq/wf2FZU/AVcO7766cvgFk9ojJGH/8HbL3GNi7+NBxenlB
G/dGMGsGD/Kii9BR4yG8z/YziqZ2dycJWVqHZfc3Q5RgxsS2k3qjDAI+PydK8/K1xtn+MdJlKxyg
y3UeMok1Vhls1Gqb6kS8/B/neg/pYujXOn+8Ijo8dKIPpWd4vDcwLhIYbxODqIda+KuYtr3ekAXK
Igp7fy25xfzPL0Lp2ToenSsz6brHchprvbaSh39ffnM7TAEh7hO3BW+vlmR+GKq0SFaRCp/PfJni
+8hnRqFV4EBq50riQNNicBWghvmne6kw8HcK3a78C8+gqaeVYDu3nXvquCSGtNNB2w52I6QHcCOj
PsXSPSNqvv/DSG0YzIDceRYghpFt1F9HYAEHymzSptRkCW50ryT/vNge7/DxOC1PcBne6N964Edy
Fi1vRxCOC/HJmzoPki8vd5EyjiW6BVdqi+CmUsZqpqUPDYrA5T52Qhp6/7io6CqTnV4vShepO9Ns
S7wYYPDgyoT+A6kXRlS1XFCh9eIYdUgGhDS4gei++JkpyPWZa4T4/8rPOu5YhbjCq6O3PVtGxCJL
S0cCRqY524i8+k1pog1oQ4BnXsdZP4mp+UnbhILyG0hA/IPtt9kP3mPhCk0O0374LbHRsRJgVUvJ
hFAUlGaJKxxr0+T8rK2tkZah1gLJnnNJh6V+cWsAStTEC11Spwfhg/r8eWlmvd7H3uyshaXvbRSD
3X2fAo4L4OR7BNiXxrbbGlF73zIGNbEZqORCcA2Br28LTN3/yi6S3L7pVUr8uupHgJIroGEeHrgZ
rHV/45cerL7uFBYK7FWg82SdWxurYMNAYl+ORLW2N4tY6ZZqsfWkOmHuL7onm5aJt64ELGFsL661
IZIOYSk16u46sK6WSVNzj5lx98qORPYCidfNTnFv592WY9Kbqxf7q2Oymoumi4jvqNe25kQys3jo
hRETw4sfiXRMYzOigP9VjipMuQiLXqZ/eV9iW7MO72hCFVyyrV9Q87cVPxTVaPAIsZ0FkQB7Lb0B
D/3p0/AsJUs3hpJ+I0/+NRkbKX+LlztjgTeMKI3ezvldJq6Sc8mB0RMHw9Gc5Nn5YwZllLfN8KGU
GWbilFHzrgD1ka+8zPrWkP9yQzPLRg2oDbGs1c48xf2u13hMLBckeoTkDiv+eDcv9frVgF5Z5Y3A
l/v9wMcaEhoFQ2EQYH+Nw9r5xmHl9YuCnxmK3aZ/qUpGCn+YSy3YwRosNxo/ACbGRfq8yqJGut5g
4oraHbsMm0uEHJXJPIGYK1lIo57uuV5Ffo37f6OD9+mzFfKO5CzKZrnU65hsV2rzBR3FWj4+Zibn
9FeVoMgjpr6SXeGY8q46KDD83mPDwzqxg6edm1AJ/pRrhxf0FxP4RJFRoW5UkgMTYeQ82AMhU09j
K702X+JTX9ZmE0lxCLN5YcdSICESMjMOkKGJ2tDJN+xHv1+VuVQOC5JHjsFqhI3LH2MZ6NWakFy7
JpmSK+iPv96KyDG6doD70QPkqj6laM1/3KS6IuKgQx/XKL3G0nz5esRHm9hSCBT816xUIc/2vDqo
LrZdF/7GlyXvoqpu6ymtlfZDhM8YADWdaGAamvAXLlOWFQ5X9oE0LmKKcsHTgHryyLWn4rsHAD4j
IkquE4Z0ClsN98C6i30x97Y8vgIG7/Qoxq4vepjmfIuGypDTunqScMC8kOdPzb4znK84bEM/Hx8j
yGpxIQlQOUVS/20SzxKwAX3r5UGvfD/taPsHTBEy9Rz43U3oSelL+IDTu3pjrPbXvsZkaWfFGcgc
afA1OG09WpccmVrOW7HoSm1fPAZN2POjO57MzjSnvRY9ukd+uC1OJq7kidGg+KZogIdPboiIf3uA
UZlbblUwF6SYAUUxX7xok64rS9NaOlaXVVzAWX45647spIdPDkX2ktqo6wSL3FzUZ4Ncrcg3fHvy
Mn7KidyAxRmHT9Ky3WitJDr97YZU4hBhlh3RJk3xtXnM+eCyac4t2otCkBfNHIKGmQLryBm+FJm3
U7pHwiYSprDMkk5778llSutPHdnd757aIHefzdVxN/6hgjaKO/0eCJrN6PPYz2nVgulKhOVWOTw/
eF9NPhNYKm0Cyx6DoZrm5MDmeAIqFqql/I0QnTS32NHD8aBxjTA1A0k17GvJAUyqtTnsAO9zoVGu
8kvQl0gNtFvicPQzrrF7cAqyisd2yG0zWaBQ1FG1fJjqtMl9BsJmtllMGdTNq9vJU5do6GwPMClL
WTC2LKcx4wfsypNexsCdyx2VNvESZ1fjqv4+ldhFzOhDMTxLDA3zZTUo4OKoPeaTEKxbqXA28KCr
rtIhaV4/eJYgw2S+/2teXDE5+Se7xXWo6/Byl4kVH8dmnd9nt32yeRSpyQTl+N7T6uXKaLH+lYWD
RchO6/W0pSTkg/6s9eyISg9i8xY66qxiFudqE/0d8QXfa4/+mEDhbrNaikta6Ne/RNKm0I4xM/SJ
HvHgGvmA+XW+f+kK7MsHEK5qe7jHESHENMs9MJV6s1c4uy3tWp3TUNAggcxgUSiVo7JhnT2jSiht
9QyAU8lf3BKqrVv/Dui2+e4qlvbKFK0Yss68mjmTqP3f8LUvqmBEjRQHUy9U19ZwWLwqUlhaRqzF
/s7fK9HqpfVlXhasFGnvQ75U5nLFzNA6mDmxPLcVn69evso3w2B1cP9fxFrR5RVMP4zjVb6sD7UM
QWc99BWv5Dbb+L0WIsS7zxNSwHNR157GbW9fgng84jxGJd8JaZSh6xeQvQjzgTUeA/45fMPij50f
x3HnDsCfrRdGXC6URN3kxpZtkaLOmIMCIELSIpZTK0TK4BMOQAR9n+fu2Y7CmHy8UalBHCei/51W
lPi+PVrxY4/qWQ0i8eLT5urY2Vr7kEptq9Y39zaHNyKathETKXE38qSAyoT/JJQFSBQU+co5HWAs
uGh+BgKqdrRm/uEt18HI/7ia/qcyGZcGKfQWk0TSD4P7mIdLupWAmH39l3TxttJnUPrhQo98WYSK
sdS/vZiqn/0HmYMENXYmYbkJNMeWIZEAb3CIET5UFxpdqaz5V16KOBfHw/N+N0i7FtsdNbTnvI9o
DYz9OlYfiW4IB8s2UK2xOMy0wqu3fYNqayYIHyQaM4WgehMHfcT1fpY0TJKAxP7WL8oge2Mw0M9f
CZdj8qQDlppF4uVvci3K+uyXtxXZOlf+Sp+nUX4v5TQQBrpJtxKg8NNTSfCca4bq0VlujYuh4O7L
frqCnxt41ny7BbiiOX/P1lvdIvqMHlyoULDJVMsjLnaBrC3+TYXZbVDI55OqAYnrYmDj9j7B6+Pj
2gJdp5rl0nH4tp0in0W1WqXZmq5rJh4mwjgfQvK06KSbCVWtInaI4P3Y5JmnhkEnGjt8Znrv0a/n
Rr0hHLGvSHmEvHrV4H5A4Pvjxq/bL9hhz9dvAt8ET96HacsWmHKY531y9OBGSqDASfPV5+IsZewS
I3rglomlr7HnpXbG8bGGDQcUeSvVWxIFDy4imE4ZuYeP6HV+Hi95K5GKVwka2SECKAm7eQ8f5s7n
/FYfwjlMslChQCSmklhdOrLl2r/FQ+y/6rT0AUdRc/ZFl2GahEO4S1q81s9lZtJpiAZMJeoN0Kxu
Uo6UzkFBj+gJOarA3xxVyP4HHgGivK1bjn2tAzbi5yg4dUm0Uw4lZjw0QtulTITnnFqjGUMt/9MQ
snD4lY+0l2HQQMOYRuHbMRfkK8iMo/LpIklqQvVw+nFd+I0omIySCkmUOy9rTWG9njCm/n5THHh9
hULMPR/aCKw5nuuYN9mO4vYV03zQaUPzb8IG+sz+2RKwanXmzKdqGV6MRZHEeitcoTOq6e27N/Ar
s2V2fEz63GkDeSJhe1I7uhxCZXxC5IMln6KVYeTHCKEPE6fQ/jZOU1JNAyY9sjf7Lh7Dp+6eQwWK
wYvqvQPv+9gwLYcVhsjR8RoJqAh68ORGj/NDYL6gmgtT+7EMK5fpechBZac7Z0JPNs8vyLC1TAMH
z8dAP+SgCb+b+MkWoCQNyzL+aSOpvuVTi+ivqOj40BlVCpLKwurvUxDwqLl8pAUIai0rm7ufY64w
K++WRMajSEvC5oleE/gOYMN9ltKBcF/tdCq1ouSe/5lpn25ebtMwovM4fDj3WQNOdr5/KlFpM899
N4sN95MmiWjlo9IxXHYqfOcwmOV0tA+6eg/it+ELjanlvZMvIQfq6/gz1bwH2YHOIcw0x/mEJKIk
zn0fF0ehVax/4FIQpqjHqh+IZebMIAkuXBZaDCzhCsH+genBsGIrJyPP1cWgguMXxFlqBm53dv2e
AZtblQ2rlVZYu7QsgxYJskqe/p++lkxBNtR7e7JOV8vlLT0Ozc4TZT6QCrLiISNqI/EU1P7Td+YD
0pqiQdfPmw64xHW/lIrJ6rJwVjJzgXEA4kCM6eM9yATefixNvvRKdSNvkLTSZ4Lu0soKmzEcoqfC
o2iiyCBLzN9JS0FnnBuVBXBlSvFm2pTNN69pcALVdicq2tzHJ2DtweR1Muee0Gax8CHVtmmqNjcI
HuPLS3SC5N05a2ZWfx45HnIFja6FstX0tydv5YXNF/Qls8uJYh5KeMnosMNjiaqH4LnBpY7Q+7qF
i+K2i8XtiyIl6x0u4W0HNiMnE7ylvWFCOdBS5AOANB0U2cNdzVEQdO7ZLHcigEfB5Fk39l9NDBD2
iEWm6s0ENLlZmEYYn4XnQcoLXEei/JLoT6BoxtyHJZO3zuwHPVylfpgnlF6S4h4E+SI8E7LFBiG8
0JPB9fmy6lOuH49uni9geWKNyT8Tx5Tq7dTBbKJDnHap27azCd01RUYYOpq6Mcl/uotx3rBujULs
eVO57X9/X41xNE90S4HODDRP8F9NAHzNP2qcCQW0SxguqP/Fe51gYcNoTixKTXRNkSbpDjcwNAg3
yZYtzWs1IPquCDub44ZGD/pryRwcw+WA/eUkVQZTb6kt8hXIXeT1O8UeAp2c3+CfxYDREUvaAGJ5
ULn/PThxFG/T+rX1ZEbxUuCYGMBgTp7x1b8mTtVSbULYVxN7O7DGHdFvBjQ59zBXvrkekA4C6vRf
jvTgiSn2EniSMiv2iGqbU3obW8LxL+Vd00sHFNaO7X4XdZKlB1fvRMRx51qwB/waJkfoZmki4V9k
JbmX0AQwn2OzqgPg7J7GQHUpbZyLTqX1g8hNSsosgPlVMkPwOqLIYDULFuJS1u6hGRg3Eirnf4vp
Yk09FRFomp8/UDmQm2kumNqzSdHiPvoSmY0FavoCBO1O8B7lwnlHSlUfO8MoW+UKNplAp3JAKa2B
q5tXnEXbQeP3h+N8RJSqP6UWu5PRh+m0gYvP+8zGICi2slEWr9oh3QJZF+jEcTvWVuHPbSTsEop+
8eEHXBRizuinjsilLloXfSZmaZYVKdp0v0KT1aRxDq5G+wD0yY9Wqo4F6jf9Sf8dde8taq/pUd57
G4F0/sEH3xQ8gL6//O6foagIq9XOnMZvRsm2cVbWSRGrxZBAfzFnqrds5UnLQAcbah6Vz/r1Y9wi
u3egssnadbKb0ejT8YTTMKdckd6UsiiNbo/AMxRDTcMw35tEuZcBAHz06U/LtwljFJEhVFTzr+/H
ef3aOhOaP6YmxYne6MKGEakikg2LaUsPoca7d6V/jo3zN+zCR0ObWeLFsXzqQFXqaJ/7jj17QtCb
lN/GiYZR4kU0hG7fBZzdAjpp2eo9UkPiTDUEkhqlyjB3exrIWzstpGnZPMxyeKluSwKMgrJ35Z3/
OUn8tCSeZhHxc3oR1LeA4uHD8VCya95ubSxfr3nJ+qYsq9H/SPmywsG1/rAEIsIjad0KldajADco
vaWURAHx4KtGV4mIp7coyXs0z7DaDak/SMpNhNMsN9dmABPI8YaDPCHlklPiHgF+7vCiav6mr8bL
4dZ+HKKWZZsLt9r8IUKSx+gcypfPmsXxfpykJ81PTVWyvBEj5yJJzIS/celtp3Z825X9DGW64PA5
szhgRYwNr9UTObn8Zp8J32Yj+JgGHqPMlS2Hsx4E4WowDNKFkwXW9fdsgGAHL6RCXSVivMysrgJ6
+oiUhpCbopbZz1K8UETdoSkZ7Xt8m6eXr1XuCzZrULkwRD4VTQruGaOYECkZSC30rOJq2aDtJ8LM
uIsGsZ1E1WDFaIcNcBFpH9b36MDLNWiZiNgj3qtx4tqQvbZD57/GEQNMEiEM9gJR7qSPKktwqR/h
IYSG7UAFojX2ysdbL1WPLSSOebXFAySqhlsA5+PqEVnQoyT1nN2IAhLAK8nRW/gmAzAWOCrGEg0Q
q4yCI/SE76CgWPbBRXKEL7QrAc3sO8V9BSUeSE9I/atBvbyqT7XWAycQAZkKrT6c/od139e7DWCU
8J7al5RidhnaUFNEikExtJKHMROqB6+FOGUNfcXMvLTvP0AnK1gSOXqjQX/Uncmrjs3BJ/7Gvs9P
sT+848ABZPrmH+2nXuSA+9YAsvBmsJW2pfIfcfus2DaXH1mQSbLqK4pRCpTzKItvKS/2hv071VNN
3g6q+uQMHqJjaGnhCTrf/GZWPdvCCV4/fGBF+aESQFFYKMOGQYGzRZlSIs6NIJMO4tZhI2WPMkpj
9PiA0TQkvUBaEQYEEagjh77v1CtJJHEyL27zSpjKoNSJkUneuL9eowjQKu1RMWs+gu3i6U2I+gDg
KjfQ5FIof/t6XN80Z4B/iN8U+rybyArQOVXhEvbUwF0YFzZcTp4VQ5gf5O5LYqlPLymPzE5S1E/X
E7Z2FMY6PB4EV9KSyBoNYuo6MGXXju1CWdHM3PIKF+i4icj8DD30lpntxqloffNULQi4xlsllaC/
N2UkGV32hq0ezMfewj61YTxA+7OXWTVQEoOXDkzkUtZAF5atnr0Y3b5MQijRC9oLgwroQ0c3bWR0
v4VRc23vN04Kbk5B4A5CjvQS5uX+ijF9vKp1O0lmEu2UpPYeEPFqQDCrwYRa4CRdRKLVP5reYSfJ
P7cfV+/nMTwQ0TYzlgCGN4ZGwaixj2D1TORWcuCM4B2bCDL9ZcZlNPqm9ay5nSbgnRaT8aDxfgQ7
HRSqU+X3rHNkax/ViGjYrfqrLJqYyhioChEm88H0yMtSjVahCUOafcz4Qg30pco2UdILzzjhJ60+
gThZQJnpVqvxdUkx9pslKaVceyjyIgibeQOH0NnliIx7NiYuP79FGwPO4+ujYihUTSbWHVXQwa5m
pnyZgVGwouxs5I7BrB0dlSwehpvhRFLff2qAWh7iF+A49ygzWaN+IwtyAUXIsuLnpVlrFNAiLzNR
nsKdWYt6LV++4sp0w0pUgLY11hJ1bnr9c2kNkX6vYLc0/lIwsJCwRzu6DSqJdxjpW04LrbMTiA3j
66gnVk2U/sf5TdN5+1Ag2dT3iHCSyoINTTZ5BXshYzWEj/i0UCtYEf+I94eY7rCxcDlSlQUm3xyM
55mF0pjEnBqGzHPy9KOswcv7ZQsJRyFe0lWHL2O/dJJyDMLvecdR77+/HkcjIFq0RyOyw/OCSt01
rTyeoYHKPZ/+yo/7Ex/I9Q1DqsGig53tLsV18TfyOWHjWV8rwEQHfkUuO/Va0yccKjegUbh6ynfN
TgmON8V3qJvjr58VtFsWQFz2MT8zKi5gnEUyE9oZ6ZjnRA4zsjOK9EjCAxR5YODr7O/EVtDou4zq
HhS57ua2NYrGIjFzNrZ9b236LiMQW5efUEG5i+uudpkeBT1btdlDycsvzYLSaCEFFYVtOlqT1k+l
amGhscUa+UmR7e3U1pNnpmDchwLT4P1Pmjjxs8mH4v/8iEv/AgqgmtpVPLQDpv3jqJTOlyOmvipo
hptZUvt0e6dFJ7GaTLGdn2XiJTwfQmdZZjpwHc9EZE8uNXwXTNtv9tZTYhMjcHnvjsyuiTxwG+JJ
k6y3KEQbfMsCjr+PxhVJB1MVNrFHmlapZ4owQWZLoutgUGUvmCpxRfeheYob8OiSIzdZvkqyG65E
1qhnGGJsXrunEOWW+G723LKVgKWiChauj620rRJy1S8nEMHV02YnfWLPV536anxfdCoKenwMmgjS
nBPMo3SqH12r0e6JwrE+Snx0YBHCVUMt7ekVzymP4ID/LbPw6+DCfh8E0lJzaxIHWt3s8JUsNFjF
BL7A94P8a2aoSKOO59TWCjaLyQfmCJlHwpOamxVN0Rm3zfV/9U1MAM/RzZ+RS03fhwMyRQ++vOZj
L+5CVcpbx49QlApCrjYpIwkV/ymd81SMuLN2UI0DhiQAjcHLIa9JIXQYHiuAmINy+Qk5eYOfPOYw
roHKBN/6wSpHdqZl71H+YGFnyOgrNxJoSYBg0+rIAnYBhPaPCEewr7o3QYnGD/rN38zFJkOhcstC
vQvSJcSFDxXVGrQ/BY6CXy4tNNHpEKJkJtMsKn7W91JBLUhsfzP4P7eKyxXwE2ir+ZefL2ys7G6F
f+bz/Ogc4KIGWCojF2Q4cxPa3DJvp6jhP1L1NP1asXlXCH86F/cAf6KSxiJFD8MXgU0jstf6rVRy
Faeyl4xk4BsWXvz4o7tCS/9/aI34RyULMpTVzWTrGoT9+hiSfO2BJz3CnjFcRJhuPL0Y5X0+938v
qq2auGmdarxtxdmtdK6ZjnUqgVcHEbfAPsoQ79cLQ73XU/9cYyvmMeifjfFa/uAoKSEnBf7/TnVF
OVYlxoqKBW3FAtpqsOJxNbWZ332HOa4uoCIjTerBOtX4tPZmPlvf/iJMEjpZhTB82nhWEEtdlWTd
mg8kj6+cAn1PXgtCWr94DhGJ0fAiOSGVWSF/3a1BB+S36vfU1IA50CIUl98QWxdShFe1J3OwJIZj
uPgtUiakGF8V4R7E8hciey81AYeyRgJxGVbnP6+OlEX36Go5u4jeE8l9qlZ4UzOjTAlFwU4b9Pih
TSqg/NAy4NFHCT7Hi1IyITBLeUcPi/7Z6EKJ+OuSyWBRNzJa+Y3CYHJ8aQbfbPK7UP3M8Zt0Jb2x
O+avgTApnWU5joLSS9/joiXoBcYGVgObdh3JsPwr05iifqR/2vTp0E2oiewhnQzDSuqkULzEJULe
5KvuCDRSBbz+UGYQ7UI3l+JOGukcRG3fKLC9WeA5Qn0K76VquCtjugtdODOVtPTO31sNBfFru8JX
eXRX0uA3Tlt+F2TCAzZwnfjereeQjtTiQPpnjPYGtlg/KAcGOJQjCUYg/D9HkzqGs9/VxaB4bFdY
hqmEwVqqxNOfsfevSneRYhLXyREG1TMYRLad+ouQibQdVRzM/XlM8hBSB6d4WTnLwt9Ws7G07R3/
r5LRFK3iti07F3l/N79zxlT34d+Kr7gZAxcoajaAOFMcC7qn1qSqA+3MHs/dOLu95PBSjqx/DBy2
uvKd4BVONacucK9WxkQBLwiXjfzseLDMrMH+AnprCQNVBFxupbW22t1Aqcl7XfyXhKWL23RZCZhZ
M2hOCCdoSLyZS2SbSoiQ8Itu2uxayuYK5hbqrIfXGgP59zkF9ndYo+ce0VQNiMwmwxtVTS+2aQN7
3T0k9C3ZzYCPlILqj+il6jBa0MjmK3s4DnRpNuElyOIP+7u2Nw1AqVa5aDSFmFXxw9tN9o+/EIEs
O2JDw0fv+Pm3Bok6I9dI4Gdq0LfIKcT2cFTj1LyzXP7n/kOZt9PgyxhkI/zd/hZefy4tFSe6xWOA
nxftePg/7aHHt5JhEm3qWFsML8BT/vIv7cb+cglNw48W/NJkoEUPdJmC/w/MOqA8a6jbUokYdfX5
1Uorv9AzxTx5nnUZpWYdXMY7Lel+xWzYPZkb2V4hHgmX/Tt2cu2+kZ2TlSuRMt/3SOs/ppd7+RAN
HkmofO2itobGY45NYRInPI3Khe+3sygSIpiImU6biX2hhxvB0Cmpe0ho1GTrDLw2lDb2kPpdL/I5
SEI6EsS5OFiRMYB4LmYA8qTpd5abK1qepemZqp0cuKS50/TPg6zw5WrVn6ssVR/L0bzMCvZ/8A/V
rCPDugxA/M6wZU9VU1EQ6pQrcSfcAtmnz7pfdo6n2MTXR3pA8EumBaooXIH8X9j0DVj42uvKfTYu
EnrOEl9lKYQ8dKJ2DuRtMfTzgL/d8nTsFfIugpA3kc5E/GpIQtxJK2xD5EGLgN9EcA6Ze5aKhVPg
IaI9IdqKo2GkvwP2FkqWlFnWVMqMb0x3kQMUKWYeTwkHLYrkU7BWLf57kr/dbaSgJ7i7jqWWA/Va
PlYqMxFLFHV62h+BV0ENdWGLeN2WHmx+WQbxHxwuntmpQD99foqlashLUjeJ05aGEI4xo0wZ1jXV
kCmZZQfjLyboTJac2SGPz63hm14H8BE3SJOjjj6j4YmtzwLHORNiOQ2ocKluPMAZSL5ssZMpD1Bs
CSNWDeifAhn5/S8pD4gb3KbPHpGwGibqt4GdYeBQkyEsoCt3QeprJ2RKrJzzWyirQTs7Iarxbzas
Gig5H4b6ZBNyFnhCH1XsMPBgTHbHy2yRNu0YHB/3QNqzh+ofFdVCViViN+AJhM8qsfap93LL4L1y
h/GvgyKEd1r3wOoSr4ZQgqcaysfJ3/4w24bQ58LoM4zEysr+bsLRNopOQuQV892XZreG1ixkEbUR
y1bX+QEWvoUyAlanP8kk7Rpviv1jNDhEeTLkUyPPn+O2caoz3IWms6LlZBXL5Mpxda4MZUEjtRYl
hkqmSWC0T3j0Ua2C7d5gF90WUZpjwHNdFV+v4Oe5vbYV6EiWwdgdQpEGqmmGPV0yhqLEUINpoIjA
ihg1I3bZr+swOssstVGfQr8fBLjArVRCpDKI9MFD8kUQRejH+oEP6NuSxm6pXp2Y2pU459W+cfFL
kjYi5c9TaAHtuiuyVQKLAR32E/FzAaKqld0ZKTtRsKHGQy1dxM+rnZEbrARKZm0Z/n0aXWfODdh2
/cfFmraCfZhkH+hIdOxcbQoWX1vxQXG+FpPSTHNPM+lAd83RJoboUW4MhwRsoR9GN+oMlCy2GWIr
aCRm//cp1w/y96fAMyoLZiBBoN5OPijS5zVGsFqM2tvnRwL5Wcn8c5neSYr+HFMrcsqXwjSMzyzn
cnV2ZJIuBOL9khcsL79gaRyrLhaV4JdtQwtTwpBqtfEGQuTQSGJZPJaKO/8DNx+1WaBLZgYel5I1
cd2TYYf7x3M7HIMbl6i4AWLD5BCPRWSYDgC4v/KZcMWTZyoAqRam63PvIHMmpN5xeJoCb4j+RiDb
VXxPnYkB4VO21eVhT46m59Ft7g8P5q4eZWu8P0QtXGn9YtS57gGrn1VdjG7o38VeISDuD+ZNZbVn
DsSlwIjrW6t7aGBpkOexGpmvOrIJF6LUGDw9i+qw03c3WueHFh1SPhFPpFwRblbQyZX8GjwuB/Na
pZWgFE1Ccnjah9nxFiN6axdUE778uW7cDpQgtVIMHWpIz4pBnYEJIfLl87dwSXsgsF1kQc7T/Zuf
Kp06M6BIcZMojKKoxGbTkDH/8Xo7DHqRy8uwts0qUQGpxQ756DpbZVVWRabD7aDckulWqsKALtuR
jSR82QVTum1YedfeROdvAp1H8dYCPTqBX1UQLGhBS+CznhHkZJi/DtNmQkZr0Y6K3KRMVcj8FiNF
nN0CbBBpNSHK9a/W3eGQ09cKxXSU0aCIVA72qKtPzNzP9ZIJSLifLoxPtk/Zr2C70zQVD4mZhPmZ
HiZTLcXeOg5qJuhZVWODldNvreT+frWhw1wXkJxFdJUvMJZMY79w/TPtb5KnZRJSP3ddwArQOP2G
HKiJo5xGlyB4Df8YY1R8R90DAyAnuD3QSty0KTQmJX2T/airyuf9CKrw1bjZHYjPNNuWR3JtirFz
a0MAeMkJsNrNrNg0NO3zhqiU+n9Y4YNVEUHkWkHdSy6zOks0LBYiWzWOupv4lzqPUgbtW1SOTHrt
DqU8lruCNhZ8cuLhHAnrofeaponBs35UXCO+G3zerrtQRSH84hbgnQk2OsJsg6v4U/KnO1K6kBD6
HQEBp5mW4MuP/+udIBkwLoyNH+Ddo8LIj0lCOyZWGpClWySOVsJRcOJuJUJV5rqYs+oPGP2jwKuZ
y7Ev0K9UM1o5WbVpwp7s3ONx9sisg8+5Y+xw2oKEfbbP8yTghGf3u2vwjnvKndZBilRVOuP3B1xl
8uf3Kwt5fEYxs2zsBNqs9mpzcSEAS57LuROq6jaduL5HZTHiZpCgy6LbTpaD/fafzEp1g0G4s/Cp
+o9M76C9CtDne4Vvu6TBtSZdJ7OWHgjMpwUob+VYWwktxHzr6884XAVp4KRGUjr527K+2nh+VLx0
RE7SVW0nuTZ6Ue30SVedQiFuoJYifnP9h0Ww+KNyl9DG+w7cUvK2dt3GV2Skz6CZZckkBZmYHH0X
b/pNvaezvMWsPl0rFO2v8r4yfAMNHe7L8iXQ+fqQmbhGMJDyUHtUtGzh5LOWgltPalh/j14z8Rza
g4RV1PLbgRzPrzpM4q5Lk1JMSZx7OZcgxlJQxakfsKs5RtyCgiTX9tK0oBkT0Y8QxJqFoc2Z917e
EIinK6Wd/WKu/pTSyKQacShpV9TZVS/A2CUPAIcZNdz/f+YA3JHeNcciCm8AAG3ev+ZUuZVIZzjp
985xtsuEqVJxQQ0dwsiPwqjty0/gbV1KdHMaSCWlJRugw1DZonCNW0+To8CY5phHqZBAXIoYGdnD
JF304sVlSVs1tHsnrOWZf0AMxBlWLLTmFu1kVjGdb2h8J7q4b/7IGk128b05P38u4smrI543EpFP
ycjE892q6D3wJ4pZBsDvkRCJ4lg9b8arfRd80KALcv1ElcHoBRpKSJ4vrtL5nvmdFdaZNkViuTI3
SOySyYRhZmkO2yZjFOJ2XwQh0CqnQX0jPHa57mVvvRY0LnTyKBb4GOIXiIyJEWWqO7oAYqIhcoKt
mVCUzbmgXElv/PihOwsQ60Y8J19gaJsOT1/tn/lzE9j9zgsMzEV/KfP4QdD+WDjcRcSovqajmAt/
M7wOcN+DDuQEOG5ztUu/1ePGMupghKLwaPn7z93cBqWCQFuDxPu5ks6qs7chnifwE/1+XxtB20SS
jFzHLqhF/003jxD8I00Jur232QgxqlNxg8LKSkp9UMxxA2sXPuju0zpBMBw3fJfM9nwzsjv0rdcj
EA2RLO+FpzlFD+wCPaAR7OD+HF3cpK7rmp/dvkS6BKnJWPIpkBzneVlCi21KGdF/v79GK5XB74X3
DFom2xEsBjrJwe9z5ex3rob9mtfJbU2750VSHuze9AX8YJ7AVvSph80UDNOdTaQOrtsiTKB5n72s
2pA8Dfumo8Az3/Nncc/fdwKUyECkf7GcrZ53hp/F7ZaHsQyZRz5hdWxNrO6lxaoW0bD18jta69fY
SeyYdybHR/oGQyxMowRabdymWX6QmW8Y3mIfOt7e3whY/VjrqT+F6/wzIrcJ9aL6X6zknZySiBQ0
deYn3jPTW3iUxbQXLC2N6Vs5X+ZHrfnVB4cDLAl6YgEG3ffGJyJ+Ma1Jg5zNYCW9xltn2ReHXv+o
/4QfUdXwi7ApcL1k2Uuw7DkvzxoFvkx6xB7SXS7/KNhsaOkbnxRDt23sPhHM5dbEWbWJO61RwthS
P+sOmgxb7TRUORZ116+u/98UYFF9AMkN3kUL+ih484/TJLMv/Ye9uzj7B7RBotwm5lW/tkEUX2e+
MF2+l8LyfLkkyLDx//FRKjuTtBNPC5Bi2CCphf6iBArdsHJdw4pcNK5Z+/zL47GkkDW0EntjTiVe
1rzwWUZ0IYptLgsMZ2EdKFzXc8/c1FlI0lBDFEc1J+ecdaXZEBN2B1OplgPLyAKwKT3ZmprYFhn6
3hB1s2jeZFsV8doq8Nj3gtW18Od35U2at0jFEg4BJKfXCi+7wTZEwKyjhHKqmKIkpaId7mIEFT7M
fjp3mkqyhFP57HJBiHdGmt6qwFVKFNyczjJf6erzEXSsYBJuwV5Zm787/gZYZdMn0bCb4n0ZxvPa
WG9oHER9b4TeV8t+iMMAT7J0+twYi5Hi+q/vk0dOQ3eGE5gx0jK/8uQ3kPRv5wmZgaZkCig3T1g/
6ZSI4WcoABRFEnQopPPIrQXX8SMIelU5VIfzEcPhFPnAAo2o8zKmqwkOzd1y21qEd434TSiqRgy1
vWCKwArWyo4G+OroReInqsBhQkRhJfkwcQ7ruCLqIeedbqqgGZRRcSVbp/GFqjt2y3CMA7WPgK6E
c8Nk5ac50YztdQ7xjXGgVXeqe+ALf3wacw14RqSpOJRqtPLCDUAq3r808UmWM/DkO6gIo6u1fBO6
HftO3xB5c0A5CGgZ+PQKlE1eAiQ1M0G0E7+VYrBu4JzP3qF8nTeGw00nzW82VFsSRmfj1i/1e6it
YGVClUeGGX8Sve+HlkhX5NEz5mr1lk3IXWdsiRaMb0Qh/6FCkjzhc1s/NEjCEx0fEsPnRWA6vUYs
Kg2EAUfPBiSxirZiODfONYfGt4TQkQ+KcaA9ONLZN2LOhWJm40BSEhW76fK41r10rPTGkgtOhpgR
R6/fzNFMpssPvJGL+MDN1WtT6GrI9+OMYreCgmYgZot0Am8w39qcOEtYzaj8chD/UWS7AM1pZ0UR
NEvrw7KITzuHFk+AuTaJ7M9LzTix9Tt5daLDMptQK9osn7/PI9t9xtNq+0uU9BwWovcjrDlJkujB
kkJQmL8dZWbJiFChzCP80YhJfSathlpZ5M6u2x3HlwYvtvo/J6FMJycdVgQpWEeouuT9apE9F6VL
JP4YeozXG8QuHa0cc4HX08e/ozuog8jkKyj/9qdDNmiksRT3DUSj6zPE6M/a2A0KXUbXN1OEnTzE
kAMKCvO4aY7Jx5UgTfUznPiOEnedUMzsmHW+SW3LLwrQ1bWQJz7tUIzpH3fAthGR42WT1MI/1iI1
/uC+AJ8ZG33We5DZoh1L9N5Q5nPnBeW5BoszxlBTZRoHN69uAq/bxT0r2N4EuwrAR7Pyr2yJHZRt
vQWHfRit9MgfgAaUS5GUIxAf6AP19voRZ6fMgN/GbkrYsqxpwQ5gkVsdh4egDDQFeY0KBXeB7uws
rqokhvKdh8MPUB03NiEajBXLMedRqVheBs2DLvNwt36CbVqvLHN7E8tj9c8wuXS4USPO49EpJ5Er
UGLz6VoV5IkFCtprLLjT2Uf61UEEk5YtPFoXzeOT5t15NPRgGUm0sWEnWoYtRagfR14EkfXuQX4X
KMTiqCAN6BSlItr+AoXULJFh+39MRqTz+8giouI/um8+uAv/U68Hln5LKFoeXAq0UsiMIQbRBDO+
WeZh8dFqZnd8xE3aDNoPYgND1L2hwM+9x0BW2blN/loEFQMlELdhro643BQXabWghphRotl2gZMv
6v+QWQCCi1ElU1egoLkl4FpE84xnGRP0YAJkSUXZKTf05TKUBWi0EUmxf1rkJDSqATiaEddgmSCq
vHhzEZR+7Ap+YiY5Iw1Vim8fbp0mAWns8goHBWukExAf/3f43MV3oNg8GHoFMm+7ALRiARSInnu2
i/7uhIpDOHRENCH6sMi64sHPinBb1LPdUTrFApSgFms9b88PpvnLoWavNOED7+OdzKwWb+AlJzHr
s5nuPtFEWrsAyc1eIhscVzPg2QeggGXmZblML5Ri2bJqo5AE45cwpeIg8wq9dIw9x7ypMUpPh/8l
2ziPCLqb0LEuAIx5hixZjgaXwBDl5vialLfaCWsqt3jTkOWNFRKDFvEWgjUpICYjv/X6SY8kTzJ1
0M/jMgqM+5XsWnyp7ih533W3mDJaRaqd4KGVAyK2Va++5S1ATB4Agro5f9EDSImqKGJOQsS+U0LC
ll8lsKF/qy10ru3HIpaD/F/XQaH0H4nWzFR0xhbiKVT+lIWymJhWH5F9fCgRInedP8A2JoGJIOOT
oNKeAmQOcn9OU9893BYrQ6Hn1NUfiIE/dKVaiFD7SGCrBHJk1acjqZaU1vuUGAFhGEabC2ulcPSs
aqYAfpmmdbrNKnuK+9fh2C2WTOEniu3rOjQizv0n+yzb9f3RyNb2d+VnD+Ul2EqSN0xqOBJnrpgO
M5gXIwgw/2v9iWzaJRNo+2lxyeVSrMeOR12TJVTRYExya2L0Rlx60rUvzVVvlWUtzfX5hnXQVNcd
v3wtbjIG59O78il2TABCVsWvZ8SFeW26JLjw3cKvBx0OSOF9h4iyrCefiRNWb7OjZSCTeIcumBKU
ju+aaGiPEEPlEce88vaoqiHpjOAIvaM74VYpTEYd/RXxpPsaSezmuKGuw+nnNxIX4S/FbNQvnCUE
o5NAdblS1inzTHG7s314TCV17vcvGyMDYmMNGeeS9/jkZsmtkpcfo2wm4iDFGXNp8SuPL+NBv6V0
uL42acDPBG/5+OjVEyUUyL34mCwWGHNwO4Zms7TSqAq9GqZ1FDGkOPleiPtjVup7kTmqoB5wsWnh
soHDLYYdO7HXG/opOFs7Zp9InFTnI21DpWiovSEky+pIk54AYtzCkyV2sgbcLXejfYRm5QrBUMLR
FqxFRbdLhzq4gktRxhcohbd9eWnCTZJVFQuaTcJtY+uXwNt9uCxDBB6fN7pvMAJN6pw4Cke11WTt
RdRNACQ/raVl9eMyrqCJnqFsusM9p2UYRZDNUjlgFmX8a1e4OyTIMq00gACtS2rQd9LqklvgyUQ/
eA5oKJmD5WuWFD57RYCUipRvtVIvQADDx9km/ckPVBK5u0TZeK6oHqC9dBU6UFl9om6vpESSDh2t
E0iqvSZXq6lVvat9ovBqNId85VciYlG73yjV5uX8Lwvowvh8/iNWOSxudIPLAPwxcOxaDF6mhOOw
A77u4FmdI6ZdjPYOXLtMaW62WXHf0ecg7i0sdLaXM6hA6oHNvKACQ3RmAcElEZkoTSsP94g66mEj
pZjZma7z/l6st3FoCt5ofjQlfpF/LeBikXZh82cVOhRXP2GgZmBMh66DLG3icgLhQAJycmy0mQtO
HDKCWGWoA0ktv/metV5i0SC1iWU9vuZOWRGD9Y5tUaGbj0JXkzu3+lK6mFHML/0b2dNr8XMU7+jm
zHRtTW0ODw70Sj7dX8WF7xzzLgeHEpJAS9iTAbQ6dhbBj42oJ1gn1u6gqrSo9m5abXNQBk//yiON
S5kDO8b/RWOVTNVDd2alQFr+CoW8boWRmjZr6s01j8GyfHFT1VCCc/146EYfMJGQsvnyp0JXIxzQ
LtffAyXztrog69Fh8gko6B30LSKjarZk5VJjAmsCMG6+7nYTxRW0W5TBhAxQB6mm4OG3OxxRJYB1
WNpLKnf1CmDFz/x02zTD0l+E5cbTExJ+1FQ+K4OhDmFgGsi12hOJfNxko608XNh9mKCKQlRZDPaJ
icMGL4ezOUOqvIUSTKRDjQNWQAuYFpwL5dNzrdY1PRZMlG24s6giCJJq15kmjwPkYbRZiL278/Yw
twHdTzlHuBZGUuKVhyc/NxbgFrMkMI+YW3BNy24FRNA0qrMJTpfZRKNa9jx5ztqFPQs4AKnlFGn9
hB2ucFnCwvux9DAVu2IR+RMEg9D3+zHB+f3CyrXqjUsGPwyu+4KeUnuDKuKjjTn+H4eWJXHCeKcK
5VqXFC3ows7/jMHpDiHq1RsXhaW/buMCb7QgQrXfFBT0VsY1m9Rzi5X44n/lqhFeoX2PW9Z9z0PS
Ehbt8SAJpwn6FwVMcQMgwQx3zIvfRcFZHsJu70yWP6U7PEZyY3J/g/mWN65mMlncVqO9TeFPAIdt
diTuMAOT3VjVx2RxtRJC0ZHbqwGCuQUu+CZb2OIYQkqJv/dDYrt3WHzGnrNIOZrqptmWTA/qNlW9
8piGBAxmX96/CtG5jwNpFEkgp9n6O/BU5kfR29G2x4T23WpAWv2/iTgPUR/+DL//U+fhW6zOYWCl
tEbX/2TYL+1zqOg1PIkgaHmDGmo7rAlP90iq5a6K5FSNqBcPat4kyIjhNZErRUc2kpSIOXgsw1El
5jyjpdF5PZVeSbxdZYJ1Q1zb/9bESAR9ydMJrNw6XhigwsRiwn+E/KbUO1W0AuWA4l7Z74fXjo0V
sJOXZ6QURbCgRvGRYYQf0/61FRxk49BujMTe2WmtjEDvv5hmoPTAia89f5dikFtWnF6/WTPiZkWe
TjC7+5JAvy2cEdv+N/GNIzTK/IvMJ6Gafs62pDJJoIL23GznMNNdC9QS9q+R3frc92YrVVNEwWWc
NofOecSnA4RbZG+SP1YAlJCtr9l50p++KDRH+7Sv5G3x/NtxzGYymgttIlLLbDWyQbp5ewZJ1Y0v
SUswI8csrpwue0gPjdl3jKr3Ee/mnUi+MDiHQevvs+9RwUyW8ChLE//XdvsW54UqdpTa14mJm6kA
8JsYq4sw86YCcpYgVIwraLlmpxgcGD5hX0jjCXxqyLFsCfGPwadBQalHW1SlQdESsWaMDIUbLiCM
ieeLonZDk1qECL2djixp3ZiYTQARflJXDS/K46xbNVq08FOTNUhnRJDEfQcdtEL/OQgcU/AbY+CA
SWY0oeF4MZ596G/UGJ7yTHEaRraAR0Pn6bUx3f4wCzmFTMN8RhIpQgo5glAsh6DCAGWv9rHB4vux
vTFfxTIjVJTNDYsZ5FfrwP3eb5/xFJ+WfCB1RcSG3J9R+4bArhEtNpZiFSl1FXlLxSE0D+GFjLD0
nsqxT9XUrx9F68TMKYwEQGhA9fs9k1+s+a+PmE8L9//zJSeoDijGi5djOZS1Mm3H6bQnufyhkRqL
vOOn3zBGBLArdszHktSOWVM/u50F2FuYtBGcwbGRrtEt9cB1MU4d4go+ZETpOHhc+J8Fm6zXmwgk
CUZUdi5WuT8ipE23V6W/dWebfUZjwXz+a67mOIKJvKsDTa03lEVHVpToz4ZGWCsuxuSYoJEHve7z
h5eZhs3us94Znzuh6k1/gUF+JPgpAmtFPSi8hADJVN5JttvU0WhTw84yGHujg7wwIbcteVvK6Cok
HxtTmZzfrXB8yZCgELReh+4iwUfVqK4MoQCWqMuUiinK140OUKqpvFpUxLj9q1IgiYZvhM04OHR8
jCzaski7pe6CRh9HikIXC/wmufvmpKbXXb7R0VDT7ewKQQtnoAYKx9zaFm6t21oicIKOk5N7zjK1
Y1sVrxpJx7bDmuPr1RqwVRaNbFRSp7r5TvZLjPNqUkCKJHM4xOK8l0Zm9hnw4ehIGpZHgbXSq8/X
2qmZ+jud7gwDyAQP+FpPx4twzC8DT71N6GrN5CixQjRrZAd66GRMY+4PIxqhwrJelwWGn0HiqXyu
icVHy6HGVp4VF8t5I3yErG5ImIPLnxkUQU47lPBH3SVzcK+RApVCOYdBvdv6EfjK5yxgcPgVvYN1
tA7Ur99SfhcoCXD0lei7jTR1fBzEv749sB2huyczDbSJA9oZclww44AHAMHUexoR+VZgeV47/kS3
JAHMEnBYNCLBNjBkldtQC/fG4B2EANMV2LiuqqOtPjsE4ZeVIhFEI1dEWaMEkWGg47hS8yzQaezK
Fay/k6VGp8QA7l/82QS3seavZYbGEYAr7v2b+JKF8IosO2gKrhQBYn55dvV+HhqwnefN7wnljhT9
qu62IRm/h5uvSIqxij4niUhNH1Ay78ZVprKuxEUkuN8AZeeqUDr+kn13WQRhyk5nI8Q+dEgPQ5D3
Z0HvzjEit7SsSfYIcLbuBpN8/LsqijNSJydBj7Oi6qyVoS2T0nKLJrudwBqKGu7K/JCle9Eg/Uwa
Q4M++yflrlom6o+R3CXOwXLFlL9tJB5q1vb9LsAC8xyig/VNnykYYBW4qcRpTuS7qq2LCo3cJvQH
oxfO0q3tlxjfoml3mKrZaZ5EYTc7CssA9IrEZ4zkKlenGAYHwRnHsusaxg4fIyGJ76ubhysiwySg
g5uiawx0dZ4l1NAKjHMG5pi0hhuLNNtfl/7muQkcVd3lzaJqfHU6YxMLoHPygQkjuIHyhwud4H2V
z/8p1pm9fuDV9yJVNUMj02zIVf1P7LXhj86C6BARf5da3g0GfolNKqtQTvhq6rbeuwOddU7KVyng
mNHcSaa0Y+3HS9rVbe698iPqvA5Sw/k2oz+J4Ece5Gksd5ZYPKZPTQi61v0WirL65DqR8ua37hjI
Ic9uikkpMnle6T1RDKkCpzXGHcgufW1rgKy0CkJgZZkhyscrsoGP9H7hvZgoYdYko1cASzm5n6Ru
9jWKsf2zrTqx7QOFSL1Ngq07gwPO1++FZAMH2Set8W2IdOZ9+Zl7ebQmjYaC+6X94Fu+ce6yLly/
bQQWOa+v2Ljkde2P51GsVrXX430+23CIy2NjsvkW4cbq2B27ajk+PexRxIsShovHL1zVeyt1tqaZ
H1ir82nY+NEiKYFVl/QWBVaYvf0KP2GcaDWTrMueACQ6/cEVDk7XWWFAYB6zoxI+EIJo968UKBcI
PXxExttw194D5g6GzuAkowYW2iAkDq9HKtd70rTRHMjikRk0SS865nzuAnX8wWiK+bzo7OFMWL0t
Gm3JWS1rTsQAL2lsPIID+JYLAHzdEjdIB0st3Boq9PG+n87HxnYvZnkcL9HyNPTTCOKckVIQ/XyS
YsTkp29slS8SG+IiZ8XVOF+uCn76G5dQYBkv1NwwYGw4DlboNFkmtdChgdRLW92sz0v0ARG63xwU
mnbFltak+QqUk1hfcSRKosGXgZpRoLFnp2akx+6WuKuavMEKyUIeMA9rPGfvZSx3iIaLiuqIrcoG
+AwN9jWIwwxu4sJRbEHcJ2Ype51eryZ0fHszTpzfwxhqyFbKxT8c5bwk7kD/0GAIyb5DGvFYBO7P
DDIYL5PDzgbHZoXqNeA+jL04mdU85l7rn3/9EF7hM3AoPDjUQgbdCcWWjm/JTngKR785AtgJK05H
fyeww8DZfTEU+TdWOemmJf/Z6KKwTksQwsbCsP+m03Jb0CS/98anMxdj3aJDdrveBCECK/xo8GW3
TAFmZqWe3+bqnzKVM4nepD6If+nCUAqPhKca+HReK4AdA0FNPORaYNTgKS6nP96KGydofAAquVgl
rXmgprYagFM7FasoYbtrSXwHPMlpzfiVECAS3nxkDuJvruLc1X3q1gKvnqKPYz9Ymss5/QGXgxDD
lvhb0HGDlDGL6o0Y9vckzQEQt4AdMmXQEbvYI4bmqmaCmAnxsbHnouZG1YxH7OBhWdUZPkYVYQ8g
9LOR6lJIe2xP+7TH7iGyYQlo1kxUHASgovcBmqF/56n0bqeO9SULBhJikvy8TTi+VpkZMQAWxIJL
OqcoZDMrAdJriZJyphkyirvrPkrJR4j2W5Mt3yfEjFkCJunqLIJDlOwZctuLwg78Z5ZgO8NSnBz9
9BUq7geJz5UdbA6xaDh1IFyGpKo76cpD/yBW/4xhJDQSEmIr+qa9cF9uOov4PcIaXCCZ7mFLrdsx
jOedHqvI/O2qZbKFyhLsIbB9AIW3FrxTI/3/bzxlbJYGyDAxHvnhZW+XQV2rXECYmwBGkDXKmE6L
mY3u1nlkUD+LSM1P1oE0kMaBqPU455r36TyWqQI/Rjg7XQwePXXFGbEe4D71N4g5YjoL/Gxw+P+j
PpBNCko9CHJPOd6lM6XxiwyH35WkgaozVAFjH0kpFM+OIa7P4aXlumZfhcptOHwx+MJipPR6II45
gyr48qJHjt01OxWk1vWw6liYkYEJDxYnBRgNAbdlRb69tcFEf4isPtR3kO8LNj8NSwx4KHlqj2fS
rf9mW07ozf8eQjVzZx6YkxzWvrHHgzB2cUT33XHAGGXXkxKuYG6HGjvVqNGluNOvLXx8O7Ddl01H
EYqBTxo5oXZJnYeIdIljVAdoC/P/qhJ6wTrFN+yhjmRi8Z8hQY0nsSW8d8M+Lpwz/bT83VT7wpDq
F+BYeDgCH0A1HtAVaZrUXkNj9eJf0fMq9b/TgbJtRKG8qi2inXE1kE7rPw0j1Vj7xPJERKogYIMe
aUlEs37R/cPWuj4HGZeL4T7glP1WaP8EuF5KUjkmj711DPuS4XgUEoTzRpC4gsxqytgjpKIDhvME
YuumnAMef+T6KK2F0EQAFIqjatROtPVH+r/yzNmTQln6GCxqvWzm7itn69NFoCc2F/zqnE90NKi/
lBH7yrJi/xaUVlLQZR8etGL4mcnwy/WvXxW6dnFIgVmiEuqAisJocBxrSPRaI1ykfTKWtSq/I2oJ
2s41O7tQQOx8M5CDEkKgGPkGkCmSPNeImli0Bw1t9OIIMMpgdYan0Yjs0hpNzBxVptxm2/2svPeV
YcF7YBk+PEHh3A5nsEmoCILeDLDN3itGx1KQwzC9AneoMTEOhRZXjtPMuecbdAq9RJeJYRx7c7Bw
CdjdknInwNc5RNW81BoCGryhypujBo8NOExik+l/dIiPgaghl5SPrGphemsM69Y29SZuN06oiTEZ
pz9X5reyJp+2qGr1+HUBO2RcaSQzUNHpjryfQQr6NA8ehh2IyhnRCK6DEBJ5KrVL8rTzgyi07tRN
WWm2QCn7gHgotISWBGkIz6vxyCU0QByDYaB7TfyS61lrIiqQYE5P7DJV9bp2tjWfcik4lSHGrkG+
+KZUpP6ho6o9w9kJpDsygnDOCsTwytRBcoTrv5HXJm6X8EqWs/DFZhdxPvdPl3++BzC8COXp6LRQ
uVH0zT6KQUOOwUgT21tvGljgj7XLc1PfstaX9/7rN9BxrwmJwagIiLcIh8ZqtFHIHCwrr1Knoazr
+JqvVvgzQ2FcayNpJzQWVJH/QkzQG8mLFonVWPNic7iA9BHJknHjnm8l9ooFd5OwyVA1EjPy/lOb
L4ZkGA1ui2z3M/d5cs0oBVTrLOFJ9bvhWa0ZJh09R7xsvhfezqUimMjyBb5VRNlCor3x9u61I7DA
1polZyzgcJtEMe/kAiR3HJ7gPuJveSYu2hZYQbDCKTlB9wa+fHvba2U9Da2w9iBK/9TCgwqejrN4
A2CPwZi6lwbqkDCtYGjRVx2rmUBa9dAmaFu00/Sc0uhtXBQUA09Wnf9YvxB1Yh6nzjf9QR16D0Dr
yVYTgm7AnYWWgnuvEglLzkAEZg4v+IaqRizKCbSYpi7cAAZ6z3MJpo1ppWZ9G4So1LwLUf/J+5C7
FVELj21/i8faSOCowpr7z4cPKAqtuT+chnvTfpcXUoQO4xF0esY9I2/mHSy4l5g72HxmtE2Y5+Ac
g3XuzqEJLavm6Ikv8P45EkNpb4C/xPbp2uiqT/TbPcN1bIxcd4CyStjX4W4nUCrbrsJ4C5q249Cd
6OIoZIUjgyZVmUE9hVdsQO2B65JYfoG6eWKmiisOU1siRRybTnmxWXPeY0zdxvAib8fD/QmY/Dkr
fMbSCXogaoPztceYwUkgjCmSf7knvGj0tBvpByuPSSE1nu2X+hSSKPEKb0PNMSdWXUlWr7rBvMDT
sXo+7ORuhzchrPswXJVqqEXQdmJhQxrvdOA3dygfpG1EAtwV8qkKG9b58PEfCX1T+IOtxSzMg1ew
dXRDA5rDu1TbDV3pskhPqlizwQ3gX1Z+twr3w9aGlz+A18egY57ice9QP8DvbkWttL3EcQlxCgSl
uLHVVDad6KG9U6QQmzXkZIX7y9c2OO5+VzFUYqRF8/p2KNxscj6EkqpSYt3+dPjPYWcOrR5D+1cM
AvAT1NwSY6aBPHCLE6zdFy4JjabfL2MPOLCyudj9hWlWv5niiXpVj8o8ti/P5tskeJIpT+qpXLuw
T3IIUnP9ya6q/cupbcrFajC+3cx22VAQBKeKdZf7AhaZDqBUJeeZbuGl4KSmIs8G8FccPPNAJykd
gls4hvNeCn+aiAL41McA+2yY/mw517ITpSs5jY4RlQtZXHcqc7KNFrTD+9HGJVzEWQ5qhbWlY1M7
pdSOT+mRnA1Jpsyo4/+RlTk0QMP01xhdpZ3aYd0pm5sBXDUul0Gjzt5gbCoPGaeXcB0ovg232n8J
n1v8mp+TRVeSEnC9+Y6xjdbOpBpFY3fGFKKlCr9WQCTicNRJLXcThcLq5PloyQ/BtmiCMbftZ13l
8c2Q7iAfDPOE2hglZhSc1cadhAOs9kityTnpPvcfSwtFFDCsCbF5OMXC1BX2om8+kUQGq7S9XWtc
NtLvAdlItQ/ko6Cu2spAuVDkf2+Pgei4l2H0rwar9h6Dj8UsFYL1vwXoRDtLVLIRNgXp4sMLsNH4
5l2IBh+rmv7mphQt8NJ/x802GLO72hIr6DA2b1PMOQneGvz5GQyJf+COZW74W/oawTWfxQgvRbHS
RB8pjTdZtIHzgnd6Npi6RD126In8fv3k011th93XwH+04yWyAdEDOf2pfEpNRhhKcwSzbuYsh5BR
xyuBCAWJsvPTI/DbzjLny7WyJUKRobMb9V7G/IbOYhaTd8CLKim9Sx3iJqEqSezWfZZ2J3z2XTcn
nmF+x+RywisAwWi49VbImv1ZczXGDCOVHNj3ZT2hbYOUvANIVYCgbRidbnE47RJuIJNI7OXns/CA
5EoMKI4p/p2fwsmUH16Jju6RgwRcDvqqegVbj2qhwElHQzGaGYzL3Rk0roaWEwjq3OVk+Sn3faM7
m8Uq4TnoLk1/yV5fQwbOJ/BUzOEvPzO7JBh3WrlHAYyV5P/2WmnKAIWr8WxMz/FLdIRo+VDZ/6dl
zpH8wP5b3kQALnjbrWXLgVzVGGUAO6EXg1NzLQLvGC7h4uUkvtUk4/db9pC65F5km9ijjSEx7uDx
jEUgeSqOhH03MCVNl5oryxal8ALTkeJqw94WZy62CYZzB45qh0g3JyjdF529CcWniH9pH4h107TA
ybBT36qM+L0P2jsM3KO9Ow/apoSqJ0I6uFvMduOB0eQpaAKy0LKgszhZbiFK0IluCKs1CmhzL5yO
KBo4jSwo8mEouqe/zHM3uatMEb64ZP1pUXOLJucyiDpzBlg5iC1Q73y6I43IfoZqj860I5wy9Am0
A9g137nuig4nlLcPtAMGoluT+iL7Lh3imsSHWNJXHU8celHTzDj99EZOjbmLlBXCdqL5T4Ea+6/7
j79d0fKduWzTw7SHa4/NEkiurYkrvtb4Z8FRPtyBSOwxiRrazy5EhGjnF5+hVtpjf8X+lzrQtHyU
DZO8RfHsJ0rCr5ku9SIvc/3VxGq7saR63IxWQjeL049arupKQ8pBvvBeM+ZubgJdaO+ZeWDaCuAl
Hc2nfzwX9ZNsvvBqvC8pZBZiO1JIKJnDaee7HQq8ln5N/vV4cLMyw76ia5imlDU6KI0NP5D9j7sV
VN2fbZukg1y6DGv49yrfkibkrw49nfUDZ2IpgMbQc4+kh2r+pYvg3ZEJIHiWPVchTQj6X6yK6Sz6
tOdW11987zLxV3joZwGqJJ96yzIMlmdu6FWCzlAYmQwVUzBzXpDeTfZ9rO4NbIua4VoSbXXzeWjT
uSn12pIRBEaW580O0hbATOSfwqLHU/keU9WCNQeERGzhB3X7z6vuFjLGMT0NV4Dryw+o1XlwfrSS
pWZXsPJnFKFvVXt7AL8EHQYTrYTCAJO1ASBHrTgyfh4hl9TRGvhdBanUFUajMEd8X/NG00FcPO1j
xNGVFDRBK30U8VBFrHFzlr6XwTlY3biq80fagh9EFhE1rwhzxOyPso6yk09GnhNdekiRTmKoDbRT
pLTA8E+Aek1bLu0DE1y1a44EeVYsVLSyZ6IJn5VMnMp1xfY6pvudJ7s/9FE7lKhpCpk7s4RgbG47
7s/yF/oSd+nlH9U3IuDXBsSPfLX6jEYvd4E14rqq5bcaLdEPjmjF1LRdKb0P4aTJkSZdQ/7gxwfD
v72xCRt6fvpgWbnT+/x2owUGi/bLzfeexGXnzUgpp9Y1ehXTUzn12vp58wIKkkF1yrSHNLa1FfDt
BuRs5ia6rC9jx+02U5UIMsNbOlfG1FDI6W62FoggDV5zEIwBAAfKgRxEyILwHHRvOykuyKSOry7e
427T85rFYnOheesJvOaz63M+4n/bcmx5rL8vYbo20lNX9OozkHAg7fpg93gkAot7qb4E2jMnEv/r
zgPdEdCVZVEhU8a2huhlGxoHn28Pn+FLvHjOet6ZQKAx7/wurQjIrJxgc1wOV3YdYJCnRAYHp7Po
6vYGDUY2iuvGNck9/iM+LdQD/9AZba46r2WpqUoi/Cc1lElHDKhpBMAm3nDrFChH6af6x93/KBcR
fNIprNISKgkeSBOfzazYA+/qCecVdgDmSNM8SPQqFzoO4tfjdDuSVjwmzf4t5mYeDe9wuCog1P0i
gKZoIvWUOkYNebzNS4HshTtkxeYUaaWWT/3qPi5daXN9AocBbJuxHGqk1BIwczF68YZXKkJi32ss
AIZjWhVQCvzrKBFDJFh2Ii77d7sKELsKANWleiCVTQr+bVthyzRONcQdnYW0tsSAsynX8DAo0Hr0
y4/u8xRp/078WISM9v4mHvbfuT8M1y5vZu3sSdkDgLdWapquJhSRB7NKeFVW4W19ySvjQrOA6Wkn
JepmIJ1RTnC4UQZpQKbi7hk7DvvJKSx4YLadUKpz5VM+KuF6Tr32XcR36//Qe5+SdGEzo834ndV7
UrW450r7O4Q8XQ+5gH7avuH4cVGEUcJa9JKOJnjsbi1xK7NxFSax/hBANA1YORlDPbyVlJqyliZK
rN0s6GR28O/E/O8CVWXPectUVzWQ7SRyU7Yn0cEF/2Q2xryaJiXo+8eQjzMggjxk/kyVSG1FolOB
Toetjju9Z0dzu3QkNKxydoBvEuxVvQ04IIe5STmvz4i5Sw6hiFzDjN4KqmnUQQdQRUPmYTiV2LGe
Gqt2aon0agFHa8s88IHkXwfWftuja493K/o5MjcxVVTG1ii633IXEUhyo1RN2mJZkY1CL1iJASC5
ITXIaTrfemGSflizTWCiaQwuRimYEuoFEWRC8HMsrdaviysOJ8QzOW5XCK1daxYNcHdH/JPveRXQ
l48KS2pwOtRPC008GWEQ7QpmMUPAvcj9QJJ99AWXpmtU1Ge4DnUzB/MxGndpvYFeNzdig0l4si34
HptqoC94FL4rBBPE77UXFVUG2gXJxkUs90AkxoxEBHJNmVqHTOVsviQNFIuKjvkjlqpv1klfViKy
BUNf5512C/WpHupKLmkiG3LM+/OkvzxcGcEBbq4SCVzCUnLQ3TGyekz8zQR2D1YVFtCx5RL78U1C
9X2ICiLuYzsdBJ0cQcEXixw4QfQHSbSkPfP9wRdlyRsTSjl9PTGsXehsmB9f8OsUpuAR6jULauS6
MuImLZOi+3zs8Mm4T862wPAdixBYuKeJLOgL9jQWoALeCZHyueMXODfGW0r6gmHw+BFBj3I+uR/U
kGxvbk5jIBpVG0krOaTuOY+ocgU4rmwFVACoG8I/v0Tq/YI11roOl2kwDotBEK53Ms8EWXEoiCDx
AZ6EdX2gFK0jMOZt7bLT58WdKXNsIYG9TVqQ9OcpRpXD8m67SchH4ekLTFNXa5in/vRe6THrrhcd
GnCsADkKKU60BEFkX64Tr0RGhXINWlpjAdG3VhsD+8nFymHq6vx+JKfNX8NrHTFPzQ3mYneCtYdf
97P5oX1O4bxWvzkDNKnT0mmP6AP0w58X5xZgC6c/Tmid+kx0/q4p0DEHC/hfoOWC+mTr/5sUuLvb
YK3EjPRzBD2n6wIlpD6Fl0sLT0ZlHYwc3U17Cd2kqh8ZaUyLCDawJFR7XsYcqGWVlSFOK3JyK0Ni
9Vlh1nc6WPwk7nYhrf9V9xQc23W+4o3QTSUwLCP5QrzZVh0tPxu1taAExWVmR7YaB4kP1jVgMPKE
X7mh29/2jL5ogfMea+6KtUzMBRAJ6i3j0PgZtIj94QhsUIUoMurJm7C38tFP6gI6l0MYjAG+9Mda
JDC3v5k7JvY5k1sEzo5FrMVVvw11wOMT8VEpV3RH5zC3HRhBeWgWxs+jV5rU3ogvU0lfH6ZB+8at
sEAr2QbnQL99r5dyhICj59jgwZmIdNB1dY9JR5P63496zTxNvlTJEz8o4kPtLTx7Jywu4TrcOxHK
cqxgv3cAfgbk60cx1B203b6/+AP8zz9KG7HglUpljMEOkY26cvQ3NT6h9lWH14MsmdKCwzk9Ilow
vvnveW9puOi/mTNrEZlKE8jvDnLnpqKLlfObKf9lqSWgE0w+h0/OXMnUCLG2Q50G5/vJExJYHJmG
WuHa9KLNntJAdCpsbXbpPp18jBKJSA3hxMPQnJsuRZRA4rlmgil//L1W3fLlLrOyIjER7HOCFib8
Hk3XQXqbgi9JjpC0yVhKgSX+nXunLndz+YLdhBZiQD+THa6b/UmfHBDpHOxHthOcOF72Hre47K2f
6ZALXXb5KXzDAlicJv7YaTpkYlwSRsLmxgWNHKU+U4xGEg7HtRvO9rNNDRGGK6DV0mncxkWBevM4
V2TNgENxIoTjHcJFW+F234dTgg1ZphsQ+zmPEVpWGbpa9Ip6y0jO39VnS5+ZrBKcicX3glPbdZ7J
YcgWng95Bl6KEOhhfJ0rX5TpLh4gE4yDVJR4dpP1VNa8Bcx1C87jIYL+4i2/ULzOnv5/9J9QVsoK
QtdQZCP4aIN2M1ZD/mhaDw2K3jmuoAJSd6mBQ5rDXSwfbC2B/TFg1Kn6gfudRPi8xwfklnWwu27k
2BMXFx11P/AqnUTipMyM3wK7w5F81y9BIubWqfd9vFA5IBuw64Y+zZ+toRCzzhorxsRbdVZF2pnd
Et/0bGD6YyiobbAvB0vpGDTgLlqk8tt7zWJb9z7WGYrgNYmMBRUUGQdLX8t/OPsmY7S/ToGAknPa
nHXYDhuELgv2HljKOUluI718WNEHrtl/gWmpYJBJrD/lUGii4f66FAHUMPWoDiTaiHTAV2UjWq3w
Tr5LIBOR8BwgvTAH0llHfzJcZwNAOGlFXqkKhBFOJVLOu6VPiXPAD79ecoEg33Q/IeBdQ+Cshsmq
HHSr7brwbBvFLFi4XR71Kpyi0/7vYPHGgIMDV8ZQc1Ho2Oa4/F7rzpH7Uytio9Bcck2e317T5ytO
Qq7ihne412Qi95iQMo7zN4MZvnFR5DxzW2zYb0BEHlBYJ6WGnRgNlUuH5e777Z9Gf4R92fgXrkZI
Za1RVv2/3CbLOCf6MS7UCkA299KpK9Bz7j19In0xVJRlK/MbzLigjkdk1VcGRmV+tRbqbAQc+zmw
jPUeDCmP1axoqepqeCRlxUPpyQs9i8DO8HPtCr2mPuWXFp1Hib94do66gNssCl2l2qUnhv9YwBKC
AJ3TLwMGV53hqD/DjUieWNRxHS6jCxEVbgZqCRCx6zhpCrt81KA3wmgSDPRMApsNsOn8y3wlnq3I
QFfMov1ZsK6kxIu9cEpJGoC2OUVIviReLFmMjXzqh1/0bRpVMlXX4GPFWtE8AkkzKJefo02fE81M
/K8SkWboe8Bj3dU+4GNyerMtdPssFqpbbn3wicL9qgmD2bA1cduCEL/Sg1xtsdF5Zl/XTJAH+SOu
9jQeIg8qeY1QGM857VHFc2YG2d4ViV2nFUBU1qaOOJ7eBwWgNq0Dwhcef0z7RJJsQCna8z/PdpT4
Tu2b37Kzoh7UDbSPmCEV3dZyY2aFkrDuNNsg8gqIhDZCflz11wSMj6DEfMe0bawAHBVaFKXT6JCZ
z5/9uaLAIusAmFt/S7eaYt8zrZBIJ/RhNw1O5SFnijNDVffk6SDrijLfHpisbMsU9+3GSlEBuXLi
B2WR2YAkrHFunJRMciNgYHZe3W+tPd4jYrRLK/Q4fH63+Tw96V2Nv/oL0WqZhw2gm2sMnsgykIoi
1E1lG4E68q5Zg3fG3+Rgk7yJxTCE8cnzhjNMWPt45h+oF+QWf9YTm8M36wODIxgO6lj0Bk3x42WS
K1uCzPiGkB6ncwB4IBWBJa/Ll2qHXP9XOtnaC+k63nJEtAvR9ry6L2r/i961BKKiSeaYQd8+cYX2
4G8FUEcrH+cOTsySvs7BiSILgvgXuoVh4lDPplaEgrOknwB6R/VIjgthJXS4crgWmySdVFhy8RIz
R9BvkMyZybHqdNgltDZWWgY+Yuh2F6OAFN7OB8MlHvn37ezcVpqFjMzaYqw9cp6dH0fM9i3tgSNc
qtzqf4atjUF7RRKWRtUxUcyJX0XF1ZeWQhQwm8kCbObJhFlcAVH1+STXt28uK9AjIf1uYxIiWezF
5vz3hGjjI3HSRoYaAunPTmuUx0vLU2C1qK2gqdYTBgqtVpRM22huHoMii1vd0qvrACH88RWzKlT2
+MrCCALqgY0bvPOlykddsF3QF2VZYDgijw/BIjywQITpgnnWVhAwP7/YJ/oWzHhTlc42wnnpO4Yl
ibboLY0R8HDa+m1MqDgmdbbPJBs+zOd0RJFdyaRNxPxPVym/E0pJ1OPSoOyxqfh1KKDg2eYdwCPi
hUPxSJI73lSy4RoIRGVl7oVoRcrOcbfX9HqRVQs9ITBr+idtveq96nvC7k6oLLrGNTS60Z/Aonxv
rgVxKn3fLfXz39/Pa3UQKqpk9H+IQVChu2Nj5rnyjj7KKGxsOA1Ogn0qAAhoTRjLSTZEFP5h7Beh
H6Kkfilj2q0tJIvgN4g6hVyQSWXTKYOrljGUOh9AafdLySC0CLJI7Dac9qftR5Auke61UOs/Vwcj
LNfGBiU9Z86H3rxwrDo2OjV/nTzpoFChzLqJZ/m6L8B2SlnkNO9BnfEJeGH9tA5unfiIJ91y63D9
Y7JmkJpadqpetpXm/pnDEQf90j/OObrjtIxfkHdfzmb7OvWvhthW6WDZkJHymR88djJpAQxA3sbW
iqWiGFNDJCtVHMaCtioU7/pJ7+0X92J/BjwDSAL1dFMY+t4b6yAqFXSGNVaD5oQfP2L8zJV51Mzd
D/UPPwPm538PuAzXI9mWULq98jSXkagxiZZGkDKsOMbE9cQ7YNtC0QTQl4G65tRdyI8F21FGOPlS
ZrrRKn0+eisCSzrv/AV3QCkjV6H44Af18oL2kCA7/Iw05ABv019GvABZpjqu+cqiK67ePQ4uMqX9
X2RSiA02fAdydLk21qfjB5ZwdffJMyS8xdx5c8cDvABTCJ7z/rhKdsnIhzCIwJsP3jw3EXNeZYsc
GP8oSZs6izhFNzBWBEXAPoQyTdgHLMiSAGeNRTRDoeTbYyP4nVgFWi44DJDzVerH0ac2JteTC9+i
UBFZemgayFrWphPbAbMOwlO9UXHwJQLJaMbsfiOB5dC8kqCexkt+JaRRh0j+2KB19ATiNmhhcTrI
W/OeZtHCoz90lUy1TBc4mDY84iudB2lezjVAHm6z3X4Nuf8XSiwoRtJB6nWHEpQuO64prWuu/1xn
i3rohckKttKHdwwFqQoqQQ/cwnXmBrwQa7Ijp7YFqJT9CEvcdGmpfTNS04xxc4rdjKywDddsd9RY
FMxDSAZfuzrHc+p8aWLj9AzFdOiQT7mWm2liWy6qtOEiOoHLFXM/8X8Fmal4PRukpIB55a5oPLy5
7j9mgPpAXlT2bguHov03F3JWp7Dgz+ao/K1v4+wHHFFLHBtFxZ26lAveMt9kKKm8Fo1QR9Lv0uyM
ATqq2WgC54kQNyhDroU6wOOP03XRo9xUuNtTYe/rH3U0O27VNYuQrO63HzjmCeX+4sdqfd1GVdY2
K3KSdjGdX4N8ACqiH0q36Q7qny5HZjPqByS2VotStAvhTyiuGyonNkbQ5s8dQfn5y3IUwENxh/f3
t+KZamx1JI+5PRE3Bu89avJHrCwloHcgNQnORxCfaIgxEzfYNfjYYSNv10YymLi0/vWGrvsdDMNh
mOtCviWxkpll3fWHjvMpk4VZ9pSAf0j9waWwBVfNvr9ihj2rq/oKLnbKiht97gawj63i4qVOwlAp
3ElasXAhnqTHrLIEAok5ijLRFTe4Sca2+NsfW6licsoRGixPku3W/MxrO+NtsrBiKQLZLFcxr7Ih
0kGyLizNmhWcN4tSy+eC96gA6HlEi5eL2JEv6M5Bx2HkXW5o5aPzoY2Gpdx3zST4mPI/m51q9ssw
bv11TkBXwBWeaFwVvMvfcms40Y8wwhnW0cHsrtKqUsF1iBA/ksFUPVoXPm1m8hz3D4tFtJAjxeXp
xna3VV53+J970WdzaY2RHcTZiZoYTjhbMDy7K4b9nAwZW08LWco55jweRbsvJnHiI0aVsBo1HAoT
MYe4/l4Qzu3rgdgraH3TmYSIv3e6OQpluaT5UlIisJyHUknLaQ264ANfiAkjQU6XTeIp3LYSLKeH
8k6EbmMpArYmVuF/kxJhV6EYDnrJZbv9gQKMAqZR+Cl8XlMuaBy1dE42vk9/tigHJKMqg629nmho
YFK3wzHL/1MRnGUQ0E7Eo6su+clJWT4JRGLlGbTDhQFyuCnMT588zftGnW8pFpay27y9UA+if3s6
G/r0iMdrcf1RN3YsOaLlh2gRZyR4ELXi9Khuq98kQF7PcV5M7/9ohqipuCVFbAXuMDQ7Ms+0Jkl8
rAXJ/RFpYOGmfv1lJjq9t3Skw44a60iGdp/wsO+6o1qRa++LpzzJJFm//s22oXBU5xFxap0gOdud
PnAo67xVwMsbSYaXrJy6d0GbOCdazA81eLgjOxPfTPVs+//IZkNGoW0/ib7XQexVnC8WpbgluNLJ
1wqcYNQ5L1YjVTajUw9Fk8zyYPICBsSJQUMVlLS0scAGD5LrwV08u/nzMXGP5Ja+4wh6cSAQhciV
KKtai4m5yIiOGUUrskXJECdltjeimW91FoimwIXItZSDNvCxn275IiRre346K4MbT3+lFvQqme6X
Og+64utlHg7eaZa5+S+qEukQPst1S9S4abQf9yIRPjcy4HO0FQC04d5lXIWPeYAMWWwXUnGNbroe
lTvgVuihk7zqNluDCD8h0b0Yqlurn+VHNu8e8mGiqubstrFMMr23I7QZ/di2Umw1aWkVR8PktFF9
2WYExGa5wjUbog3bWwgRIWMZnhoPTzji0JJvrSYyEYcGnPBqWjf+s5v0ZQ/YFk61mTf5PW5YGYah
wBIm41Yn0Cik426Jh7bwJqbiDd8PTOZsGZ1OQhEMMfRjJq5XcSnz1UVw4OOnkjrHTUb4WzwZ0sBs
lCByRM8NVJF4Jh86e6tkWR6N7390TCVJTn4ujwwer+bhvSQayGD/XwWhVCkBCz1El/OZHEWlUf4Z
tdCFBjuuleQ4y0QfshKBIjXfqnJAQ2j10RxLyZrlh1TLF26hSbLpYP26TbGMBwvjpzC31/gLpFCQ
in7kfg6Qw45vp/Mqwg1082woEZTQkUJEzvjzDfgnyVXtvFoPnRjsA0E5Jf91oFpGsfJG9aIhgtBj
+UqeRgf4SHFf3THOEhxgQ0MegDRXtdSBvjxlzSRj1qsXDUrRWFYyXEUvlmKRk9UOzdHS6I/UlFm0
pFlP9rDjl7ZqIXF4CGBKJSJHfmMgH+awyKH73Zmmgf6iDUPZ0BsKlx9xXc57p0dNnSKFuQWaQUhO
E5h/XoJ45FBuAp4nSeSQ5+rwYeyd97WWAVRwni4Zs3ItyKE9SIqgTB5K66Y7cSn2R0lRITwDlpy8
gVP9v1ysUcQhixBeoBhv4PmZbLFDC28znh4rhabYOk8Wzwcg+38f72+SS117Uox5b8ap0er8vlWR
G0ECd4JMd3mK/4WaknGvhX8vvMjtDZmWsnukCBASVmt9iZSrWMVetZISG/mg2VCzWMIUKl+z9r0M
6uQ2O131ahjK0LCVUofMKO3+hDM0YP+7Ewqk6ANtNEM+WdWrIYA5U2ZV9i4LBaVbMEgZXRt9/srf
PnnuqfcGgswW1o35JzXuri3LIJt9u9Z0g+sDNEH0aFMCuHxjccaeHuRy7OLeHHhzC0ypvXJbjpZt
b+qmOj9rGnwEIyvRv8kl072/zZP3v2ZpBPOy7VknR3ntFPdzH3GcFr4VBWG/habmSrAzZB2G/EY5
0xUKYC3/bMIW2TOB9ruuaoMIKEhg5tJZOw6q3mtrDvCVpaXVXTXWCjUNo1i8gYO4YLp4esvYtVgG
3LbRlqCAgIN3iDXwTI2e7GTt+afhzdixK/YYIFsWDHAYCpBOTpFa8BUF6zeZca8TGDt/qOs0JMFa
O8WQlo/uz1dvLAhX1cIYl8ZWhaNewzZXZz/xjNJnX28gV+JfInr7+3lgHftO72P5LCLhO4Kx/SnG
1zhgIVpChsnHdvdJv+sxt+lb3Fm7D4RQVlkqLaQogb2uki24tHBRVNzYwL0izbWcLYIb9pq5ZMBP
cgF1nsQKDCewxlnH42W+B6mKrN0niwAwcW3z/Y8WowNXwXwPe7pbqzzU+OrlpZ5tifdgWcxA+BRO
jMAev+0aqyA8C65Gafq81cOYVDbKxzZoRpyWeHqFW9mQ7Txje8GtrqxiA0Tx+SDg4xJeuR/7GkQd
Rv8rQlBz0/aREwCz85SzIJ8h/eoG15VFpHLlz92n9Ev+fYEd5xD7OZkMXPnOgwH90I6kAXML9LCR
WjmqZTftjAEHuEMQHXTY2aewa3o+bdy/n+SGysOUjh8G5b5whBEyqn/TKhKF4oKtz54KqDtCXzdP
qSggvZr3jj+Op6+vtnzZzVXG9UYg5+35GFJfIE/cRGD/9vn6YR6f+ckG6HokAW0E0hwGjfojEeqi
nOdI7rmRcdBSTlSqDk9yXe144tz5fMZHmwQ0XXGL6Qm2OCjl3fUyhHBvJKSA5EdcWAJX4hawMyTG
3lCcxU4/Y3Y3OPGQ/f8PYDYt7S+El10Qjoclgt6GpJeMmOkWGE4QxeM2W6jfZzzgtELZVnhMgg23
wGJ6wCYWvFTZNTSgxnerqMviXub5didgWFtzhLFzAMW13AWX/iquMQI8vzVvUarvyRV0eTv3MIQu
vEEh5PIc4tL/6xXV6igdTQx/I+f8fSLQZWHZlx33ilCHhphtonWhH8iLZMjteerfzYk6Fi/Y2Ag+
GHdV7r15cigMrxKmbZJMEagyehGU9eiGlk93YPbK6ucgghELGaQ0tZnp4kQw1vAsGJxy7YW3laSI
qqUz+QInOCYZ7DH5KUhM3pggZL4i9NcBPgZasW89p8EMhjD4rinCl+GgKYBdjIbJV2wfByvY+GDB
wEsIa5MjvNLA16Q3AIv8CmX6nlKMJ4nKBjN2nAh1o03Ru6G0PbB2PKNgB3E/0HX9xA7bS4CO3VK+
DvMaBPa9LgT9F5a3Lfo/aX551HgnFLrlJpsbpG2sTVxRwppt5dVEJJo75HpW/1QMzUcsio/AF9YF
h+Ekpm8v3rjFJJBu3m+Vb8gJkYPOGlS0E+F3PuFNtPtoxBBGu8trPYvLPUbJMGOScPrc8Fd9oDmz
SQ2FlQy7m3vg43JaXRWmAoNeYMai2LsZ/5oxWemKnlMEZy3tq5YD6meLEXMwP1AvE3FAIFMiRwJH
sAwayRbeKecYbk7FS5SD4H4LI6NsVpGoix403qMptXeRp5bsxgKjNCPTq8bMWXUJKHYaHNtL1mEs
pnxA2Kh38XD2zPo3fEhTGGq/dj6mWiANmmcC9eJjUcTLuzFUcu5/AJDz0180rxZ2QXdU4HyeScL9
d2I5ntA9Y31FT+RY2rL/tm0ly3sJ/owTyB8U/f9utCslF6ed5JR02M8OuacjfRsIzzxZ9f1NPdUV
MpVbg0rt86yMoQIA9L7ZBVSei89KVApzqKCMs5Dlu4n2v2O6Qr8KH14BbFZQ59xO852zF1dVtJ1C
rhcx8t+LNNxfr+BitJ2GtFabuaKhA2dUhUOpiwSRcdGmsYJQb2DFgAl9VYPvZJn64IoAcC1gambl
/2aKyTeO+kYyZn+ziIOw5cIdxdohEuu920e5gEuDZtFiHh5+XWrxQhErG7Edo/0enNSEUP5zhYEg
oiyBv4REBTDgq4YXlthNgqM2xkpqsoY02ZOqi3y9a/s5ySzSNzWNkrLV+xdbSoLh0pUZUqUVD5+U
MhSq5fs9ADRJ3UlGNxnoY8pLYAZOt+BQjIVbN7kXMR9HUvkWi3GygKAOfzstuVzq4VtVPJMsj/Aq
FAgTFFUZhCYFkf+7jXKU1z8iwfHz9G5e7DjPHoEenqOZmaB6HdEx3Dw6Ny/cce3eRplLwRF2Rny6
JoNdY/3SfV2QkwXUCh6S7Gju8JfwwG8KutPz8gPT6b4VBFKe+MsHtx1FTZagzI+hqf+Nrq3/BlSD
/truBGl27QTDrxaij5+meKACxZ9uKWQ5Ox6VTFMMDX3RnI78UffuZwi0fV2DKlLsbQBALXnbPQ99
Of64cODWzGdLp/HjNms2IvbPPnN3rBDNENILmmWOEz62/0y1mgt7tP64OPYz8w1Ionytmx7QtaaC
4kZHoCGvgcDlFOCjCMrZlvilrzPIoV5DmVreQQMH2Ebd98BM5p50sNVPz9XmiaSm1HNsF7qgv5FU
0qi2/aVjDFSd7QDk/j5gkcH1rSGOrlj8mtSRmGXRe5sFW2UotO9LWeBcGyHz8AU5OZj4nivsNfLq
OpQvrVH2qPanyreGt/zkBbEyeIpjV8YOiDRj280ZXI8oOJOBu+CRwDTsBRWOfaYmOOFLPYwJr68j
6nfFoDV1c8E7QMSvNIAoNFQQQDwaIQWwlP3RyHpiUl/566Qpnpq/QdFnReSosCH1EwkOMjS7PaOL
KtIs/bvv++6+8+KK21DAFLUQ3n4cI3jWkPiaOUDSW4D1Hx/Q1XNPUeiCL8AUgJiD+dQw05jnXi2g
Q0Gkp6ffcBeNiiHrLZpeIBkcAKkUlIHGsdrba902g1sbu4t4btMAELYCk8Gc9c/M/0EyqWNbIVOl
lnoIdqUtn0KtOxEDuX7rW+gAi29umgT7IVTQ8CQDK06ujJChZ9jgL1NIO6FN2MJs9eKf9ThpMBvm
oQ7ABIJxiUwJKbOvcsVtCneA7ahIhhhor1xa6q32jFnaXGDx3dViuD7QzfHfHrDswJ5Nt9vwIUYx
VvNq5qW4vgwShEAlv5pL1cATOwgSFmw2ctK3Uw6hOLHPCNOSoF2d3ZO4G8Np6YBhxfw28oWpVqNK
gGjAJ9HOZRaN9aIrkGD8wQ+PF3iLdaC99gMNcXsD6F+K0PvwqmCoKw+H5DwW2ZDR+/N7OCLISR9A
MMdUdBT8U1Pfko2RQGllVbx6ule9eApnFCG8PJxpqX/ZZfdHSr5EjeZI52nfa018o5fyWiq2n2nf
lV1oN//kms1C0qO9vJxpw4XVwcNSXsB2lp7kFMAhomLt5kGNWcHDA18+mnyJQp4PyFtA0RWcPlth
V4nTMAZSoTfmN3HEBkG9hTqWvuj8Lw9PAzp5MdKKmgNUYm2inI3PFQTO0mhA9cKU02rYNhIiWKuw
C66qzN9Dy2vkZXjfznkB/lTVholLOI79dVMlPwSGP2OsZZnV/3Qlafz04LQLj2Y7Uqs95IPCR6Vc
vlbTgDXfid1IahLXRucFfN5yqo1BH7xBE/PHMaN40KGeqte52TzfSZ6PpZcZLKrzWHZKWqGwZvcU
DZEGP/Rkn2nArKRsKfYSpKy8xprBxkhO5N5mV3IElUS50YSBrTQiuxYJggWD+UMULghTy/ldxoJM
cHNYEtqgWHUe3JX64Gr1mmSZ5lxKtm+CpU6+OajFuk/HNk6JrRGp+P0D2/hS0sVLb4ui3xbaInbf
wxf/R1roJuEDL5SFltStrB8KmaGGKk6XQfKS5XSA5dGwRwrm/zYWxzCc9qctrkphfOglK0hJPrqG
GkfLneRHeVnJfeGJV2NpJdmpnJt2Z+AkbBIf2jVt2rijwt4pPyrPgOVGBzfI+CscZHzVXmN78/Ns
GZxh+tT/TumtYzWBcMLmNEaI+ZSo5XeKIgf47b0dGBIfXhyRr4qTmzWisEnamWBH7fBnTx9Di86j
3lGbXIYXWDX3OMb6dklRvPPOJhfk260G+ZVwC+i6K0YY/cNaTCM/Sna1TBJIwBYXiBOiBkeNhGLb
PXN/WQC1GlCY1E9tRxH8ZjzAZdIhJ8drCADJ98FEHcchBqBeDSQVJcAvxI64HbIgUOAKkh/T1w2U
ezJa5mzCNd4xD/n2KJ7kHybt+Z+cjmWFGgWI+yiiYIPpX13zUgF/ALh5cADAfD9ABdAX5S/xs8n1
hxIw6Z3UhQfjHG6U1pFfFmsaYaHuO4pRBuCg9D2T4baNTDxzAYJ6jmgrzuSKC8fUsvqSuLNDobg6
fi9Zcs7tV8vwjeVzIgR4PT8dcBElgVN3b27E7ulL9i6fZfEbEBkuv8+DljVXswStj+RDEbwaO4Jk
4ZZ8LuTZAtPtOK82RFZ7tJoZqOl0GxnYdaeAMRIfWGVuhrWN4zraz4p907SYUy0kcSc+wJAhzrbX
6QN7yoYY1mdG3KeTMLC70cGKwDaAmxRk/WwKaAfFuPbCZFTRw5UW/vz/lFt4LqBXrRaNFhow1FMa
lMZ95E3HhSlDFqyjTeLKwXN7pwPR+8hUa0SDl6c5J86IF2QwyreIBVlGuOMH7WiK7f5cYz1wu80P
4TY4vy5oegPecsCxDLhbEygK/3WO2TGZ3VtxC/3vgM/lJJhs5g8QYN7yXJybZqr2ddv5hEbeeG8S
iDSSDwiAVqg7Dhy/P13VnK91VfWvt4gdlhjaHKhfUqiEjskCCWOiuSrbM2EjTP15QFNYqwbzSPH2
JfDBAWZ72EFdNw7ctZ8rnLlmFNv4+rHv9b5NT/fdRvBZVwiYjW+SuePS44TdH8WP3yx+cMbCxGuA
ueRIP5aS/CjT6pkoh36wqk33WNhQ00JIaoUQRbT86xo9HcUMRS4Y8kwiMytYUo5G1bb/uESUuoDH
zAqiM0Voc0tTtkoXGmQ9+2iFkVMSnoeUx4lJ1shn/2/suqHcqN+ExSo/XZszEY4K56e/Hl2JMmDP
Tx6XLU2petYvQPh0Qz81Rb6aoPeJwOO3R58Q9oXQT2/+Ys7EWyUmcWllMPVOzAr/yAgPk1nSa1+Y
hmEoTdn5sGBywhq/LeH6zZRb5ZZEQbRQKTQGFdFkTjmPfPUJADXMrwRw5Tz9Dc4vktS+0sjpBqOt
Caqzggr0iegdNHNuLUDlTLExcfPxh649lnp5NM6jUlLXNiPYh7HbfNuohh9kMybFneH4OVdA3i8v
dA5if6OP3YqQaRti4jtPRR6P7miWxMUDT2M+s+gS+Z5x4GJk7vLB+QR1EfipZ6MwfWCE9Vg7YQZn
UR2XFd1nbERcRaUnEek0FZ/PHorNXwGJ51QoCztedf7pvnxl0bsimtnh816jvOjWOVz/0c0DXv/+
PkMJp7zP1rd6rxP0KW8EkEjMM0J7YuGhntRXgOFh+pz0kFhjEMnU7F9Sndc4v4GDuG1c+dj3ahyl
RMmH0csibd+iIq/kXDCE1kX26tZTObZKMG+UgsOtGpBjiXjZLb1EL//cF3BIGCfP2J8qia8n9AGA
VmTVvOLzLdyEm7AoXi1I8Wa2BA7W8kmnpdpoZhi6N0S4xcatRNyj8eQetfDdZzKzou1yvsAwkJq8
cygcLD6THouAT8I9dCbp8fGzc2Qw1cUPPSu6wpmF++PSZRdi+3cS6Y5xxs0V9Oq7PWkK2Lpc13VF
wZK2tfXfsTy0wuO/+052llxPOiSymA4P4mT1p3NQkgoHQHO9b1R8nXhhdjkt4hd44i+NsXhPu2y/
92l/5ZNzVvIHMx+RO3PgqJAFOzktX6LAEhPNDJyJir4RsHFkgb1tP/3xH0vSgw2xy4Pu4yUIz+77
J1p0Bu/HQRGZ+SJg+3T5HcvAHsWxzbXL2dQDm37jF1qppmTHPFSG5RD8B26Out137Gq8UWDXI7f4
+0TvtXV0PkfFjoIeI7AC6M5Ae1kkaaBtv08xItYSITUznNVJN9thcoSIvoBgDxx2GF1qExkoJBFD
jDwZ1XROq0+hwE+ogrIU7lBRppKwX7RFu01/bsl5GKW2YOR5gNWwXaRcinYbpoH0FDIA5tuxZl6s
FMjCc/tC83RbWLIkR33aOqL3Wuek2PNCg5IbxYh2Z26UJlHvS+P9+SwpT1OxDVEBlqhBedV7VbF7
Z/GH0UkueAicHtVimVPBdM6M8j4p0rAnVGlOvoFVaXA4hpn+ITwR6tmKQSrFnSQ3v/yLei7SOMh9
C/RFFMepwV3HpR+2PyOLrA35xTap+u6SJ29GtGDhZnoPd8+gBNHXLco4Wvc/gw62VaF0OgdUkVbd
syxy8KhFJnjiXxKpHusl71969U4ejd09N4HvzVRxUXpoi4TWrcTA/jUDhTZVjwrhFqcsW635UcBC
yHQdbaOjw6Wn38RIINH2/pYErYPz3SUL1bxVvXN6i9MXUVQcJJxDx1T+6ZHrlw9wf/pGBJEb9pMd
cjI0Yvji9wd1svo7OgdMU/Am/G8ZWaqO5g1aUwL71Sl6rmHYX5PwjBQNR+XyUKRGNu5kD8Ys0sqq
Zg0rhyMvZl24oPNX9Oa3L7NPizefGyX3652dB3qiVG2dOgx8AaVImB8AutWSFXUjSpntUYJIRqaI
gdIU8oG9c2tdlCIAXFwZX+avgnjVGUscJkZDLyuCScsUN3b2Xts9m41yNt5Um7ztPQ64iQzyXxq+
WffA2a9jkiK1uOHI2M2eaQyG3wnHsgh7LrHfKgtDTVWsBVWeIfO003bXkfZ82FoIQg+RAelfW3aF
hthMI2AIuSCSrb2Krso0ThGIiSxGhk5OVXJjB6wqSaj3XWi5iMk1wDy/CVlU7eZtsdNIp0OEo29w
oh+D5j0i4AGdFvz3nSP9QEUYysUq7jz9JgoMmR6gWTVARmheu/L9kgYx8G88MGKnP/Mv34dqVb07
/BlQdzfgEtePU4byEme9MDJy8XnO3eCc+8ihtdVEYDsocGjs/oyOef4csydpb7+xhz3EP7o20ZcH
hmlZUEpiJ1nuKX05vFTfFGCyEmpu7bsIaraZUAXO93iWBFZ2Hyn6Fju9DQ7xohxEuS4aHi+Vl0o1
xLAduQwiVjtmV8/BEhb2VHrUWVeY1lCiqz6eDYb/PQKYHjfFt32IQqpFbAGWKSqwabioeD9KH3se
EuLyEEW/6xKm6D933rp6Gw2Y3dUeuIu1mGOkJU8wyKcmz1whIg7tbEexHAOyHywbP2wZ6iQid81x
zK2+NPp8m8rWq9mndS/Y7xML5tZ0NlYT5lmtbZhiDZtu/aJsr75TniQQX1JtWSfMKccu5sRTgzzy
I2oLnnXgGLmUPtZTj360LYZ2dnD7uTV2o1yQU7ibHCGv6C9dw7TZA49vwentnlkpZOoawzJXcyMP
wybHOzf+Q68kvwcahocar0xuXLxrCkd4N22J6sqVaxw9+DYZuHCw4LGLj7KjKocchd99r87oeEQC
nCJxLqGsyJ6XUUmt777fo9/aH9PI71JGOZ1sWHauAdomJJAfm+qEjWfpf0FU1vZ3sZSHuuu/mXpz
iOGaYjbAuoe5zr1QauRI4oV0iv0jhkLl5PlM7RbhWl0ARyQhLyiDAzb2jtDvy2cOQXXnXLls3zRF
AR8bzl3w8W/HUay+dQc+q6/vQzbxU2oWgZ3G61FfjpvQgzd6c7pZh4+pQw0AyE2LMnZDw1B2UBmy
JOMa3UfvJGqjbQo1DP9Sr74TGB3s4WLavb89qmt+fCxTLDpEUK8QnNcY9wQni6y5Ei3w+LRc/qZk
6lwIcOQUw1umfeGuag72RrX2HLl4aABrOPNhFbt1eztFcRh20R6ZJQmIxA7DyWd1qZdIncu9g1mE
FeBPtrW22hiR9/KYikuEdfeRUcohRQaX6vZ3LYzrbHA2+5lh+R+CQqfvIme48vL+8t6HqK++seV6
ah30yX8X1Ow/j3kGKIb5VfabGdfALs2BiXTYIBX8c82EFBurgDQeKIbTgOJ5LY8kODmgs4LivVkS
3nXdAiMhBjlMR7eOxk5w+X3FERHmHyR0qEOkFBahGvgxKoyTtBey1R91PfOLrThQXmRLqBrxCZON
dcO+rA9Z6fjNEpVhM9EFwckqv+QG94pq33QWOjeNr2SZQEiBi5rQbrN8swGOvKPy30cScX0UHn7x
2GWiee/7XNEcw5SQM5NMaq9PQ8dqdGW+u2TWbULtaq5kKudleJ7mhGVMozJXoylksmZRA3HFUnw5
A6qgYw1cVMJvCd5zxplLHUigB9SritZF+pC24sasPpaSk0mpcJFH+C9C+O/aybpaR9vNpZ5leByD
xc4Qhzqx1tbdQ1bfD/OHaQmQtLZvxC025J9NmJczabJVqgQdp9V45qmFhjs6f3Xe2zAjGF7wIcLT
gvOUJz9dfwMY0aA/rYEILUDPCNZ0/9JyGom4gD/JghfcfUxTPgG/xHFHaGjytgjNOKafXvvpE2fg
E2wDBYPaQXj63FJ4I8jXaazrzpz2FdIzYTupFT8qe1VPATyPFZEaBVqq9jcve1c3kkKXlqynW0Lf
GwzsBGCm0OvQc2pqxfvBY+71iIxhMqxZzsiR1gY+tqcBmGytvGHJxX8JVgqGAsgD2tKruu5b2xeC
zW03z0N0W//PDC/ZAMvf4v27z2hANOBPlBEb7d/SwX7TeIuuoqPillMYqDP2dg03I5RoH//yDAwe
EC/Om7qIw7LaV3vb1+FOUb3fuvquwLmyf3maIAA0M4qUkK3LntvAakmGchgpWQ3tZX6GC+0mGnkd
Q9IDG3UuTNXqI+EhVB9+x6O/+fbg2Kiw7qylFu8NPtUTNslgEQUw8OINaEZ+632WXKNmFMG6OX+k
0pySEX4zyRhuUxpL2IOooEPg7v5mk/cWxLksiIKr75FVUhyAAPxB+MuMKUpcS1lrmGxdXt+hPFRH
I2wvPaC70VodjBpKHCHw38iysN59AEBv7GLgmyOiUn4VOrLzE4wADcVKV8Ka/ifPmYgBvYKREVWW
hcFjzy2KqjHCA1fYCNSoQL7dtLuQvkJWzu2S1fRffvWoOiUEKgurIpXCgRNRRKkWX4DCOw1SKBBn
ZSXUZ1+dq/bQckNpcW42Qr3+WsXUxZUXseL5Xqv2r230W89IUbcb+ZpwPvpK4R3x6Eyl0fKkIGKu
C7S9OXehGmzc/BGe8h7CeeXk0JzJYIXAZAJ3tqNoMwsmjXEIEe0ax50eW9yhSLI/yObtnjuK2XSf
3hBpxkuo/EebKGUOzh6y+HvWxGvuisNdAHNMhXNE9aLOhIFLWzm+GQlnEN+2XLxCn+i0fq/WIEAd
PfgYEsMnBws41uo7vD4IJZ3D+qcwQR7IozkyuHgBHM+A+d1kbF4xp5pPrqtrw1pzBLnLdjuUHikd
MYDc+yChhxJaePFPhem0Gd0S3/k7rVxg90QA1lrBhbG5EOjnxkf8UDehiGi0vBQLMeWhbO5Htrhj
Cire9cDBcGHsjnyadjS9HHUeBbDiUWBB4rgJbtlNxgnohf9vbN5Hp6/ZFmvmbQn2wE7xnblelnUT
89yKSmiMBDGQbEKovP2gJsHtC0qU/yHo0LG3sIMeSHmAamH3fCwTVUkzQIJV6HBIgJGufsWn/fa6
48vfpDuDdfFQlo5O+uZFMiPlbsnS2aksL7z6AMfob+6mGpBK+QgPhfJ6UQgjATO58IizWPw36Zcs
1XZ4+yGYeezm3u5wQVTdqC2+uQ47okb3VaN/9yoLthUyX5S9Kd+u7tXaSJ9/G6hfjZ+sSTSuNXr7
Yo0XTKrmybvWI3hvvZj8NLjEzf9NQbrSymfDGusC64d4PgfYcTG573GhnHLT5+qhJ4qtfcwJBfzW
tUKxJaBKn62RakwG1Hfmi02qirvi1hMNEfEPqA/vsi2aVT6MQh9bcAgQmaUJFirzi+/naYS7H5Xq
n/OtxtygDoScC1eJ1g6OKmmgSexe0fodk6t0AvCJiTYyHMKcURsb7vkzv/MeCUsugWNxfbf+4cwW
ANdvhrcGrFZXdvYWzQSMWZLZSL1r38JPmWN2jjtU3HQTl1XFmp9vPi45qNiVwbOd0M1Osa9tpGzD
Qt5zfDP+4hGbcoRcANghygWbFoI5A8RNgeVXApmlYP/CiVSiiZXWbB524VV/hDYXntx01R3rmkHC
vLUnrHsU0IGHm+LFX7xCfRSCUP8HCl9QhUhMGiKliZYktYIxJiZFENPkT8CBIs9Kz0rE+w+khfu8
Drt3BVhb4USC1PlaDRi+cwd2GYuZ+OD2K8+36Lgk9ZR3Ld0i9ZGr07U4aZCiVrSDpbY6rkiNK+7t
0P1WWV4dkBYYdN81OVwQz7ONThL94Pwxkk9BC0wDgwWvUdzaGwWc57YawVSO/fZqiKPJi4YR0XKz
xhebJ7Byx1Zjdsd6VLYe/9/NORgiKO6cAOApKYXa60Im9Rm4wxi1Fe6PuGiJbAGkQcCVY4nQcerQ
cGOlrtcdYpOdF5jeWRAS2JhLTNrJabHPO+JMgpDMWVrFKCHbjHk4r8r0jdGljD6BJURrgKDauVJK
y3I7C6mQT5R34wQf4Y07lQi1c2OjAmZTITOjRd13koOI5DnkmaDg4lF4830BdqaPso9jR3GV+7Ds
1JHDp+yGweI5kVVIluIkkLD1IL8qyp5w2dy5tpbKzDCcGDhD7F0+mCM7wzVblCf3XVDjjpz2Zie4
cr4SzHu5lijLyIGuMf9nTzzachoV8DL70rMGS4wx3Al6nFh8JxPIVVpsuQtTntw7s+w5bhxK5dxy
EZo3a5J4tN+LWQhwSWawm6m5hrycOz1NFlgRkpPjVPOcNSsrofsHy6ngcamH9BRzadQLBaMFINPN
TpXAYk0HnhE8clnEiqSqp4LC1MtxOIUYY1wCU66noHf6cQy/T47txkYa5cSKb9H2KaVjajWknLfw
52zriHTS8jO7SKvj7eyMv5Wlgw9y3MsR5FJLwMG7JsLmEU84R4olKnUiuCGmfddcaI1AePFl9HN8
HjUgf9gkkCkfIpbTg5IW6W4uCyoiUwWZeFy/Q4oxBSIxUgplkRmRsw36I16SjNUQjc9/mUkwp/IN
+KjxzKDUl0Q8h/zYFZJkwM1jCC2fWO8GXh2BGqPK+yJ1ULsGU+eiSxuR6nx9z5UfiFnIBFWdWizB
XObvVB4xmm2sRtiLSeHEEbPxl9ClU//huJ5kzh/58yVidXSrf9gqwv70+7o+2M2usyRD2eldaH7m
quTvotd4ZS8N5geNzc11/9nWkNk1ZeGESNtZytmaGVaus8q9jcjZpgyTfL75ce0RytexEC2eEbM4
aziztrytXVtP3Zek7dvmwF5pHEFSZBNl/z3KqwdNCmHm+dCqWRRR3yfKax+WMFiJhXIGr8uqTVra
/P61Rqn6pKHo6yK+VZ8OKVhgADWaHafU7JZTqyothRQr3g1cXHUEd0GYpS56B4hLtXkXe43wGVbB
HLcKwmJ8TtItnTCl8ruB3+c7bPqMEAS7KZhUWFXoKmbjTSdBno0bsPASOzEXW+hX/6W9XTfQXgmA
S7tvil+IivOCcI8BcK7352XbPRkmz1D2Yt4aDULVWPafOl4CFecBvXGW4wkYgvJJqmA9llnKCCF5
SkFtzBegOnM4fhho3KWO9gOoFUrYU0L8ZX1rCpuzkTt+ou/gTwffN04ExDJcqYZh/kQYxNrjC9Si
GXkWv2R0n3JmmRcufzlGBUtw+2JuZzzpQ99vMm95/b7tcgNkZFzCi7jcCo6TipbjQC/z/NUC5//K
2z/j5WHo/1BEkiAUVoHIKC8YkfY8nTjxsfNgpLAQsQGv9XePl2zJbO3xgbu64bHJ9OhkGtD65RCf
yscxrMljVUjxqGJjSz8kVhJdlNwrlnRncrxfeW5DDLflxpEC9AtJCg998lI/J8ca8lQCwAKfgCAe
ehwuCyIPLsV3+RIXS1SWYlDVSHD9QabrMVYONSMb4vflhH75mPCpxI5fP/amlkzCf15aPjbPhCCg
MZgOhgN/InWtCfxa03ja8JP4GADf/VG7JMOd/W2sF1cblOEhUOv0He5y+OVcbFswOPV7JrJ8e4PU
2KdCMbzmKHxU62gMqI/KiLHiYyMeYcQoDDj0FwKBHfh529YDvQTbCkmhEWODT69EarYt3hft7leb
z2yMk3SlLmN7ZhLcAFbWeXZ5s4PAjibqjWNsOQPrbal6ON1LKOvMgb0hod0nqzQ6oAsZ9DkHg92X
YkgPLTB09rzfeLFRJICa2viCRHxrCtUMcrNJB8tN7zApPUpsDsRv+sPxmG2r8VVfFO0LgRRkMBKM
IXsaR55jWtWnq+S3ouW57JpungmcxwG4B+w5HCIw+hdX48ivAl3GgBRNjqUt8KfDwFeYiqjAeEEo
mEXZ7H/zRgwszVGLPxs+5nVGJ3ezuzvir7ZqV58kaD20tC1SnZCDBdJNszw/AIlDp8uXo58+aPg/
XOGv1fXrOShcnSZqU1x7IthUxFUtN9A60Jxam83bT9wv/lLTd+KNtTuG0MngNeL0H60N2iAbh+Ua
sHzPM68bUOnJzNt0+OVbS+OYFQtCRPS1bM/PJvhwZhM4vq6SmnHGRqBrgsGMJ9qBp6qaIAohU4hg
9skW8rQq3cqDHa5AgSbPLV4KlvKQ4Rw71geysPQUcEWb3EadpzX7LEXnGF30xLVHDGF+q5zIlRlv
awY7a6SmjF7SLAXIyJOVvBXzpXQNzsdJevOmhiXJZka2ibtm8bJzdKQoaHRWMSGOPbHqAZojEiSz
sZWmVTXWfPWdHWf3ddXOCxWiXJUE4pCHRvQeguqDNjjuRy4SXrEt743K9BCHjI4fKJeZh5hxQMjF
r21eynlRqNSUMWljfJgSooISBkuHAijRLAaC4gqhUWNkXnU+5RLAKAbJxZDaU9krKtR5rml5Q+fK
EWp0L9lyFmgMfdgkGzU4NTHP7BVAv4A/jO+9Ji8bTgk6xXvNn1G6GQsMXyPD/mGyTXL/hlEQWjUT
qfqy1MuWdVDdiuQxvFIy6UzPhWo+2e3n0tTdkavjBr2P6mofnBKNjzImp+T3MJWgx3VV/LL/P7O6
Q4x9vnMAnoVNeUVFeZHEQWaRo1IB0ZRxXuB5FjOrYbLubBRX6Gr8xvpHLNSUH3IBk31pOj3hVhW3
yMfVm4LxZLlgg1DDMDMmOh+iCSuDdSD3fnTuvMH29rQzFltfgaibih9wvTke36I90tw6EBFPh5sA
wkuNXGPH5UZqIaXLheixkoEZL7iAyZJxzWf6p9mCg7siH/kIF/uwsgg59/zQrKlCiB8Ruzvrt0e6
Nk4nHBVNm53DaVB+xtBp9G481hCrVJIvs4b5Cw0vXJnlK9LsQH+bSibj56csQCPjTEzVWengr+q9
yGAR3RTpZmWElKhgjr8mpAc1fCLtiPYHQaDWKdDM6fEW7ywkGiXvDUs5UPj514UsW+1YhAxgYLqf
DPzMUfgwSGS0NQH4t21f+5jQc0B9FpKh6mscXMQmL5WElEM97r3kQLl7sDIEGNxLtkG1/qqOtW8L
LVceiQac1C//+oJGoR2PkN1qICK9iq0O/UIQEUTiGNczZFaULM7eRPIwT53znGiZPXfbmDYpMvx2
iu363iuVccsx8Ss1kIW1yFl/0BammpICSq0XvD7VDlLkFfmGWCQ7gKvi+r9egRoYa4jOlNxDZacj
JBPC5egHk04gxHGzax/YekHtkVJlpBIc7ynpJwlhECcmx7RwwTQxBH8tuFTWtGGk+WpKhD+AFGnm
pkDTosx3Lz91n4lqVXxtwMYKn6cWkMfisO8fglEtbRrpxH5ch1V41z3EacvLxet9osxpaxMT7Dqr
nKdRql9MIzfjr7saVveGLIrieGLhF/Mu5DzE0vkQI5eadlpMjbxK4Y8BUOn6sTaIBNTDAczCevpz
SW4zWZ59T0QF90aBYYZvG8DZc3bWBqDwGyBcTPnU8JHJuKnNg8HtAu00exk8EFfow1bQKD50Fzj4
lF6mqWzf+CGKJK1yWn8IhH1MzJ4DCjFplqKwYXvWqttn/3Dw3vs2baAhSjz+VhoU2DhUqKHciEmV
r6JiLUPlVL/uqGGUHI9RsjQ4w9eOSsG5BzeebXRPHWHywOivrGWXEx+KxneStzexylpxS7bZc7En
rF+NHE0WVS1YrquKuXixiTqSHzJYZ+kbVu1mPVDvQbXSms/0vS9R045IBmK8Iylp9DmeEFs5C/0l
uCpRs7oicPFry0GVSG7RUGHmAOJ1fDdQqCohi4jhlBzCMhB6xkf0m5i0iemaf6AR0eV6jhP1I9QU
MStpiuexDQNgs8jWXWMhh7e1tuGaLTinq85EipsSe+YNu7QBtoME3UnQS1KMDbxDlbOarNaABVIq
XqR7h8rhJIoRPRiKhXB+0d+orQilgy7j2e0Wul82CdnGWmav8ysWA6hvUpFzYhHYYdfyg5sriZ7+
EKZsyoTO3uFCObnCF6npQBSBtBPtco/4DIqbpCWrD/C04vI5Xbd/b2KOlhugEFqAl3BusTkfvOod
jBf8iqeoXtfndK6h0mJO1cP+ZI/qlgTqo7zrF4p2e+UtOan8HCqBe8RsMGCrDEcQHGPj2iXwGsoG
/RCaJMtXzIP8o/qdEJHC+A19qrVO1MJS+lwMDXve6rhVm51mAEiuyTRP+PS4y2J5JILLmQADFv7t
Hmf1jibvfR2hW6r5xVk84JB11Egq8pqEwKcsBIRn9YF4D/t+AjNnIpY8tlXskIKdxbOp633TmsT6
6/DY1buY126k71z4FoJVcKHnuMRkeRuHW24RpAhF+EG/bn99V4/v2TrRChTPEVe7yIrxKWE/ifUe
84KAuoBIv2t2FcekWMSRoBIXEJbW1YyRlI7P7Xer80blZisSMc6jH/S8p6/+k+97dptz7BN3nlrL
z70t0vkiViIb0d35Ua84rk66OPCcKUt/EkZmES8F/M1z2nN9ZkdDZ00y8IojV3S8I4M+mTuRKcRM
MwWPY/rNYDGAeyHDxEayVEx6kti9ZqpOrVkMKiOdpXlyn5uAawfJlrbdzT14eqIidKaLRllAWyX5
S2ZzZuI5wb9EjMoxctu4mmIlnERqb+LCudtVvlJ8idj1nf/2Xtu9ec6LlbYTsWbUO7zo9syTND11
e1gCF14OFvivDhOYPR/pgwO13y57JF7oMFWLMn+EcZyobO1ZCzmh479sGvuR8t5vOc3j5579t9/p
8x8655TsRjSQR+qRe4D1+H8jT0ChyIt5NXxcomKs16VMvhtDE/yk228lP7pVK0+oX9nr/PBTcCqo
5r08L2AIhhC/Xl7ChZ9YGVGnH6SC91rDjq7e/84dOi7+SmhUuMw5FVQu4MbpnhGfohcb3NRGlcM0
kgUbIncpLQOqSze9FXdSDQP5maC5iZg1aPsDi+pXSbNkJgrUIEvt5M0g2cXG0CiuD8x59a6ZlS6T
27cUgippx1pDSS3M+Zn4QAIFXuowz8JUeO33aRL9G1nzFbttjZf+hOLuevUdzf/dCmbm0UaR+Gfz
+CC7WHRPkccqKbSSfkmaq8JDlJJgzajeGEg3QYvX9cOLIDbosSK7XeAQSlcG9hvYQESSHXwJIhv0
cNjk5ecivYD0MFTsSN3/1Zln1tAJ+RCrnnwcxPPrfCOaT9VGpoObSxV6bncbBP9ZzubaF7YDGK0o
G4DcW1H94XGWftpnOwTRV4txZbwoBIoK/5SyLZSjvgXgO5YhiUjvAIqYuX3oYMtfhOvsCEcKpsSH
9oh0vH4JnnhXPG+FAmUeQOfXZC1tGuf8R7nhwgiNILDwt4RxH/SVlIV/upM/SYW1RHL6XC1gj6J1
INHDgeEWcSrKwIlaCqiUAcOe/fg3lhjktofePzHgIbzR9X57zj7MDElyraAcA8HDjIZmB2LjqDY9
pjkJvVxZmHne3912RQ0JuEFQi3OXqgcSsWFq78p7FNYpcaJEyUn0ye0xCwZAb2eIOcpPz3yYva6z
foio/umLqpN/Y0RahZ1U2ZoAInhXvIC25qbqzZXdNPr7kVp4+65c2PKq0ufOC8nmLEHFLfJ/o+At
PAxrEJPVGohK66FfV3gYazFWJLVPIokepuG+V9OT2UzXTGcBWa3FJS5/yidxQxZpcNHRmkOpsVQp
+7LzmQnXJ+5b6kZrdzcVwWGLGTku9beC+/j/uxMuMBDPivqSFkXP4NIbWrA/UaeVlqoa939lZcA8
PJnZlVMULF70QPbyqJBBTDd+C5dxiwX+dmr4lQ0mHiLZ9ZIjZZ7rhEhlPK0UQ0F08rKDT0o1NlQ9
EELpWNWbI/2Oy2Lk35ubsCYjwbAjLdVy7WrtyPDRVGX8gqE3waYx/GTuwfl/5B57wGdZMDPvNyPj
8nHi0+ynEzx9JwBPTfk0Ug07VBn3FAFu5DYcTCcqrveCqJmD8jwuj11o5KXRhH8IwBywREPMmmeh
XfDnv0sBhHlCZbeKwqr+GdnzpDp1ja9/UdcsI4fQ7Ra0mbXRlTGJEZJ/iYBtCs9H7OkmPgOw8ruk
jScdgrQlA/q1Bi8uGhWwWxdFiraCVYGvblT1pUZ7d4M5oT7plA5Bs81gBbALnEbNWXbpMKqAfpiG
dook69oqnLUxsy7AHlEpBxQUYjgEB+rNOlIwo+yc/12CNzSIzzcgfbwRYFVK+8KsoXr5KSxVdYwN
CcuStUDvybfxa74/f9ID1HYqV3yfbw49HKHUi+2nnO4JicJmfoLQMDnvMx7uOz0zMz3LQ1daPnvU
sEySjLcx2eSElrxBaDNMchKPNlOaooiuu28MGjFlX4TainDifw2zothnI2iZQC1VFe1g05FEOeCu
Ygv35/Frid3mSC79vfd7Y+Co6MDpE8BXl8dPEbkC9NMRLpLGucuZjepo+gW0RyqMncBGryr8eI+2
Ut4vbyj7Nmd5x7Ugx3SfuxEDnbpDqwXkuG8Th1aDVK5y+ZSFatocD4PI+eBHj14OrFpxSqj0Lx1t
4bU7PKfMOOzpS7LqnT9adUsswcBVQq7VLWHnjU2gD+nHyTZXQv+SQz52gxInFSxyWOG6J/NV50XP
5VJjMtEztsGBEAcmRl2fG9mde2iz/ao5ZMZROvaFLr3R4sFR2HdCBZdxNwQxwksPhPt5euyQTBVN
q5vlzJ207XIQY18BRcIUzU7qziBtNef01St/u4Y3pNKngezm2Y7JvD+8NXikVNtHPF/5QSAzDlVm
6cSTF/Qc/TvNvRWid+daPqIRSozvuNg8YEJdCMenxy2IXnDJJ3EgSZxUbLlj/5k1f5k+QcpV8vBt
w9gatDKwIyPE/7XXy6dl4Oeex8IiOTdMWez7pXIBGzPFuR/9BfCqD7Xy/Rl7JF4Fd2W7oKbAgxV2
0/u7vYLN2sJVkBWcEFHbsK1A5STxjKYjhI0dfrvpiC9w7+jjlOJ2LU2HacyeKjwFmODR0bMyDYfk
TABAbo1QNzQrgXOhQlcoHQmQSBgEm9nKHjjJZpqfta1KTyQi1lcUwL6nQ5TAls6o2Ajso+A8LjAh
0Jth806OXwP2GOkqP5s/U/1NRTgDgvfOb1aSx9W4+DgOg4xr+mQ9e+vu2e3QrZV2F+qPrtKl8VWc
QZAUXq0W34Ex+2EX55muWOIw3RtHVg7/Ueo8QUOkcI82Txa95aXNdYzpvaFQW8doimVAmRSgp9ME
22xnSp2rV2VpUVITBeMwrG4Hy0xXOzyarqGCMIZR4WJMSJH/3JBBULW2XRw4mF+f6xSwG6TtwnBM
bIY0vgH+WaR90PuEiWjkl50+Si7WUdlKZu8iMdyAV04QUN4GfkFIwk8qQP9XOBEsXntWP6zojXdk
H6ykFmL00guvDdxOKs/ZnaGIVourrle7hb9aO14wU/ik0k8PMPD9cRPiCaCjCZw5TUbI1V3R2lA5
h4lJw25DFc4tsvEwOrYNQo/SVt6TGfsqEpqDp0THZ7eCPRmhFjHQ7kxMvXtaDjATWG2D/3kl+xxt
t1xnq4IAeYgNQa1c2paqazrAjiy1d9se7Pf3N50lYDgKc0FdS1FH2MasVgPx21mg/+MNRucRr1VD
9hOiiT+Nk68beOaAFFRnFQSvHY4SdMttqYPNJKKhjE5vx5gBYC4A+RlizxHAci8UU1S7Mgh38fUn
Uce+TI1Byj9fEdKhXJPLcyxI53MFBfMxD7bMg/bjMeSvmzFsLpAmg194t2Ri8gm0A23OkqWVYgDG
QEIAPPBHEHTtBCRkGP8z/k3lMWdP06vwJ8okXXtzePK05yeynjcQB5Axx99iDquIwa9gwp3lbzeh
9a9aDUek0j1dgugSPZznxf9RmgbBV03xHt+H4YI8VuQP6WU6coQVYstPlUdppyP1LX34VkLHJOip
s9eWPBrj5/eDed9LwYuT0IKADoJI5nrqlu3pYnE3xEh7W/GelpwV13W9IDqdxmd3K525ul0F7nx3
AfGWKKS2gFDJijvhpm6Xq+l++WyFo9HVWwCFecGrEB3MeXpUPy7LBdQvHXj5vtvUTaH//Zbk/hS/
mJq7ozOz0d9xRKUi8DvAAQItQQaafhlNy6fEr5OXYa4JC178Safrpe0sv79b+R2jKYtjRIvOC45C
M+3+yJ0poaEAsYzh+9fcnvCN3J4EnZ0TcBL9dAtYIIUgjxpF8TrdQ+690y59IkBTElKoPU0zOus8
dV/AgEjb6fYKYeIdm+uGhJ2My7hDHz86HaHF6Sqjc+QdZUrQtDQmeuDN+azGgycL0fzQ8Ju7nToH
2H8G08JDgelUcdcTu0c06fiB89z1bnJKtpHz2+MeI+ub4NEoRW+kQDqQ5JiCE5nwsDeS+s0QVpSK
JAEEkvzxt1azYAgZE3yLm1Cdk99bf1CYZqGPaU3847/2ewaH3mm8OjTtU6RPOqpIgz35/7c9lviz
GIeKiv9R6R0O/G9UASMn8o5+n4wbVtCgY50SXedpbyVbSPC6Y+KH1JazNDuqusmyWI5sD0xyULxI
lJCqnG+o4CW7Q34KPTbH/o+VpWtssPd/07ME2oyytW872CwaNUxjpwYZ6TYz/H/A0Ro6M1M2375j
xBJiSJQCqBRvB6vRpCtiYQ0o1xD0ZQUwcD9jpF/RuG732weG8fRAiBi7xfj37jTuIektA/5G9J2/
itpURiJZ57Un8PePgfNdFTboX+Aq4qPIuOBrAbXZHEbJNqK6DkxXS4rbkMh+K3NX8YST7KR/O1PG
zVijtE8uQObYixaMzW4DwtzehCvmdTGybgPjwBCDLNnPYO4xtivEyg4w5aqX8MqPZ7fLIgrBqhPV
Bv+b6rf00EFJ2CRG0L+dK0s6qJMXQEe25kvazaceWo8JP9ujjMLeczkEKha/3xTVCdQUhkDAyM3/
R1ipGOgn9buAhcdfvNqawOMu/H/nNbsiS0//6Hexd6QVj8sXkJGddQgm4m0/XBGqb7C6USWZg7GJ
912o1mfhU6nwOcbyjtDcLqtzdejKJdfsS/Nv2oMf+WIoSUaoCn9u5Pl+3GGNgZLMz2kYaVVIdZON
NMuYhuYITxuJj1L9BCekHlxx0lVScBMn38pN0tNDwhDpvqmqX5G4zwtCnxmUO9i1VJbVM+cdN4hg
AF7G/GkoD5HpSkCnq7/6DeowfOAh1k6wWCfL3qSPxRaBCnIueO04akQIVwaxjZ6E9pCDM9s8wnLr
haQ1ZXBfgLqq8mVZ8E5OtAqWhG/O3mkQx68IAV+9GiUy7bpI+LVN8nbt4CnIDIwgSaV/rRavZhqo
2QQebdy0ta0YB+SRfbpZstgAx91QdbYQ/5E2/HpKeXYeAjm8pwYDrzmMU4GrlbmkCrOz5Hs/K6cX
fB4Q+gHCHUTBKaFJ3tNirKTk/wmo1F4cHrB4Tn5DYYrHwrQQnvVG16be78cKABq/upZCiZxfParr
LAQs4v54Ek5ExKwiRRdaNDd71u6jRKMGXqWiNnAgYvIvaLSXv78s80VgwR69Uz/RjofE2Ps9TW69
TiR/jaXkEXC0i5o9GL4w0UZA2l3G0oR/H4KTdwNrkvm/DZgeuXLBJxdp4XGbpniEWYUGHghMknr2
DlL5CTyYteLFlRcckUj6ujDKAKNTu6EB6NE4YvdRAEz6sflk6itPmEBo207/gfoeju+CliR0IDfP
zm3L9AFZzF4fYno2aTkupe0JDnjR7/sJctBo7jaYOd1h18cmgVCyoo4REM0g7XJ/g5pu2CWVCLgh
3EHgOGTHxqrBHROwv+QxQHctiJWfSRww0N2PhydRzloMn6hHlA2Ob+rDAGVdtG1YLZKBaiwW6epf
VUfXRwcXrEsmA6dPmrvSTkjNiQAFWleLNQvenKwpzPrFEjPROiDWZ6e6xgmWpshKKNHRT5mnmxY2
iJwE0n3Mw9Hi48SPWXE9cgwbdrjb+Mvuexco4rqAiDBPSP8LsXqeDVJOsl5Lc4HsmT175WYcPSas
FYfkypqZwW82tbrAx+9Nsx9uWrrGN6xRf0RDD3Rl01kz3xX2FHEMdkGwR9bRJkBR6sJc54XfbIoa
K8w+pJoEB48xA1tlqiFl637dscHCNDZZD2mASyY6OjZJuwLGTqOHsNkIVTfJ1JuJjwHdpTJDDFRD
OecPzpAHMWVItGiADiX1ty1gkDIQMfFl8zjRvhyxcvTYehQtCjPgofpxsPKDR348UBPzKouT09aF
mOTy2/xN6lvOr50NmtffOIUi5jJwvSJBX0X60h+2ly4G0dGDCKXlTkPb3Qknqgqr5IlwApFcXLzl
eLRpvhAuqWWYo9j/v6aAKIjQhf/xoO5WGXx7yBSzDR6X6Y6kgfEGgPnVOfX2O23RXyRdPOqSu4ER
pVfiuACNf9m77hJntrOR9vq+6YzULGXvIIsRVXUUwOKtT0SS1RDguZ6D/n2f/sWL9W8bH9NZWqSE
ZWb3jEOwvxwj/AtTkgfVwcS2omDFhN20rw3QsEbvoYBIaovIOBJIIAO4CTG4SiDHv+02eF3PdUEq
I/cbY3ml/j6kKUb1vwEQQUCagwfttw9y0fFRdYPkH4wO4DyfEwtrWL+5z/hhCpE+zjIpUgCaNuxf
ol5El4gCOGTn1ursDh8YH+KHIPAf+Y8dI4W2UhgHAtp3qFax9vTaK2v4UFVhPJiwqevXl5lv5IFr
+B4TLzzhiX8Cqw+yuwyTjVtHsRPyhVI8wlGrOMhhCs/1otpgt4PPyQ0AYQeDa8ufz7HE8f3sKFUg
uIB8ymWYb9CTuiVM4gU+ltUeGcHs3R1pNX1IEhl70/tEt5izlW1s1bpvEosnXR7b4FIAT8QQFvfF
w5c0yN/PT3fG+vbbAwWKqmXhSZS227BhhoyvbtxAYKuQEVLceG0tJGQKxSrQ1PpVAcOr3NRYTg55
H0YWiZMtOQhK98Re+u0Skp4bPmBO4FH4UfSduaGSsW+G3Zzd+eDCRkAQIvP0ja9k7YFnStQM5PB6
h7Nn/cpbYzNqOfnlaoLfu2ZUm8aF6O/dbygYHdx6OeMoNHCHkGUMmo5pDmmZQCnNQKZYHwDslQMS
46bb3GYnNaZX/7geDoh+mS+3kJWXkz+ga8XdVTvThdjL2uy4KzZqdOV7XmcErWeT62kSmmd6cO9L
U6bAiH+jVRQsZpPO4kMp5mMNfLby1Csk+EHP0J6V6GD/0xQ2KrjmBVuJBFP/RYM4o1tflBvvgzkh
7lW8IGAETvbU5iaoGwVycfGIVlo8RY76ZHlhLFH6WyrCO6kHYVBoBx9rlWYMuaWqkf/7ljQZfJ5z
z/FnxzZxZjB/LEPRH3GeRB49+pI7ackSCvY7G6OuYFoe198rQob8uvy+70LpMTirugcsKIjbkJHP
DLZDBgMOQPq5Eyr5DQ6MwD6hJJfJ8upUWrmhCMbZGSL2u0SKgGq0h9PFh6Rze1hSjqmwsr5Ga9Oz
N9uh/zcmhLGP06PwA4JNW6ykMbPBc6TwD+5SpxTSXt797Ed3xp8lHKJmYghGx6lfJwB5CeKVqZ3E
CVKi5Re6k+vmFM7ZyOLpSZPxVF3mCOFZ0+twEy2GBwqtdnrczOma91Oa/fOjVWfa++/pFEwC8HBP
K93NHGKeotxjAD4Hy+McrdJubQilYVpIQqm8xfXQqVX9HzND+8RGKhE++b7YCqEWlqkLM+Cx1aq5
rprUeK8yCiaDMb+Nc25BB+VlZ4GeUizSOdpEItnlhK0mx4G0xRCf0scueBA48Be7MvSKoanCdmUJ
vY7gPv6vfR8tgu0Ku1PoAeyD/xH4MxCwRs62GGwKLjVMIKSS0GEwc9ebPDBa0YcJYZUHwr0mKFfb
6moh7de9kkxK+YRtY3Aa3rK/++T2B4JCCQX2W71I5j+8tQcNmYVUBxaEqy0KmMDczdUXrtZs4XF1
fVj5STwABAD9RW28o69NgUZ3kMsp0Whi2PZHOGFtJFwYpDqoT/qTFgY7hMnBobh8+lYXuJkt4CDo
pmyVFzsBGBzmnTsFhUCFfBQdglcUskYA5McpG9gA8QmBebcGL0c0JyoqJ5sa8F6eQQvoqhOEGmeP
+nTgBuq9/HbWsGfjupkNcxe0NePBrH+MKmbeMlC8PCoSB1VFkyKmULe3uCwML0d25T1HGUv+xlmP
zEZDq/I47fNmYi0MqNOArLNmd2DAS2UfWS8ZSMsM7zTKPgWEf/WuawDhNtnESRHE0/AK8JLLlviD
WV6H6g+7RJIhnnOgomWMMj90TKERlg4PFYoz7QiMQBqvHwQgVbS9KcEEbOX4VgJkwNJUvuVzc9GQ
UHh75c86w3SPqv98BLED2EF2fIkruNM03dAHidjPZap/uvh/n/5YbTrdYjDO5mW+EXP7j/dV+vDF
d7WpesW5oX+nucNUGOS6sEeah0nXDuGx92eFq2i5YyORoOW794e3hZDs5AKj+Ya0awWwf0vknl+q
8qofPNzqYJ/6sVAljG4W8/miEXP+DJT+g3MnCPOBryAPma3ZeDrJXlGaRzLHSwabpdekPeGM2H9d
yawhXvVjU6sZqZa8+lk4wXujv5vIEnweqt14DY+JjBijTH8PHk93kM01rI9o7O8HjpgJ4CoE4KA1
65SmlHvenw/QBKAjn4/vMC3P8FySFHPEa5KOBTvMZ9i1q2OBLU+HY+JPkQMeRTpx9NNFkOJAOrij
II/9+TyeHX62Ug9F0N+WHUhlYCqe5bfnp/2k6xKPztUsdJqejrCVuf646+Y3P0IiGYx4odUI01nR
wtAZnRQvkYCNAm/7PF1fjrXfuCs+CIOUZQhbHE/HUWdH0Ubi4LnV673/6eiU1nUDveB5e8T3rZHC
zAkM1j0R8do41RdqaADj/97lMCjRxJx2i+ILqWp44/0ALRTWiXxUxZgNG+rI41i5ZAyQCAYmhgFu
CVk+/VuBUmzilKvozU/G3PXdNuBcNZ0IGCxPgXZB3s+qzPglnXIsxAHWTTGLLsFyVpmKldXAltkU
w7EK/blX8iM7GzDwbvTGwm1oCaJJVE89ozTfzWnbE5XOISp6Nh6QAtSE/fHtE3r5J3tvFVj5wkra
0h8Lb1QBpCgEXJm/jgrFXQREJFpieS9lS/sJenYPhbK8NFz4io1kd6uiVeO5S/Q3E2uvsO35870d
pOzyVDnqlDVucIUa2NnkCbkuCiJzebKNJ0qeH0Ebupp8zkKG+BdmlpW3IZwMDxgXOWWPkBqD3XOT
FOQ38uXYTgLgBLvK4xwnN3ABOj8S+am2W0diTwkmzP9R9BI4Li7z61ZArESwyDCXwpoEVxejE4Qg
kUVSNN5sIMuTC3Z4UwxcylAhDy8S2buuebVhpN+XhXetvayimNGOh85BPN2DYLeWQM4PWDVYxIam
OjMOdKlNID9T2rp7Juk4AZ69991N2UmTK0zDIfI/vVPHR0HDMte6ddvHJzIkY/VcAyzRQ5MpzsqW
ipMiXXuEVNwCjszAIJSfOHee8tzYff9ksyUgnP0SFXOQ4c/plXbAOc4pPYyCjML3l2RkCpSBPCsX
RUHdJlgOy4+mMg448S0aYKQwFc94ungbmdDgIvIg5dnq5hXguI3yI11g93f9Dq9OfxMwaaLKBDNJ
7HCmRlnCrkaXIdX8XwsfZM7TbRhsoHpygKIPDlG3A48daCXmWnWFANfN9OUU3Osq0TaZajmthN6u
O9NtGZxs3ocZCzc11vVZrV0HV621j87Sa2oCgZP5bqkrCIX2YJCIe1sTwF3pDBI3HzXrNBPeCzXJ
WI7BHHSlxF3drVX/Oojl0YE3XzwwUweLBlRDRTebHnaK4FlFNy3+162y85zgUrMvb9F6iR+IlzPS
jE4DP3754V69Da3beuF9UkT6+n2StgMQ91UukC++yYsPulpp1x50K4omVa1u2IfJlzaUNGt8GmTm
hSNvhrzpBzmVFrLK8/oeVQ1gFPdwQqwJCc2hDWTxfQpdH6s7q/K9GU+ZxMPOrzXTjeKCCkwPL3VH
seQXOCek45ViSI8/pch/Mpay9/LUx1c0u2ish5S+70GAP8WZU3KWCdn4808uAclCUPXtutTiTv/x
E2V274wVbCJl5m2wn9jWs7SP6DZOWs+1slgEYPZ9RgmTOinM5Z4aRjZt/gjA71cCPrdBhurCGSXF
JKPO7qUjHrvHNA2/ThNv+vynbfasJt+5J1cGHvJAtaoY/lxHL/UCns/XLW+ui4LUX+WqWuB+FwK3
jpS/qZAlKCelUhxZZflJSbZmz9X2kNYc0542+TmFQjS19iPbn4R+d3DFKFoWndczVlXlWF+07NCW
9EDpD7JfGJ2xV8bz4Jllnht17jDCftpEDhHsYT2hkg+5+LGzBsZKWFKY7yO6wnFVGUh5zgvxofX0
wBH+X+azp6boAMtP/0pAeNZOLNOOujZTB1euGt0IooFHcnc9/IpjuXiuXYuz140+9MEUad5cHLGa
PaIPK1TnJtYKedVl5gdz95nTeN3bit+hYkb1ANGmYpfkg4tIY+UXcAdLxCbdYAqh8oDa4/iq+MWs
wot0YKHhyvQ2oPWmPEpPsI2eMD8O1mUOhUWp1EPg4/pHSxdtyuk9Sxbl/LWMlqtCrTreSWl+AKEj
BuqzWRBrYjGeF+vqDA5/ss205u6y27a/ZJOg+ylHzqZHXQTnKx3hOTQ+++pRX++zanCcKJPKAoVS
D9gOdOi4g9yzPx/Y5xn2iDGOEoEzaVvASF6K6Ldzxt/jT3E4zXyQ5HFJtGgjs5kqjaFyLkjAmM85
LZ/1ygMt/Gu0uXg5v4K6DOqkA+XtLsB5wGHXBEZFjWSQY47UCm6RXC68p3q44VCr5sIDFTtC2DvH
rMY0YyxZbWoy0WM1Crp7i9vdDF9sG80W6eSjgJWYRUbK1+Lp1qeqLGuHNSUEtH50hqIByyGnDY6E
IOnL+RNba93SX73m/9qOPpF4HC4hxrgPbnhvEfMaMXg3NwwAqxlraqI1XUR3W3CXHf6kAhf918gY
fbgmroU7qyDSDFjzD9aHEPY/hQdnCaPB5AZnI+G8OnXboGgbMjWye5e0Oqy2b+ZWTSQxkdqW0W5p
GDp6ggoLLI1NX3oskQEhXfXZrLkUZKkGy2SY++X5fsz5cQOp2MEVgiHurMuCznvSrN31yBv6v2WI
kji2mTeC6cNiKsiRERCyoMQl152gp+kWdt2p92et7sy8g+vmoj1DuuuUpbv4SXFLPmSsnaJ9haF6
YHRqS+U8SmDtcI5fvV6VDSn6e6YNQ6pQMRbaV6i52gL6VfdZo/YnNW6AE6zxRS2lmgMDZgEYbZlK
Wx0Sx01AaxPgbnHKpIltjfsuMeuTO19Xcrzm3ItbEMN9fwPiTvTgiR9RlwOYqEM1EAPO9L3Ea/2g
e52UFeeY3VW8QuRMb660PCrj8UoyIwM4pU5y2LSq8ZCCFAPOce4beKJv9NIhviSb25jvZz3zA1ws
3IYlieNN29SWiiP5GzVWD0CIVVXf49u7hpwaiUVbqzyTGe99GdDbeofdwN/Rpae1yR08sWk+Cht1
hVrD3CbleXSxkAaDmPweMaFChE7J6SWa8n0kaUTzaiSmX6Xxm/db23fBW9wv86ymKuty9sSiL/CX
V4s28ydTAo2/DtPmyF8m7V6FNthM9RbgxaGNHFfvjUeLb2/ZwU5Fw+8MEDEtvFQoee/1FoFNYR6M
sI1VBcAM088G7gHhn2uJQWfwV0/gDxXy+eIfN1Sp8GvGofVXxXp5lv69CA7sXXh5QSzws9V/T0JM
N9ReHYUzZtTE6nxN0amRX/aU29gp3AO51QIVg9rYvyyzqMfr/4sTzoDSqVeikE4kFYhcSgIzX+03
TJ2B9Hsdsv2FxEHe4DWqZUmsH1G8I823jat6xzq0Q5olHApbhKG+e9psCe0k59cauO0glTMOd+Rj
n7PdEAxLSQExeKNyzNWQNVHcfUe8p3d8qKB+87KgvzpqKiLN/K3K323/colwl4d5mvIpQxqBQ2xc
5z0q8AF9ZV5dU8N3SirKOYa1fMX/3gK5akCoq51cVnuRFftL93Q7kc2MSAx8jn1spX2JhjLT/loO
NFbshL2G6YA0iIFFyP8HxPfsEYbg4tPqGjdjgJzlP27wLxEGJ2YBO0vD1V2Ox5lE68oLgGgOOW9l
qfdsXmMcWRLNGDBivN0soxTMEOI4J4hgLr2m0gcQSPrFbrfnTJFrl9aXqr5tJm/z1G1OOclds/hk
LLEK6vGW0tSxhiYBzFQsQDH9Jel48q/lfcvWESSfRin1354kLKEEzvu/G3Os1rBp/hITM8cPql5c
Ifi9R8g5EMuwwLGacKSKf6uEA3U6zdehh59sr4btP0AV3d83sYf3YXO6KxPGHBu46+2K2wm7/9Dq
s920RhMGz3NjucOoybAv4j4XU/HGdxGNrjK3EFU16WmI4ZbOhGS9Jqb8K+tEEsUCWa7hVSXJQvlR
32MYzN01OAaZ5fsIak4NdkY5LVa98gvgaigHwx2N+HfTjmrDkNVqgKYz6G9uKm7EuPuJ/ifZ7RZV
AtIjF6qowLxL5Ypod5rBU2nbbatVA4lQXgkaSLSBURf8gMJ6n0Bwl8qcmYHldmbS/wca20pXQhB2
mkosDAD6C+FTRnoLVoAer91sD+D538hDQtHq9+sIZ8yZbjPjuGWc18NdXe/TOPtlLEamCcfJjMpo
Om2hrdJHW5mYP6aKCu3HHfKPMsewyESBMWB7SklZxWhGCA5vI3MVTsqDiLRcc23rWN5Vs6ZVsDOt
rDRNFleOGC/1XhbkLj7GKxwknYMv9gBDXYurvqhheE4xC5ymi2HOmp9GErCYY3rKFIswsEwE/tuv
1Sm4JErg4h/SvY340wqBW8b8PhrMwsaoKqQfsIUCbZHr93Vra2Bu39U8m8yLNyV+QkCOFJxorkei
goG2xswdDEsp53L/bsWgvUS19UtfUWThNPxHv6mRSr2fotEeeqie8sjmHUiCkSpiIZtEO7Ri9w4L
qR1tJEC4fE5zFe/tynYEJVxlK6+FO345sUxdBU1bzFbdnPed9lyT+bxCIfaAAxIb6R/hf2lAS5Fx
DjPfX9ReiQbGQ4kIRULke64vi+I2UP4UnFqdVPkYy2F7pxgauze1R+vg4SneHdHZ4aAjIJqlJNDv
9ty1vIXJ15bMeeAoL9aSeQuwTZIhTbPMH1PedAej8B/0uGOGO7sY9Rtqc0zrcdUTw5JuSou4iXhd
ynRCqoLXC6FDXPJgj/DoJ/Bfkls8RB8zbQ49LFRfOjAL8cg150n6ULxuSc9FXqrlRBVL3qZ4Dvha
1f7kvsCn7SusdEjNU61/rkQPQn1Mxb4FUuYNQHpSUEyT2Iymfjx+GOjoNTyo5hip4s//M3vCdOb1
KH5pKL4iS/hk+XJUtoKMRCf4VTo1PlYpjd/MO26eKw3uGeTOAJQkt3Ak2puyamBCCjbIKY+jat4f
PAlL1AVqPbRWYjTrpL1CS5J8ZfB/vVBf8v1uhdyIzM7buI22T6EVpiEuA7IqzqnFIF31q/08yLml
xCbIBwVJ1EmbxoTxykdNqH9h6F3j5mO+hWq+lhWBfK7zhm+/scdPd/fuOdR8RedgOfm9O11rByp6
EZ6JxEd3on8/cBjNn5Y5X6DUuTT/aKlm++iJjeO6HX06aMhXSmCYfzKZxerPxQoezbsYg2oivG/x
soWazGkAXTJrtpCIFUo8eixxQA3OS3j2X9Y5yFGN61KBYD9FXhhSJzj4fUrab1xFy/NSH7e9C6Rc
7JBwYYFidiag2It4ALI7fuifr9jl32FmJG8CSMwnAiamnWwM77La5DzjZVkzsAptBB78ogBGa3AF
gJYIapPyaGqNbPW0OQOYuumVDe5ffLT1sSS98Zr3YcNeYGiItzzrC3+KBBE+48xuSop3W+gHEOeE
ZoggYwnwsKs2PIX7cT44bY1lfIkIkvlgTxv135HDm6rGUNUlmD29nI77IFl+Ts18GPzI/4cmSaJ9
BKibr2/eucHv7wju0Eoyfy4Dp/GzuJRs18V4tjC6/ZETy+/6gSoiHnwKJV89Xclbv7+AVG4cnOYI
7utbLk8zONpjfu53JVbjs+5JJNypkhqa03Nvl0yZnI4g3128yf3NuG6TiBZD/KFUtwGSKnCc+C5O
7slWeYi6V4yYD3sQbHUBM+IAYnqYzYIOydbITbRG8pIJ5pbIA5ME+8mkgpZbvt6dcdqwViAtIsjJ
WiM4tMjAhlqwDfK4K13Ths4rBSbLN3ZJcLf8AIVSwZWf3QjF6oG/XWA6eEDY/4o5NOoY2UIvmg1v
cy9/svGIsG4RDIlPzq7fN5VD6groyTbI6Hbc20tI1dX5cobB4uY8inEjfIhqn53+2ytbLLv4yTOd
eXx1rtYb3Nq90E4gmitQXKY9OVLta2XT7iL+j/UaYuUY/vQrCLk75cnQ/oox+h27o9qutNsSIhPK
qiNNmwFPrnN2w1B/j2rvEAswb+JCRa4mNE9xi4Wk2E8R5SfuWLrVajfz+DV/TPd0UgWDRPRHIX+p
K5g2Yef6ZyEBkdxhKgQe+DvzOmn4VrQrZr7M9lepopluoAssADF1+LVxkF7+dfdIwvwXCs5EjF85
HJ32pTRyKrxj0fSUoCyz0Szvnh1A2HuOtG04JqfLOcGYOoxmbXuUgXbt5M20mnLftX5uW7bLnVc4
eNqKawWbImaKTtkBjED8Yhq6MxAck4y96LG/BrSyUbzs67MqYabi9aVPp3Du+z36JiaPtRN33qEE
Z8aUUg5Arg2dCC502UAsyLY0XfLyzh/ssELct4bLP5zMkp0dUWB6fQySO0Mb09njl63CxaflNai6
/A2ahMO0+wkYJy90U1frUHZFDlNeX3DwJ5zH66ST6XDW7OUc/Bn1fkfHCzFMFJwsnrQSOconl2lE
DH/uAR0QprY7lL4xYc7BaXyglJEfsc8Wz9+2mXhxuwBsTEvByNvBFbG73VrcXUWaqIpL3si67/qx
Wi6Bvo1DxDeoB0bWoSIwy00MUo6YhuN0Sxi4B2TZZzyYEMrGTwC7cxsDtVqOCzcbiDDwDQTei+oX
R4Edcy7sghKj6YwdRSqAhXJffrbjgcY9Dr3rd13lkxIZI0YL2/8jyEnkKgfVLdxKaAn24ZiJm9k2
vaaslZRTnq2R0C0RnptmKUh1J1npphVUnKqsRo9GeBQxCdmUPRK+T2S+MJc7QGjp01DnxforIbuI
EDF7WNoKCXc8+2YqsiS8hb9HuXIrwGLzoaxnt7QdJKfuvbGEX5TPohGrQ0WEltVXP65USqhRFMKV
X9jMP8VSnkVzsZs0kPI6oS7Lj4lrFqKOLjBtknKhfKyOni6ImBTmORHIfjFH/KJq0lwSTGKFbw+Z
HZJ73pE5TucTlvJsayXWgtI7fKkUl4o48qfdEZ+6sZWYOjYWrnS3exbQvRmvD8LKjuQWJXG2uf7f
60ECJqjeDiQRHnasIPMbtuzbtzAeS8RAcUclFTmx8pe4erIATp8s/0lrqMAhxDn8V1XW/8WjvQ3X
KxKoJe/xCOyNvl2xoHrjagyS3mpAkx1J8OGxAG4qlNKffKR7KueLrAtg7ingit33Qsxr4Be1iCbc
5oE2ISlX1y3Ieec6rwIYpPRFf/EAcTmW6HePt8Y7QLgYLMiN8OpUQMkhM1y7BLT4TamHF5WZgPPn
bI1nkjrOi8yYOqcr6rfRNcNnie/iAd4s7aGwajrA/t5ld5lTDiB5RY19cLEU3SOfPnwDWuR4H5Sl
eOLiXvObBDyHIbeETNuCFCCZWcumNWc6sKm3UH1tweoXiBJVwp/HhYMFEdlIX4t0xk/O4InEIorq
rVp3svLLsfsh8j+/B6k+6zs5M/Tlk8qjNAPcd3g3+CUbr8ft4N9G5qDVMIdkWqm7b3c1liJP2n/8
YZDEvjNLS/a7iC754IzIxn6MBn0pC4RLgeAYHsgqj6YX0W2rIffGrTSn6yEqSlgDeGVwNQx4rP9a
z5G2YmnmngP9h85BJpI/ocdA2MqAssSy+YB+/4u2Lvyp74SpWCL0uuUrDVyPK/VT2gX44F+rpDrO
7whkPesMAlNGWreRGgi2dNys7gKX73/CS1BBnUpe9bY4IwzuLk89k5X1KfGEbgLit+6lKJeFeA8Y
KiWd+TISJlfRt7nny3vDayFcfxMOHz3+8MwtetIDNiBBOgzkoSXO7htgZNjFo7zF9fO2cHNZ77hs
lKKHLgh0ZTjJ4UDCRrFpZPVIXyNRkz8C5M7wu9Ak/JnQtvX4BFmX4nUsRTg9HIXj09dxI49tn8v0
nopfikEblsE5r71EkZoRvHiNuy4XI27tsbIVWpOpvTxIyntJaVY0FHbanATNJC4Bzzz2QGwB9JMc
LF84qrbsyiY37I89mKDAFNqix8PH/5sao3uoev7e5kWDwbtQBUzRzr4xJiyakVsOgM8JB4fspp5u
lYfSzqGOdqFO3HboKnlStN985N+WLTtFhjgNPt/WSrXwcjtc8w2CAkFqetAMgYNoSO/AscRy7KOs
5ZrfhjxrvrFsu555kn5q3HCqdQYoyN9YT66QM8iiNyqEdj+z0FGPW4fOcpXa8y32LKP2KdJwI5u6
26yMs5wt/0DW3D61eyxsvTQiL6dz3oy/r7pXLnOZ7gl+vFefbdmFmJPNz6GLoKqa0+tfC6V+nRkJ
0FQbVGfnLKPwi8K8UJ9Mb0wxljKLOxVMgI+X75VX1+e3srOHFOitGOILys1ZnMPFpPxz+WrCdORe
h4Dw9o+0rWUUOxLyj7q13vInbOWf9FuGyokx5U8BpCVV5O3XCLF9I22xUnFxYkKaW95aNGLxKugF
8F7SfDm+sqcB/QQYoaaGRf5f54Xrau2+/SMjSTCi59d7DhgL8P457YNVj5wLbJ1nIZdWLKIXsBH7
ayDHMeqRTpGShUIRlcrBrIdY0mvm9fH6JLWuqbp26TfQECb+Htl/Nondb0LHm1Eu1Ibr9cG8W0AL
nqZdUm3FUi4REWinc66Y+lGzAYYRMlTUL68bz7hVbQKHetGMZr34R80hhLTx5EGeHSM15GkvNq7n
y3i19zczj3iRNccPbuSSJHNOfp5cRYFZ9mTmsko7niGkfAup3l//wEeTxkLKBcWW26AjyNwy9zd1
p9H48gmp+zs/kenBvSqNCH+mlfkv8pIwesVX9rwaKUz8DNZYP1OmsBfl27wd6cbDVhnwXPh4E+0b
tjxGhWzZoQHJuagsAQzOHYXs3asS9hciIm1uWONiHg6BZGMJXt2I9IxXAjtvHd9106+TZFqgR+67
g6EedljX0V4s5R8rSpI6a6DMmvXwc+3Vfxqvf0MAygcjBQP3nLh5ocDFZ6JZjc9ACcTN3heZ+lKk
0C6/v8qEbRaIGy9MUzQxXx9VGspnhOmWNC2IU1GhopN6qyuFanrk08y+VBwMshKXpnaXyhlgUYB7
nq9YbksNhUBhsVe4W1q+BlOp+KFMh+UgmaZoMqt4oUqcSNH4JN8xW6ymXPGHmIhHHZbU9+0ce/nn
ZgQP+BZSrsYYe4hWFdaZ/UxXv1hEowMFYMYHg2TGXJlISRCwq7q83hEXHwbtVSAI53608SxasJUf
bp5nCEu07mm3EdhdSRrBw0COgYVM2e8fINW55WBYe3yngKkuASPEtkPhC++H5IWPIaDj+dugtDMw
2Q2vWLJFPKHt41KAqt4nGF3EZkM+GVwTRGmsxubJ09wbtCFYOODaJqTNBvnF9sdbc5pjxZm0sJOF
hKjfblM2p7xDMqQiuWDHnLQ0a6TKaBhTH9b0lNRmaOsW57f+Hd9qyh8Qw05v7dEUAimZdbTrWvGe
/0QW1hvJGi5IjbNcgEMdJvzAmh1foYxsrb8QiHk7yv7ocG7CfsjU94SyjRRi+t041J6Iqt4K1H1T
VArJpOEIZFuOY0Ng098edyPUTCPYZKqbTHMrukXRQlBr+XwzavlCISYlzAmG/Y8iZwiuDbCIrkKK
MHss8XeLUdXoxtSg0v41pJZniHoEt7hrHLfXxKrpNzsccICCYqwZ89WWFDB7gaP90oksMG+y0gf4
yEhB5CduGI1HU1WmhZFpzzVytNIzzwVPJ63EDMuV0OKHMCMKF0RsntZoeKOhgiaet1vBprvt35qD
SL/N4VDLhvmzYoXWdOKyk/yCh5dH0MyvONfpyb/37KZ8UO+c8ZbAQmLOvceeL95qJKK4xxthWZdy
fSQrcORaRiitREOQgFyosLzcw0ctMUNISjziE8PphgQY4c72Nbj2fB+c6uX9VDwuAWN9s0VcSsEL
+GwehIYg8v43df4vJizdSiVqY959mNyoubOHNatn1wN4S4zj/wjgDXF56ySfG1v/zAihk77sDxam
gfz05Nx9VS+HAtRr2MKecmbkSjoLWHVEzwiQ+2jVaJdDXPSGxaRRVXV+lfmgwHY2qw8Ohg2JatVQ
IgKRuM0RSVEcvlt5oCXXDJBIOUlQzcht4F85NVuJqfhH/ahmwWCYMQ09/5j8c/HKE1/6g6OXNHOy
mnlunjHy4SdFQG8oyq/TxSwuYcom/iKHwlL3vWpNjT7GnUwIAtQ9R1QNiT+yj8rjBQxzG59c9fnf
wl03JSRtb/bHIb3qYjNuWAu/D0IDN9yZRFBMed345248mrxl5ZfcKY8cOo8dO9H7t+sbqFIWu4g4
3yzygAKkKzp0guonzwWsJRCQ3scDGXA6NGWtyQn3WueSPtu/TrqXfNm8TsV4YauGiiq/OSMG8WIR
bbh6zac+HN4z9pxw0iV4NK3swYtpJBXrUx4+dt05TSNUIvkCzz6pd7AEjZATvzuLIZ3Lu5HDidPI
f0wLUUDDkjd+J213Qs4SZ0kl+eZ7ObAI7okZ9quifFr+YjhZlhMqwvROhZEd1/jdc7S4zYQ1CO6l
OQooi4mt7HdyYYg3qEwqNN0x0HQ47uKcmFQS/1HvH0aXdm+1sZqyyhHop/SctzoeGX513CU7ZMXL
5PDibDrXshgDH00nLZYsqEf5eLSlHIiWO6PqEl9OneDlzidMyF9TZRZVgukbG9DzQ5VpgZjDe4UE
wjtoA+b4waw0SvApd4yE4OsIk5Y/5ojwpS4yRHhVfWD12nn4/TD3qEg4lkjYMDUGseXQIWVVABMC
egn4QZS6dU/WKXGao7I12YcZmSxZchrDgV0xD9Jx7ZOE2Ky7uH3gT51USDXDpl4fpyr2Ixk5uE6T
PfihkVSPDSdJFCMTvUd7NLcBpcsJEiZtfAdnzHjny52+7xoOlE7oNvB+RLca7USxBELNnAhm4UJ9
xUwsEwzLXtdZZbWG0WAwHgtVeDUvrVa/s/rk1G0KbJCfkrOLGfry8VYc9fg5rr2cvEkOUQlJr6rm
GRfkha/fJhvyiZ57nx6whIudXO6bp5oYcNPBLkQ1w9tpKTCeLoBZI4sgwXtr1DdNW+Ja359kh9jL
11rr1P+Fp/wKzyg/bCMPn0M+M8hkQE54PFlYlcesa9WON7mCyaJqE2lx6nDHDZSB3BYtCudlVEMC
4HJh7eAIUjFInmly1xHSr3FxxFGadRY6cX7WiyMgoohxQiy7f1B8WV/LraiWDuAB5v/8TlQZDEhG
Qzyoimo+aJ62ziAMPRI7vLz3c4c9JSs3jGRtdoBMAaeeWdBVvDG90AzVtEuibr7poC8S5wry9unF
ap4I16CVpdrcU5E3KYvF865igUHk7S1q+xt+Ej+Z1k6906vA3dybPdlwrVJuKR7mLOKdXERmErt9
k9Rqjiijh2vLB8bIjpA1h2TKkTIJ6I0cxQu3CgSz4YAa9mjnJJdhKT1W71B1hbPJKXtWlE6Scjjv
a9c3t7w7K05bsapWE6ARknCbonsGDbuhtiSLX97oEBahweW4MIzAA9b2HbC5fbxQhUhT70v7uWy0
//H/J+u2/r/lDaDcqQmnqTVJECslA2moZ8rZeYqZJcMB0XM8jCJMvwQT9oKY8rCWskYYw6Nzw4gK
0I0RXhZGqM7t06KGjvOmvfVkJXmn+M+GU1fYSyDnvxn9wJn/Hct2R75EYRhORHOsPJ/FFaBEenmy
bYLvd+dWVF13zqKsmj4k+wLqsoNPbYNPuC/oJ+eJr0oUSLkbAWGmZRid+YiFKp6jMTAr5euNyQJG
1sD41Ev6ULJQ/Pb/MU6jWkPhXeXe9DW+zDdF+PIahEpq/rH/Cen62n1p2DYjZQW8Sqna7skqDY8T
ck5qVFXHokvQen30A+uxr4enCGSDUJUSb9MfBxqkOe3YC1nZU4+Fua3gcJEFs4iGpqaWXsBgFXXm
TLtjZDJkkiiyWsEILz1+NxKiUCUxQoZOLgakUcjfrjrcIomdqy7i74ahivrIMWW+OwkeIXhouOu8
05TM464yND+nbJa2lo18XB4/Yd8eLCGFEVUmhQcPzU+mOCXu14stzzMywUVtxJE4Pb/0uMxqcA7+
IRzHkXM7Jzved5rl3q/7dA6ACXK1jjR0SrKow1X2/3bRrnfAXLzXFpCoO3jrgjgtTBcHA8WeJyVV
2S7UXm2wiy/Z4FcWF1yJNILOvVN59VYXQ31oWbiKLaOB/vthDH5FL5pJ3wxabu3SgoDhhZU0dVIL
z93LKZ05ndMllCp25UCwciywbNNEMtGGPZ7xEiyLp1pmtN/Y42olw6uA2PCbrnG8m3ItXKNwtCls
tJymO03u6CTA/+ZtNYsVzH+55jqdoIh0vqt2HDYoIaq93rljaJ/Mz/V6oBMwPCkmvCxbQNRppb2s
z3axoAEriHqSQyrf0X72I9IXy7ttoakLqZUjGuuZ9U9YEs9cSDmXvy6ISwdKEnql80wCa9QYxp5U
Da2K8QEfdwm7JxAsoAbX6bdstUiylKlWj8huFtgpbE+Sy/khCmkJvV3VupLl8InXha8MOCxNHDY3
CQqELO6ctvzizgxehbNaQc4Kqy4V9CMJa/DE+ZmfGP01QWfqzzYEKFWb3ZMHRgITqLNSsoqPIi/g
oeUWPlHnJXBCkOufaamKy0uch6L6hrOcNrNjn+kZh9IAv2BW0GWaC91puKyi/SRXxbEBOkuFS83S
YxvNNO7oGIoh3ZGa+PkQXaoMd3+4BlRbDFGM09teb6gv4s3KFIaRb95jwRg0pLLkgbAUrzzMMUXa
6gqcw7qmrS29XSjUA55sBKYGBgbnmgx5aWHHyhha6ukqb6JWpDp32SmP1o7gEsI82VvrR/mn8Oin
iVCa1DuVcg8x0DYKhuxmROggCLGb4S3kZ6ymNU9Wd435UWsf7OeRcvxB3kfHO6zqQ1pmUdu11L0v
YkVcXtxgk0yWgCc2e5gW2hFP3G9ybN3o0StZW3DIVpWsvjt41On0SFBxCEs8QWeCPsV0Me5Kp4El
0yiyRiWO5Umxc8tKNzPy2f0pT5wXxG8v4/dqM5e41EiLxEKHpVwtj9GJIC6+nHfSCVh1SQ00/i5l
w/6IE+3ApjF6icg1QCyJOdTst8agmS4D5KwhYp3znGqA3OAcbuSzs06B+UJppLm+GtVXe1CLT50P
eL2TUksL7dNuTLnpBZtB5e/MprZ9HlhEvIKAmsh1EIHj/2FbofZrGIDdWpjfhXvjkUW3OPsZkzk9
cenl3aNe3XxpEUdTW5Np98hUzuNga8VE8IddMf3hlamTNyRGgXhOKtoQxbruRoVq/LLYAYEJEPX9
5gd267nWL4Miz3oMtN/Dk0aiSSyFrclq+mA+YVGMaiOVcKNYZpbBnm3S8ZkMVSvExtVopAC1k/WO
TH/pXKlkC2v6GS9c1JXoiygVyfgGc1OJ3Fae+P93XhvnmINo4rFBkEPuAgUujjB2wfTjzFrkZ//u
5kJfKrYD94DXQ9IQF7DTFET9lcOQ9YuUQE4n2F1uPY5r1nOS5Obwr6sA3lDRgZ4pCAVQOUuLho5+
/NtPD9i7ICu3DhB52ttCsUMnVe21T1pEige2nsMizUEvcBMvmFxsulNwLU1N1osN3bcxJZSLDDmk
oOIqJ2UNqr2LmawIZY/PUIY5y5V+p6aMwn0n7ItNFLu/kDFe+T7cDeiE6zYDHs2kUnSPzHjO/bGi
FAWgZmgJ2xrWDG578gj3JuM6AE/y2uOw81iB+KTcGeBmUDxNYSO1xs/fksDx1PW4+s6vGRbtcOgR
LchAEF1tty3xs0Mi5XQmJl7qxkt6uOyS7O6raycaJrLZl1bwB3H0N96p/lB7WcBZ2efLhmLS+7OD
w21ExAR0fjMPXIB2h5yUIRlvq7lkry0qoZwWC4d4S4+UvvWRHwqdACMHtMXk+zdE37jO+Ms1DoRi
I1ACk2cebzygRd9i368snymxdG8UIjqYttf+hh4Rhnn8eFulFQTtHlPATT2nsCaZM7OhJI9BXR0C
wn2e/u8R2jgPbsNVktTOEpN8EknIxdX3VBILNOdalrrtrC02XAtE4HAcdF9hSx+dWaXyayjle086
C5snhmpe1QHsY2GB0VNBhT/034KAlrbM5WrEMIDB58IZuOTcWQKqGB30KP7q+Jty4cvYZKZnkEnG
WCFLycDV4v9VKJO2WTpq7nPGkFmGkJJXIUWUNN/JUKXfgHP28KReaR8AAaZq2daklppoYXUakkrk
IqR8nW7I9eiJRBoS3vjsFJvg6tzxarUhQjHwFojGj57FbBSXaHOhoMFjmxU/R8QYX1xwnr1tftpw
n8niS9F17u1568kGGt2TZVu0qJDe4Tirzsqkthc29CzMM34YldxWPen+EGk2I5rBSOLp1tiuP3QL
GG7ZMGQQy2WU9n+DLg4SlS5cnmt2LNiIKOCjdxpT2xMPTTg4QiTe6rQXZpTLRPXZuB4fDCDQxv4s
PS0dVZfd492TQcROTvz9wqNq8fZwCmXfzl1E5zl2IZElPDautAYeALIfWsUZuzHYK3HyLXI1Go5M
Hwk0fx2M0AU7XgSGFV3lQHUWEZbiTPgFPy7Re9VWWKIHTa7nxiiC1muMBnPihMr/FylvLTdfO1jz
dTL+jMP7CWoUpcO84NN78ry5sn8nNdSjFoWOBgfsXKfsaIRY08plOveoFIDt4/ar16G2vUXB/dy1
NNg/BlbQl5snm/tP00VN2XUwaWeZ4tHMSx3e0ElPnTGzX2pu/wSZPWiP/dXY0qYV4dhDEfFD2xL6
cHp+yFx693tMeMORnVWJe4otSSE4ITWMQKlo25/O68EO9LZjgNHIYvrmoXV72c5L5Ypepa+ECSbv
bVeW8kB52YuhyrlrtPC6s5vrMscH+UDUxlgCG/jUdu+O9A/spbA2DogXs8DybuQZe64P+HxHY5Vl
tltAHolm27nmMXWP3eqteGe4Ryk4sbBgh/k++Ik9rNsSmd/WUhKxwWCcZ8F/lVpE+g60fRJHY1ES
ThgVajQNqIL+DAIcCOgAANk20pt0LniPTpBSRI9l1JLlqkRZEsCllTh2IFtvo9WlCrP6EU3+/gIn
Cjv7nFVSaKwSoVDWWe1v6tKNJYh1Bowb4ae2i7F7NmsoVGSIGn2K9ubkmqQ+KZ0phcVuJqxso0FV
4WtWkb18q3sPQe400AShqLvK+KrekX1avlVs2CpQown6EWj6fTJThm1e/ERoAlo/ztuNuuXg6iOr
8rY74HUqZngRb2A3ev8krBE462DBG1F0kvilBUgPpzSvd8QeBfp58k8vOAlIXHBEL55gx1ha3Baa
ne/q9EoJ0TTC28sga8lGea2GT15o398XA3eeBrqSgI0po5G3RqehB2h48bhYtm3oJeA+s4qHdkjG
VQLygLGYvF40kgZ0MxD6t2+UpQ51wA74Ij7I0Xhobn23Dp03KYuDgjlGthONyPGbIVBT6NkSOdLW
D6pU8w0rmxfTa2sdyKZRIk8o78AKLMlW493GqMms6lYb7ovfRfDyHQPxeSrVYx+jpj+ajYTM6Rmk
us+dwhr+JBmTZTfJbIYeJuOqu7Uws27hDGHUjYBCWL1oRgADx0KYJLSaZ+1Qcggjy4VZUw15Kr4U
8Lywqr92q/DDrEHlDliRzHiM3gz4Vq/Yos24I5SAy7nJFldpGLL8zqWRJ0dj/7ItOGkH2M9Q7e2H
lr3YeNy0GGAYCe0JmWzqUBUzdzvElE69OgdEK+Wk6fWxHHVmALMtoDbf9VldEbneqGPyTHixmTCe
haxKS2fBzj6A2/h5S6mJ89lbMcwc7jqpAiU1i3b+0BH7RF5IY5NGU4OxEbFUtPojSngbiGCjGM9E
G5jIt7k78ULdpGiy4Xm2qzj3EjWYCDPj2pXnWd4TzaJKSv6QHNbbGRjUg5jEiLTyuxERXoQ195Yz
tJzFQoGyfPaLF3xPLfBYUYn02ksdsEnusaT6VMD9XR5Ch8pHcWys4a/pnpkBRWuIcvK/Xzb1EOql
18IR5M6d844i20A+mnWL3x1JQZhjwaG9AWoMBg+7BYM8jd8ViNqmWLtUnGi+XhKdQB3h/ats0wIw
g2V8Wb05M5IMM5m9PKqrexuFHKAqKpKpzQx7rEqhb9+vlPuYWPG9JLRbm9nwRB16t2wjostQfG93
wQezVC+ZtC5KXUVzd09kQqik16iADk+xUAOkMjJe92h4nBx/h6bfvPpPRVLAChobb2uUqTSMhpFA
aaYpN9hOfqiLmVTUATY8wXZLxKnM/P1gnMuu5ioYyTDY7+0dhD8PhGsUccgns4WdCoetvn8j1ICU
fiMSoYq5zTXms/YwVwQnnv3INVlaRdrEx/houUoMru4h8kiOeJIdXxXZME4ws53t+XHiO33f16SE
ZBoxf23OFnnv15iBp+Y0iNg1oONs8pdJEnVDDXmnVN5eqq9IjimZTlEPCFrw3ckR9ZIW9vP8TdLc
cYezBn+em+vBijw/fdi8ItV0leSV1EJbqcOj+3WeIV0QlEBvA36vEdnDSE/TmZA3WqxpHsMnjuZC
StKUWbQDHHVPF4BOfkbiPmCKgJn7RkVTwUXu8y36wgEkahF9IK4aFunz59YTwFgzrtz0x84Lqrun
az/Cyi04nnsNpUntja1bT4qvdX3/O5mpGqKAzKslp20cZYr6o/Z2w41rj/SiYoqeW5T88ars0X+8
SnOjWkHCS7d60H6QtrNUH6zJ24Fm/SjKrMxxgsBSEZotVubMRimwh6ZxyfK0ocfU4oYG6dDeuAaC
nQLdms7KkB54q9r862vBeZOS4qqhqdQtOeuflsXs/wLRDE5fvWM9Gxw7vxhCcBmNs/pKWQG87vD5
dcjeenvy15AH1T9FBqXk8NAI1UiulIcXhutjoJI5D6u5WWZolsTsJs7g5VjLxHTQvKRPkiJUXhk7
kuOv6Qgg8cUAVmHWqv81jwnSj0WO2/J4S3s20BjPF1dCJvjc+fEqqsQRDY8fjE5uE0JX4LYswqTE
cgx6Qiqzt06z2lGBCyUmGVLyEiT+KaQ2e/SF4JoLIHh1yFjdAUJx0I6JpdKqKuS8Op3vyytUnHm+
PqoAYDmnXrcrSlV0h7vxzt5RYaF0EganHucL7bVQ1ppohQwsZfTqtR2PjomaE6s3ALrBMgwN1SxY
5D7qUOJ9jz4iOlG/jYNRVsZsdvB7CbtlsSv1O33YjVfGJR2itYxNGIVNzpJBL4RHUKQC3ogWW2ip
JYulOmLCgSeJdQr5xN0pJEYcmHkhMrKGMVRa1lXHez2wh8d42RoTvYyKhpDrlKz3hwc9jdJ8eJvB
kAm7RlDBMY2Bv5R45zYiD5Phav5vxHfTwdbFZFtw3dg+eDCLXL1DMdy8TVPwTMahzKBaR0Bz52t3
0xzp+p336AODREowP/v6DZ9axzhKO9RnWT8zsdeoiSdMYDhLta/r1vRTL/vsAwR/X2AiSGo9X6g4
Hmp7+rKli9+mFQP59KdMNV9IX5Nn7FABRZeX+p3gehTcBwp1Ebc9JUk5lBzAsYtiq9I9d2BjE0lX
yUZ/Vax8kBAztb/D8UyyNOzSWnrOuODi02EJ4qlg6kgXfPRLAbJ+u17aXBS1fbjPTmg7fVickpKi
ILOy493TxsYEFrQj0nR2UOJbBS1drn/HIncbHJkcjG9Yyq7fSv+zVUu4d4/MjEshyeeV6d2gaOwm
p3TNkn0FMu1y/FrFKHYUpsKgyx9p4ubTKuHGRPcER77GLvYXhSG++8FqSpbKQBzgFBoElnfP0PyU
6UhpLPqkgX+MBS5WoJEwhUTj5oIaehaFVGf51kJeVihwL8KdgF9oquDRF3e2ydbFjGz3M68+HZKI
lELO6pQeVgLxOuhCsT9Mr8gjvSRmN2Ft8bCGeitD7X1Zm6/X5DTscl1cZrJ+froGU6NwuUs2qtoo
C4gyELFh4Mk1CgGiBVOvZVGrbQ4nPT+xBQlH66y9K4uyEqy5cijBmfBogZ+Y3kHZPOAMt6O19L9D
HfQl/8REouW8R5rTSFzYYQOlBUp4fTwlipS9Qro94zwtDHctNBC1bfpm3vszVBU9Ou3/FbzzrQYR
TJMhHX4E0nEtBRHgrnjF1YSxxlVgnZGaFUpjBn1QPuAUJolcG/QYzxeoPc0TVfThL/06E5Vfozdg
LnKaqpMC/VF5vY7EDZoKEJkl0BB9PAREIfQlJiZpeSsrspJY4w95NCWAANhqyE49z62HeJa6/TrB
iEmNTQk6GCEo2fnVJ3mbVzPCMFNuveBENmKd0YL/jLp8jOKVMMLsC/da/9h1FfHKg26RCqDIbUyy
kNFqdPHMfgFGm8HA/7lmI5xap0MgXUbPu429L44jZ40fSkO1qhbbc2YgUwDU/LdDjzSnO6hHgGyS
r23v8i7LQu+yNmqees4dDcy1Ek/X/tuQqt4LvyjjvKPZoWKu/TBg0wO/MpSTjcspJHoIQxUvbTZ2
GKm37GuWZt6dJgTsCHCHYrhyoZ9NCQNEK1W5/g4u92bii6NlEFiq/nSMzZW/0MvgckN6ONgulOUP
WLAqkWbSbPyb2ubIbm0OMOfFltHcNjn05/FT5gd1rS0VPi5UpakwBlh79HpufwxJtgbtkb5jy8Le
7moTkaXVkX5X1YXBKudYoadcHQvy9bPP9/5vWr5vYb0l4qDOl1aPc04276UTYTPibHmsEzEi7FwY
vo60IkJ278TW1mL651hqTga2Qa3O7F9zVaEg7t/nlsueIcs59kAKI876jiemD09JS72gDx6t35As
rCu8qRuT3KKWNKDUzelaQP+MuY7rU18uLUyqnS0XlCVaQL9/dGmnMO0i3gRENKSXSulQLXHcfHoU
ts7RB/0EPiRmSw0/6baJHweKk+vyJgH67oXCM1oTWcygFCry3DvPTpR0dc7vXRHHnApedOdYrAOJ
rUchPEVRnFv7imTo8bZRzWZBgLJ5T0r7Bx/eyrDgJaIUcm0pRhTwZhLqntGE5yzz5GReTQ7Lhhp5
M2JUMFn62vQXpZyrvSu0hS7rLOkEPOpjwQZAql8OZgx+WNr/nGQ0U9kGUN1hnFrL7Jd1iuAxL0J0
I69OeLU6EscJO3CiiGEDlGD9506SWWsZqSvtq/bVOYoqwqx2gtmCv4lPOf/TVTRH670zz3IFk23Y
ij6IgdWXZI6+Vn86+QwzTaxDnUMWWA7RzPJVVU7jY+gMwTolweW4UQnjx6q/8L22gDdqgKOVMe3a
E2dYXNsMbUbpXgEmdY5jV98MZtXoYngfT3XOrDaAz2XyV8mOGcGP64BC5Oqdu6h3oj49bI4R+mtl
DblVFlMlNE/jlUOA3TZbwA84aRbpjNAkyuJ1PQZg2+j1k09obkAQGXWKudnP1sVghALf9KCMd6+e
YCJhiW7nZueYBWXAnn+S+UvUwBcCysAumVrFDwXvHg43AMGX1LcqNplP/WQjzM8kfiO6ADE1RBww
N5ifzaI/Umf42e7Q9ZF4SuhdHrnMMcJReUrc4ddpiQOONYmmZT7vj+PnPfedSRf79fqIJ3Z2g7Cp
7aBsRviEU4NyiYbUcsBn/St5JZfPdoVGWbIcbfkrJ2mlsJOTNHrcf3MtktOzjudXRb6DRGHZy8K6
D8mU1kkO1wAKTxa+MzeePWec4p/wM/WWacZ2MnLpzWXdKK1QjoWdjEU5tN8PZiAROX84xRc7D+p3
qpPwzFQ6FgM+lsuGsli/+oQPU5COSLaYh1G4hzmkl0Vn4843JUhb24O066Vy19va/PZ4QEPAyhNR
pQPEq8X+4cAghLLZcC8i65PHwpy58ZRGaxKxglgh7BcnxZgzqX7jZvbfMVlEizrDv/0U3GEjlUyB
v96Vsc4NzBKTefi8fcrq/b4jbplTYyxqxLQOisNQLz0UQUltXpRs26Q2xtDsB8pSUCrtJ4B7C5RZ
ep1gzpTWOe1qHuO+JNrYmeqEvyxD6pC4npGrMoEd0bBrKpAcP4UxYhwbGL3pZUF6NAyLmYtDVYng
qGa+LD2tOqCX+dKkExrxDqjnNanBnd8iIZVeC4gbWYlny2eIlx/3mbTxg2M6ge9MQYEclAIpHuzR
8MQq4mlQVJaSk37Wumzaed/DN2Z/+Bkq5YOK9kmt42b4qhLi/FNgIMgQiv+de1khPkBSmEz2lmxi
Zr3sGMYZl90ZS07HI2CPVSC1onI/o9T1Jo88lddg1ZWqAffSrkPyYtLiLusX8BhSr98lbDdTckPP
JHH5EsFGaC0U3DV+27GBFpDm9C/JeTro4kNvEPSckt/KMsMs3vd55qADd4Rx1CrnQb6y/QKu1QYT
NWB2jVavtXy32Td2G/2NnIFK4bOTbYWG3he3dB/cWd3hEMPW3cwN9i4dEC/2ViiNplY7vwnzlr9r
+VaYgQB1cfOsQKYzg4bXvlw+jeqBIduXexuWKpNo6Xso/JAVM2WMkn9FFDLzZ66ILVfWLR2JnkXZ
AHz2llgzCcfuRyGkJL7IIT397ZZA1hxxplS0QgtPR1jNjdsVQl/DYzVau34HofhsiF/Vu5G3GEpa
UJiAj3FKwfs67vxFdAQNHAVrCUDgOWpgzddoVJrcGpM7bmAYyZcZOnCuoLz+A7HlQzj46Q8IyFE/
8mp9eD+WD1Ck7nKKy+Yo5y24i58Y2nkiVKO+rCB9LBiIBSGL05NABYJglCrWZgKJz92iysBiiIJ3
5rdobgz0NV7oH3gDASZm7fDyl0lXzqbDXRRkRzLcpckTMQ64HWwYeJFxHX1R2oNHWhDpcZLzWx0f
hq678Z+nxmwGMYEuuMSn7++RrB8X7DcD7QRqV4MdfRQzDSfIvaY+sXRBU1EPL3f72QkeJ2hb7eI4
Kii/ACFQKmzLL7dJVmEENch4L3akKIDxdBtYJsx1VGx41U+1mh+fE84GBXj1yWZtLbdoOMdj2rLX
4+uX7QCj2OpQklMy9ISUTBnpEOEu+znx1+iiAVaJOdTJM0bPQpBH075gOcM6pHj1aeSp/dPkJ73U
0IbHQGtU4X0aJLr7xNGgREJ1hVQ0UahCQf5dAE+fPh9rgM69OfXhAmVKkQOYhxx6aiE4VGhQgSN1
7bSZaQaFjvACPf+eDYG2C+798z8AJIT7NdzGqBirFE2q1BG3UgSerORzgmBENq6eCrglKUiiSR9g
qHPD3syPnG25MJ2Y6XC+kcK0S3nxa5xxaCwd9IraZr0VQqEoD0g1PlI7p4vj5zxQVznh3tLBX1I7
bvddD5iyvOuudwsaC+y8hJJ5Q4TarY4I8MRGkimbPMybGbY1YtMAwjwTuznjKYrI7vrd02ra5Hkw
OUUz99SPdalqVPPwSo67GuQoDJ7qH2ehTjQe6LoztFOE4jNT9iA2vQH2hC4Vz4wFsASRvr9/Mk4C
ElVTJaBts9CCq6IW+9NzbSSPFabBkPVChA0fdLg8NBiDiPoT4Z6YNvHk3OID5PiAoFr7koDvFeA8
NVkjq+9e5eGHLyxf2N3EhsC24WcGy3c7BQboxXSMa8UUbU2AUbOyyr8Q2flzYcFygmGMNs2wNuSW
0knxsdIH9thwvd5wSJIGAKj5hUDnLhuLEnqdR4XFfxeGmk2VUybmWoQBs4j2cURATlX6ep7kHYWS
D/el/mnIA9FdfRSIrbcu7aVRiH9W3/1Wa7YkqKMMfNv564Xu7QNEx/1Rl8STzdLHrP/xdU7rDRou
zfASiCGQ2ZJ8+Hq4mDqXjLDwmlMuFkhFXPtYSJr/pJiDrStShRWrOb9bUr+6d5ypoVFmXAzhNnp3
bFNc9VA0dqypLIPdZpiVryY2VvUCOSUgrABBN02gDRgmGQDs7KkaTg4h5kQgcXbyj3u7tf4i1OYZ
wln9aeCYLcDyslESV7MtDvjXkPyW59WQLVmf1JY2D2hKmH2QsY3XBGV+8zj5GXoy9omrqbxsAYwi
rh+1KhLaBz6ATSBVypA/J2YxslrWLMWCFO43XnCwz8PtUJlbQndQl7n0lnBXn3P+8/U09EeAseaN
mEIJxku27NN56PFB4sXYQJJ6J7yNtLeK/kx6s0TIUSFash7ba8ik+PMP/RORGtaercvSPWMWi0nT
5ttV4yvweTZVvof2kpaXYpwKK7k4vlYGKQpY0zibBdO40nZkQgEs/qg1s2ByR0mscnoGHGqERD4e
Qd5zc9RWqwRqG1DDKBTYSW28/1KMGT2T1nbvzb19soSp+uWKGQxM/Fxauyh8EQqmEzPh3ameWC5H
bXw6s731MU8tFLHUW8yklA6qvrczSIW4pVgNpuGq5Bx6rqj3VQ909uR9uRm+pCCS/vzvszsDI5qE
g29X2lH4nx3iwtixiaHI8eSmhZLdcxyCmyk77fZWIieNfc+C33ZyvKrrfoqMPAEjbhWspMnANUYw
q9MPhozSCdccQJd4emXEPOH5gU6gzdEPycoTZP85umS4xPCy5n+GGObK4HJHgl5PfKjtfh+3rKHu
rsVLSCwELZ24qEz9OXXaqMkC1dpuifLH9Dd6SdJNzmkrzJXWValosKgOyjz/ZhNt8w+dap0j8oET
3JaJxuOwsquDfSoLHNYe0Nok79zZ96G/CLcsq5cQTPnGZSt45wd0Hc3/qyNByL0bKPo+BHcyKDmK
cgPgk+D1agFXVWOVbQBtZqdW49qwAdY3q+EdCk5AJz9YwS69uI1nEDaYH+r6yn6wWto89DMu0hX4
WLrEYdmQ3O2deASWFspuDVURtXn1Wfih6RjwQFLrBisiUL4VT7Ryoy0OWKLUtJCOY+Pad/Kqs+kh
ZK32KPMwoa7Bqk9AoL/qxIIvgx8Xa8dnX+E1QS6WEcjwxlPboAMdRvNI+RFNDf38aorc9QZw5bEl
XvcW+yabMKUkf+FG8dz7qMvhlZm9wXWSvD9+sGTKG5aPZvAYhvpW95lXqXPwPp/YcZkSxzcnD7mc
zJLIFVWK1elv4QLqkr/b+oQ9cHXvDz6e24rDDOFQLb+kW1VdVYgCfQb47RegEjDzKOBW+/JVdygI
XcWAM+gl///eSHT3HdVOwBQUe5Kmo45gn/ytqHJuHNP5mbXoOFjNwxkXn1mZ2lFuJOS3w2EAdprz
PYhI0pIIv/piGsMHQ62dFiruKsltvP1X/D0KDrP7KmBAqdxDBdA6MzSQuRe1lHqmw734DD1a094i
jsyURaf9KUsXlEqGtiXxESG4TMN8zl7tjXpOmoooX3FCoQXMQSQQ2dEweqtxpYhxa6agruM6eGD8
Z4rlYw23DJK/5kZ6W1iH8DzfIIoxFL57cIAC8yCuK1IY0cpHuAa3/KXFSDvhyAzEVKN246oTbexu
O1uVCjm30Jouq97jRXboEwdb9xFNEXmj10uIasuW1yW+3YiSD8492r+PAyVPX++OcuYRo2VA+T8r
HRQmab5s9y5ozgJBeU1atZ4uFWCwHtLP7d7Q2YFD6Fml481qJmsvIGVssPvCTdeYn5txCHl5rgYn
LT2+yG9+dc85cvQ4s3lGoAgu4AtVY+/FrRaCjjsVkKkA5PvIzqYFxPPM4kFH+eysydfW9lRMbqK8
X9uhEJvJGSUvk+jSxu1eskNlFRk4WNbRfh7s6YeivHrjJcsphperY2jfYKIsIhsjSiUxoBx3Lx1k
8n023CnQ1pV68XGlGUVner3bAhDPNCqQqeXoiN3RimWPoQIJcnTcvH6QBQ2soWk2TePScbCqVFy9
qYstEBrEjGJXtUmBRxtcsyz7Zmzr/Bf4N43xl447pZR0DJn7uau8eUmWBXu2Hi1vKbK7NJz09drd
UvTMzpx1bBKzHwdmXNth0glLI2Gaf6i4ESowx8nu37RvMVInXSqiiBbgrfBghT0L98at/4VFJqw2
w6I4aSUrr9ecW5oqt8aPQB6e+E+h272b5Tm+LOOu/3EohkRFluDNAaWMJCK3Lkbt5qsdYaRQ5LRK
QFyVcEe+UY994fIrgduDTjrgWjx/11lsZUC/29SIeRcSJNR+zdCp934B0H5KUeEPx49RCsQW0H7E
14Juw8vp368B0t+NiemRFFNGXgboTkBnsSvJZjlO+F6+rgvO7R3erYPHcabjuEtawWOWVWebVy+v
6vOU3Wvg4lXdghFHHU9hJ7PJaqLeJIu8G3zrAfkZl4lRbks0EWGnOx589IwdGA3VvgVMXAdnHvA8
r8K9ltk8FaWezZxlI82Jpesf91EiFZ8RskmY0XQIw//cADn138/OZGrWlR3HeE7M8ijZ2/fvDpRH
/AMdBmJY9oqCNA/RfvwaxuS4B6B48l0zz64av4yjfzCe8nTfn60TnZr8TSTedP7/DqzpKBuxYqw8
jBNmAaFH/tr5qAAO9aYa3k9uO0bEY1MGkYn0V6svrn6F8nSLTLhf+7RaVndaJavoqLFzsUGf05ef
KsJ+/0H3PLAd1TN9TaxdqPHf2uvgeDHAIdBOWlVcA0AGSvLhNsofhZIjRPBKbwHufPibu9m2by2I
Lzn/0jFdO+2yNpPKNpuQhDd57zRiCxM3vcTGDcGSITsYRdtmFMN6iq2Kc4fe5+yU6g9t+lwvrrx6
/0zauqW85r3Uf8cx9kK7TNWQaUPhexrFyogt6CvP6PsUXNxNJkf/7yIgUJq00xGmGeLRIReoUyDT
ULkWB1CQ5s5eJBUELeBVd2abmhAcTnDFdTsECEk88OuZGAfmpxmzov3aCpbZ+daDUgdnJvO3gFAM
Wb0pgCmOEv3EfNoC84Z66luT0m/fbAc1WO5MXyD7V0As1ewo5lTz+ZtPbBSlZkpLAsNifP+zxxv1
PvFpFowunlKbHFU3tqv+zlcqSrA/hQ1S3vkv1roev/CrYAQz99bI1qs1LT34Y9NVJVF0IcMdtYXh
LkbyGpi1OM9+hEwunarMELDvgHSsLxc9PdmGNVJO9Pjqs4VHmTkpenh38eIScAf3m2Xj5m7CgM+/
8Cc3v/w77lEtndnM8AOIWdpjZelqEWmtGjG4EZpdFu3nwKYDqb6JubIVdZnWHN7ZBnZFGtERB/c2
EzsFflD22iMRZknO82FF3zrifPE6UR2WZjktFVdJCyjt5uaU6mUnzt8ThpTAWt8vPKlg9iA1rbCs
LTTfoMd5V0xOiLn1+4vK+rw4Gtj0wPAIKl8EHzSRpI1hnuvMnP7XwBtqYp9b46pAy18Gl+DRoRpk
93rpDVUFMsDoyn5myWMKVeOA2WfmM2U5TN2eibiYW4bJ45Q79PE8MDmQXNTi/vWLXdFe4sTjoZdJ
Nbzaa3JpIWOUeyWfjIbKXj1WcQwrpZHTjiEYctcu//PMT/RwhZ9JI52LRBfqj1CYN/61VH+60Mz8
u0FhSaqntQBqxKMO/xGyrmLP4RUNkDSL9WlMY9ftul16uicxir2kIfgNk+G6TiOR3U1MWkncvkXm
5nH9sKtSbkimLeIiE/6FxakOzGw5JHy4Vx7NZ+WZNOOEr5+Mg3lHZNwf1QwT0i/QMQEp+sVkquPs
7l0OjOLRlSiTuipwXidL8KiOKrehzLDaTxqHjMBm86SdNo4GVceYVVTw8a0qE8CICcE/G0KZE1rZ
sy8cvI9K+1U9nRfHK+mbiVfwgUhNZbaJI10RNuJI1mAy4Ef6NcAUIrVtABlLqXQtB1kwk8E3GqFD
NRRivjLiQjcQs9gHfm+jY9VhKhL4/H3JcO4TQCr9plLoHXMVuu2Ev5CzuxyqDm9K0aR57uwVnd92
a9eJrO8QC+nLvt9qAherV+n8ST6fAei+1oGG+M0lE8uq9B6sV8feH8byvZwDMbJvih5x+hFRCbUZ
YysPfOeoPQqiwXq6enGogKI9y0znmIc+LZbyA4blpvp1VZrNB8EDJF6mzXnz8+igs365/iVBwqZx
PQbcSdDFs7o9BM9+Bbe2lVnVaCmUNv30j4trg4Wf0/Ao1OFf0q4LGoRR+1TGZcJEsuDaciPiduSE
hV+E7GjWNz9ekXhDPGfHbkA+sG9Uet0NW1V7A0BMhnsRO4IeP12ZFDUNbNzDqCU1qq4chwWe5jRs
abDjlIZDjenZdoIDq+sxXT7T1zTACBZk9XIudP1kXFY+3/5/iQ39pWoJYyl+Zq0JP1KLlNEIAl6D
69R2UCoNHl25R4aXFaWtWrowRv9eBhexHCzicygSpBlNs0PbrVgxbrpJJ7uTuf1CjtI/gGJeVxEn
Y3cYFeZ0HbICv4SDVof/TbviQ97H6blh+HrC372jYTQa1en5uHVNtGfvzXtB2ZSUd0XLphugBtF0
qLWK7IYe7KG3tawhVyYz2dI5DWvtDDYbPnKVoKjTMzAWcx3BokwLIAGiyB9pAqqO8+aR8ZgbPNt8
o89aSPtJGxwJTn7DQNYPiyJ0KCf/Vg3eTueIuRyJO4Pjo9+wLEJJD/v3AZ52eVEkWelq2q8ppmlV
GoUicsQ7WsFnrLsCFoiwc8v02Gj/SWtB3F/ufmvgAlE/dvN/cRkbu/iSpXxmKA7j7dVXpBrMwtH5
kpwJDTX5DunMyHTY+GpheC71y99ltlV3QJD24SVZnBqS0R83MOYeueX8Zr6+5nwhVhehJi5BxjhT
VAEwuz82kh8xlPP+81feECaAO2sj8nvIpN0H3r2fWVC6x1treKFWkqtFuQIHWVRKjZ/4GVqFDhC3
DF9hfzOQ9B0QkCAce4cMczJInnI74is4OlxQXRbfkYWozJItnCzX1vW23Kw3Frc07CQb5bbiHE7w
+rkCZYRaz3oRK1o1QhzTzyPzbtYDUP25TR+0kwFUFFkUEX9hRCIioxaviP3AKapjGs+e7xaesS1o
9Xnk/Jc6x5wb6jKqkF07IH4Vp34Tmmipv2oaMruVd0BW1/OGpZN7IvALENG92ugaEja3U4qHUN/W
I9DnCml4R/LjMV21YAuGodfJ1Hx7/DgvZu879lwm/xwRYGsTHhqbRa9izN0+Bfkbbv969KJOiBdH
EOSEehSP/kA/BURJD5uAEcgh9p/TBZrnpmL8L/8u0coLntvZQ8HHfG/sguqt7P/tfL+Iz8oOIu6R
If4kH5dfnvTdqrLkgbbap6n8ozis5XHWsCm/lR8/lqOl0R2Rb9tgzxO4/FvrOuo5w42vC1ZMKtYj
W8d5aBVhugczE0wd/FL/qfByI5xccSqdDatme8qJHj9rBsOMLAe0QzVWNG96CrqwYO0zygFbEYkr
VCx7LiEVEDwA90r86/6vek2PEojLGN18hJcH0igfqF5Yzxe4ooKVXQ1uaEnji7EGbJLC+l79wAuT
zCWF1i6/F7m7Et+Z7Ba9LbIpO6+Z3hi1yuRYrQM61gibyQbFP4iHVqWASz0wJvo/PlX9/ejA4fve
WIq4IxcsHAc3wq4fVqiaYRsu+raR7Sv6IVRuGX7LlD0hnxRz0UAW6yy2tPMENlELtGvWBpAuAqQU
Q6g/h62sTKVUa4m4vBKJAI1Gp0tgV60QTdLr8DbOmeMh2g+iyxVpPYrAGPD8/iPJV0V+BDs4K4/D
bJjFoXTwHdb1shw7B0GmV5DrNoMVGspEO8p3RoKgpJl2xIZJYIJ/rCcatPezkZCGkw+9Un6npTr1
xwnyFi6QrU5SHfkgE9tR3A4VSxuhe+Lnz+csA939o3gYuyMgu6hYSGCPE0U4wdOlnDgBav7ixvi3
+sjBPujyfKE3ZGZVBuiyQ26dNgodW2pyxDlR6g4d8I1b9QAKGYrqcFABHjffR2uHg38W1MRRcEkj
uN3qRVijVslSKwjmOYsctRS/zU0PPXOWTNPAluO1MHXuvP5KrJpBfNJL2BLxZXuTBU5ji6zF61u5
1V946HEcuYU1wuuhHOj3dVLy/4ayJ/RNfLTBGOC/+PZs/+PjYEn23N5qdCvas0KQ/5jV5+iyMeBC
PkejuY+4E2RgZy+KkIWGw8UCDX2QffVE0BikenGu6Nf5uiz/i3TQPfiJVxzP+PkBItinZSfVVsk/
w8zYcgbKhJa97qJe+nTq0nngdOsdUXP6FrsbH7mSXGqERLC4CYYOXD0IEakR6Jr6l1d0cpY98O05
U6Y90cbWcT3NxNBfv6Ql3DDj7Wb54mS3XpqG5fJS80Uwady22j7UrsLjnfGw9zseTEIHKktueITJ
1oQs7tTi5RpSLOo/mRbi0vtBb1lRT8tbSDiJf2lordz+9f+ij/oGK69W18OJQ/TQIy+OKGly7kc5
wh/DOtgEy8hCJulqW8H60pzm7XfkChd4DqjWcNhgBKl7MCu8aD4xpry3MEe03g4mUSvfCZOPZXnY
07N8QAPRzoxOEJclup/wcLjVBZ6VDyUCma5+y5S+erqBv428gL3Hlx/ltw4Mng6wGgMylNFPA/B5
MFy9JhyYQTjICaEE1ag0ieQQHN0fptTqUvqeaknmsnHK4dg6W6pUgtg6j8MJGq7yD3jScSIWWs54
53+6FEtoFsF26+6VBsJ7RPzfZq+Tbo1upaZXLdQfslhjESuWD/vbZ5YbZalLUyKwDpfO8r6Dqeiu
TM+o/yi0ggkzGo9acTCfE81o8dDM9r67U030nZm3dPZS/3VoPi4S6kZoP4thuIvfF3gOKilY0F7u
ApoTfGL010cms3JLQQWjqdMj8edBWZtKw9VRFC56Me+YRd77zZnF1cLE2YYj5iyGhVT9Lg3qo4z8
N0790af5Xl4cBO4paMBD+c9JsdZq8L8qoz1g2HgkVpLUxvkXVItrf86awzEBRDmAmYOZPUvPtwZD
rnbEss5SUhGl4l8oQKy3Rz+ta3NOIKNqaO0tkdBeaDJJ+9H1xPYP2ccHgUSZjbn2Z5Tw3sPS3YHO
6rOxRJUASIZa3QJ1RCmFyMHdkzxFWGHFr4qEsnUm1tsOmlpsQfRJlHp2qmVFHbKw37ZPHU1i6w0F
1FlceqFXIZRnwEnANlFyBnUocJzbOkrsXf4vvr9ENbwksEKiL6Brz6PnyCoI9onj81k3JzawRRZx
NBoev4UwGq2VQRRJyUFHeNMH4mBC9uwfzC6KEFKlJKFJ/iyPDBowGJTErIvILJ9F4bZTo0iKpVcV
TLHC8l24JgxtJLmdV6wSg9xUFPars7HL9SAqWFk8H6xTD+TYqvGKBUSyLzSHZA9bpOtzN6x4u24z
MtMh+flKzcPbDCmAg8s4NQbgTOuQLCPQ3+ATc3ljxyD7cLkYf6EB+Hb9RtOBOPUhR7iJX90rVhUB
owFc8kzZ41yMK53Nvf5dc7msqxjim7ua0qtaHItxzaMzqEOpyeAOkbFOWMHS8zp/0nIqdKc1eCrv
kKqTCUI4ikAcSijD6Ed8i9xb9gAtiAtZaMwsmwhBSvWwtm21ajmwnxjjapTGdFuFW4tVapHu7Ker
6VLg3wNxjqaxrNMuS8j1bzN+3D4zAIZ+rPd0HbaEDbYURrMVAfVMmQtRwthTxZOnn1BK4uIeu5lK
wvB7+NKxJAp1W59Qf9xIq11EItqhALHVoujPEWkJZ+FAyPs70x4I+YyJblYE233GUfRl8G4c9fCb
GFxfXoynolhiCXIoXITN4n1J6KSAzBAamvSnTcpq/nzl+b1AjJa966JpZMvUbKkDd4J+ks8obNWO
xQSTzqVo9zprPvCKYxIeruwV8GFjCVu5SMkopcsgknJrTlUK0qCeUDp+SH57HIppXDM20Ky3CN8n
7vhs3idpPEGm/ZWa/wWiB6ilCH+LMsDEsQDAJ9MSK8Ckj5M6sCK5btYp3ijAOgzmYOFlulKjfiDg
h4tSHxlr3phRJNz7Y409TvACy7FHbqHl1zdKTDN1msWCqtLtqoNetp1f9y4PM8SZhm85QnX4LfK7
i7v74KSINVm/cdfixgC+M80PDVfQcsNwJP3ll9m7LIbHQ24y0zADbv0hKzt9Z6aTR1XSJ4IiFwhT
iJGUsCilagcdQZt1mcLdJbD4N9L/nS148TUbzxlwRSND7RUvHKmEfcPhRpiMwrSF2nObnqRGEcBb
AyMQkDB9VUWWRM631dub3NBDeJbK/g+4r1p0XVwMr0y5rkdhLwsGIzZOJ6P0K1PuCqJtXHfPvGRM
4JDG7yQ5h3EYbf/MGJZZtasKAm6sNMwqTcC/t5m1rNxutJi9O/1RUI9X9KjMDN3PpkqM5TDWSwVI
GtU3EB+eWu9jhBuU2oyBS89dDeSxEqUq35Qkh8l7YDiKI+Spjyic61Hktu5uXZ1Y+YfJUIzNElA6
EOvVdbsp6VA8Ode0ZakPLuN/fD12eVoa4vMTb8g5XqZD05H23/xaPMMO23wWYd7f/Zvekd4y1Cok
fE/aTjEhZ6Sze0ZnrXUNQ68R5MKVOgEa6TLA3GSPK+RNxkxZG2Fd2xriHJFcJxCHPIBPxqwhii6k
QziU/WZ6xlYT4CY0P8wwkzTien5QVZNkqW4pzfPf0FqRteZzmNdFVvON+/qn1pc3gA/51VJ4Mpaf
NVB+7dVcgs0xBxImQAciUbgI8fzSNqMDLh/4ifKk3/G8KSaiIShCOETilz0AlR1YiC8MmHZ6JDZV
AKs4cPcZNaGvXrtIJGghiMZEczzFMAsjk4oayAl9khbBFe9Rdi/xBFhIAaP34EqyKMJie4cMff+H
VMWxgiTgLuwGyX0SPZ8iwdwIY2bWaqf4qB5ZIPHlDhrjYQS2soA7PJr6zP6tCGFo0gV5Pju6KT8+
LP21lTpDdIpWcdzaPS46B8AN1nibiPTNCqPz/cE4E3QVM1IVF/5orhyR2XC3INbYVMSzCxroJbyk
b21MXBC2bpK6wmRwg5Ms9XveHxIvn8QMTL75Spz+IN3a5hSfHaXfbigrKKsGRgyoxvpff014DisY
b6Ui9RMivy+9sFQPxS0IhpTAnvs0mHGyxXzmYbgZ+1jSqRtHbS91PO/SMxaZY5L8vrERIF+MUTCN
UrzeBaSvVwFk2/1oiSR1yDTvtSEXRDa2da/2wC5Fi59vL5ssfhuFged66/r40T+PxCJjAo1MQPcC
4tXYLiSUASpNu8Tc0NcuZig7MKAkz+miXo/kFxBx/9I+MtyaMUWPDYlX5JUpbk/77cXmVJ7qSRAJ
UBfAdPvoTuBavwYPrM4Dnq948Ku6pkpzYOedokK8D7arf3XggxFjUCNHBx5/o1zAzrGBqzZaNxCo
hv79gOqmG0qIpbxntIJkavTQfXoUJL+AlSYXJLLjJy8xDELOKmg1+d7t+6tDbgM6OExROOz5tlgU
EhhJntjiOCcerih/0JZONzzDENE4Ieko/0k4dDWljCTCAYNO8ZRcCH85MU6wwOzaNOU1vHY5zn/E
CPB7o6b/4z+yZvo3oW/ugMczgozK3gRiN0aAL1FpWLp9gbgP3QtQwGowrs59p2tKXml8WhrFJA/F
z9mG5qSYkU9X80RyuJXhzkMJBj8uTwDOv/QvgLNTGYkJwjZ+Oj7uDxwTOBPpfC/ogSgqBZVJeQUB
osYzwsNztVEUbp997nIzCh83kn7je3u8FEdfp4z2ayLxSzo3icZAzT7C/+7tJF5TFY1xQmrqiLwR
aLMAHxs4hY9Vky9C1GZeQVExZlJC4rb1P0VDlZDy1L9GWGOO+G5SE4PCJiL+I4lbL4eLKlEkMNqp
C9AvbynDkglLHubVa0SScM70+PdE7PpfW+qaaCLVPyjUjLk/5TGdXC8mnbY6AOYZC3snv2NoTrKa
llNi3rij6rLkUT5LiIZ5wNujZfy+XnRrau0YL8PXpf+EbGDJTdaRcD/TLksNxBIzxy72Blk66f/V
F1QyEcpby7ysAJmV8urDzPJOVT2LbbNGs1UWvwN3NiB7zc0IXAP6XiHehozeySRQXVT/XD4jlxH+
HcA0D6cSjS8FBCYsCLK6wgnvw0GP6nIHwviUn0Ukd9QZXQcbn1GEGKPIlcnP/r19xKmBbeAKk/RW
MHc7vIbsTQAprvd2q/l/+HUtG6mvVw8BE57eVc7FPSSV5kA+q2OTrRGQ3Vdx4QGC/v8YlujwYSIg
URAcruP9QEHTyEkHcIEPKRpey9o7y5e66MHIzmpNAlPT83eJn4rt0cRiSYsmAYGcKFK+Ufl41cK4
R1lhLORXsnHnrChgIuuIMcOQ+EZWEHqmDudqgCXM14r7wyybHSeeyM9AYg8Jj3tzXcIIZ33xgJGS
QrlxFDjXukziTby9GSyNGTZJbdkpHi2ecwvJBetKZngizasxFoSfigbrrxLGsIBzbKTObsw3W+e8
ZdkCNQOGr3w+jY8YHyPDI16vgL0+e1rBC6lKYFL5VKAelBGLJj3POYJE/MbrYO/tN33uu3AGER40
9QYJu54MEI3Hfv1mnzAXLZwkq/rY9St1mHnjLIL1jnC/f3ZuWd9iZ+zeWbDoZeT2v2PPEz25unHj
pYMXnuRWautcDd4CT4cYAXcwqwTWrcvo+Wh8KnVLI6YVUHzJOuNXvTVKsUeVTa7RbDtfLUHwpUF1
Zsyfpo1qK8MmJR2s7Dr/W8g+VJSMx8XWufqL/f5qma7ZrqagEdFSryG0bxg81t/lClNQwtZtnvzb
Z1a5RFE4OAuLI/Hw5WHy8DeEfEHWPe+A40PQwtFSSdk3NZ/Rp7Xvp18PrKlpOx+3P3buWM81JEPW
qNAApcvnCyTZYVcfGrCo1kyQq8B2MR5KI15+3AI6yjERS5GXgR67HyHZxYcCIUxCxte+hg/1+59a
82b5lDfLL0Udr4K64bM57KrjyOpd0nLB+nAVHJYOI+5Nqxs5mJykBAF+/6pouYGUaZ/RLaj94MOE
hX/n1cVPHU3yPnLGr/L7kqe2uln47wSlL+XPKsq6n5e/miElwYxVh07C9ZiDxhiSBGPisMKri9Dp
xLVfiAA4BUIVk7l2F7nP0nT8CTuypxqxswbYWBkOMwfp7HS2ZRToGfNW7D6KMSuN1tUVSby1AnBZ
xy+eIu1YFCBhnRWaea6xHnzhpyDA3nD9Vr8AILJ5LVXfBPlCr86l6HajPwKE4R1QyNHMZUisqi9Y
YxC8eOR2NebHZFb7+XgtpVQbgjKlEi2VYd4mHDy590ZwQo9Bd4kirWVkWYToz/EPYs3/Z331jOmD
zZdIBXSRxhoF87f3A+E0R561wx+FHZT8I26FgBx+z4Y4bH6sWsDdEpEw9S4PM/4jNAauiYp+v7Fd
CMvxva/pJDlhmaJ5retGAxFxD6UFtFmuoEAVD3EpfHljQPBld/xAP4FxMNJt1N+gSGf78u25xONZ
Yr8D3MHPVwTFwwceyTZWbQRtjZLFBeglyKBt064/RWKUzWFFSRaDhScUc3lk1K3cbvTYGbEzFlLn
r80ilFftiUp6htajnADAPNeOjDwGCNbC/cjOvf9aRuVDRzJk+SLzsuwVt55vwwhrAvNgglvrF0qj
yQveoTawGAdITN5mUTNSU+pJiErxshpiykTiCZeBVtrXndZBWJo/wc8aJE9UvAuq8FhrEG9HAwcM
T13DlGZ7HzBYBdvTV1tINaoqZKXFsM2oTd+rpmb7TOerPOITMCkziBY2zb9s9h1WsBMD0hTJz7Dv
zoxRbM7f9Uw1cGccBGHrOc6MeYs/pLVIFxMTE/54nYC8w6PRY6WBPDbqtUV5KqgOD8etTBHxm4TL
VTGL/d2lbzqGnnjzq3+USJlxHrjG9jc/vcWIuX0zeIYK4gRlRqRMFrtHPVlqwpHzM2uc5qsLfzRL
DSDZsslVlecePj9bbhh444d3A3ttQLtbZyk3S9dGYdgo9a0LPYgjSjzRXd6my21GebrZUHYQoKPm
OwTnJkyGWC1urbbD9MOevVege9fwnE5zwIkkIQoTco2pwFlALy7qWeKWdoE0tFMvGwwNIfMVRzAn
ma8Ukr0m0g6JQx58Ez8RLUnMc6d+IXxclwFg0iNrPSzUBYf6j/8dfnh9MGHTc6g7RiA3IlN3ARDT
c2JLuoPEF6yN7IERbJaLUU4/jA/S1oOmD2fRpYoP1nEKFgr/cwjbVuyja7n//7hngtLPgU0wGdfN
N2zFujdDwH8oFd0MZydP/qzVUC8qv5VAnzmFj4ABvfBwE8VNStRLoPj9abaxs9aHMPJbiiAqClK0
Hkzwm6QUEidvdaVcwVwPb9QWOjJkQLNLmHGldxSleJU3x2INhWTnG0w79KjvGDOOfqZNDi4K2OVJ
CVWNABNOMHgny6Ap3U7Y4Frlr0OFzgud7JflUG/6wYE3F0n9bfvZ0I1TgEvh2ptxLFsHZ/V+733B
3+YIf7IwxwQ6jSuZdgjQtJdDYIOv7dNCHFZWu8ruZUVrdK8+e2qgMHUbBTgNwrAkXDxXkDr3Cfxg
eihpbi6Q0TyZS7RS+FHvRPZZGEOvEDh0C1EFgCCQ0l5R25v3ly8x5A/OUkYlYSJuWs5mWzFH64Ke
lsCnBumTeGuDeDQI/jLq2gZJRThOZgV6MLTDqYZ9frChpLqnwJ1uu+4e4Chx/KtC4RIiOQqtG6og
QBajmjttMJ4pnnGkrHztZhD/o+cj0Kt6bcQB2NvkkMFwGMdEdLO4TMaZEgWKKi1/9IMFcU6YBOe7
g4H2iv1y+h7zk/Vrzw4qVjBLRoE990+uYm17Wew7lNfoodixSTanNQlFsi5FiPqxFMaU93C0sp29
bc0l7IbiQ5kbIfxiKPiLKPJVkyoX1JVIj2tgsSm5w3/B0XWsfB5VsW2PxKt4yNv0zLAe2OoIfSqp
p31VJLbCuSF+Jk5f/D7Aucu4a4X7i9D6oAKGCkjxrwHiOY7jMsnKhHHz2ZMGbksuju4pguuXkEHv
4Z7bpH8kHkxL2t9vmzKqHN+aPF4ZSq2ubELy9SfXqQwImYaMcdNwgdOOCyroirIKuUXKo4wGPrhV
NpAE/aN2DtwM7UHOQqD+bxBNiR/7QKMTxyZ4VpSy/fefucH550+l5SBZldJMVB+ueTqdiBU82knw
q8t71omd0NJHU/qzVRrdkI9lVYC8anOhJfeCxQLP+rpkssoRaKJNRCoXoI/fZw8kcsKotIGYYz9d
dov/iYAyz7dC7KzTEsWRKxSiiBKjI+D2HErclNJdMO2RW/63FgI7mdHf8NWNtW/wN0fTGdnEjmZ7
R05Zk+b1+du1nSkOH8BKzGK7XdDCtWpSo8osPwIbKxz5d5XcXNghbaDGcncthcviH9+woC8dzRYn
+767C/kurdJ0fLtUSH0kA1ApsIf+DchWAhugMK5nlCW1Uk4YiXpVxgFSMHAFgxZPjKTPmRVmRtcz
cFD8UrJWDScBQgLqdC8wPq7okbtw9bPvpOKVgQipcMnF7yNBozgyRl+vbxl4vFxM1Znjx2Noh4Pk
SgrxDisd2QViEJAYHcGN5h9qaX+AFLEdaOWVl0Tks3hPVVcGJONqe1C5tlOPKv/WbwadFKeFleUU
K0zPyrzdd5AsRVux4T/a9uUEQl0+nhprFyBIIsZwYiW5VPaFsC91ulA/nPHJwFNbQKHZZFSIgBDc
wDD+v6Cf/YfY/zRkrr0Pg5b1Y33WHWwcR79xJJvEZ937PkDpoh5BU+dgQzbFjPXUqgcHapwA7a1I
GD4NHV6nXYw22knb1e0lSAcO5UkxMEGZmVVZEZAK+fdO2yUzniR18T5vWNwiNV7+qq0dxKlfhDT5
G0UencHA79J3TNrgttjegM6lQ873YX1VBIEro1aWVWuyQnhHkoqNjSDp7+iA0Alh4hyK7MFkN4Bk
dDYES9begwiYHzjblVq4WBGPxYVlVdlPMEEaQAszx83qwElR8DbVq4mtB0Y5T6Y7RfXGLLF/3MtE
JAqKFt2SlOY6EjyF1VYyDD0x6xc1eZaUdDoAGnxAmuU/bNaEdZ0+5i5F5IdX1rD29ms+x1FsA9xt
f6ZAB9nvdWLbaJYNRPpFZCVFK0MvD4SpTnAogG66dCWa2Hv4pxY+G2zhccSlmCSuyFeQAn676WGW
RquXsvSZHy5sAT2JE5rkRbyXNtJxGb3i7S1ThFoc52eFEyTDHldgKiJvsLrcxnZ6FQZjWNgPjKoI
9rrXfyHep6wUZlPgS00NPeMD3zvTMIm9KmgXE4sFmKrWgCUkHiVzxjAnGcRP8rpgrHDakra6Ouf/
aasZCLzjCU0WOoQ25UDPSc07pS6Pxy77Upm+HUJa5pFwqzYuerCPZJ54ZkTW54kcNJKSyE8Y9ujm
uGPNfTj9SEfsjZ/M0ZlOxsxMkTcOuv5DaSy6UCI4jKz5mdasJ+SSfNf5PvAda/k0P61i9F5sf4yu
+5wdh6e4drL956jdqdndpKUaj3wtXOposODmfCHVzmB5NwpxO1augVehAIJSZNgSPzkCLJXmfTN3
5FswB2AVdmRKj2wW9lrjGobP3U3ld5Y95geF8mfX0w14JX04M/O1pDC6J9giIuQQRTQNGrXV66bU
qD6Ym99p3iQrIWlFOWL8VRBqzO+1pdFNwa/Hazd7zjUceXMTshM9VQr2Gl7esfLaeXdnPeAonifB
8rSUZC/uZKNyklDaF6a2Gz1PQyHPReK+muv/bEZnhwm73hmZ19+OrvNN1HgpM2c2L1UA6hMi3FOT
nlQ0KTBlhccpyeNglCLYKdvL+4SSw/kBHJfc11ZM1sWwT0ZKjWmhVo2OJybaqfaYGn40ZFd4S69Y
KNCibJU7+fkMtLz8hvmWKEiw+nDpQ5bzXik6Fe8T1hSiPyZumEKDY1fT6zj3rL+vDzHpOSondyba
5L/HjFtPKsMbXn8xAMh0yYmDsRMTQUFwZpsPXrJ5/K9En3LCYIyJMpL98nHoavjPreiWh07TZtf0
1sb/jEJYPLAaxQ+CQqr1V0womImj+39jmBpLArkM0u3z1g4r5nE0I/ObhhIchVJQMcsziUhtQcir
tNb5yoddKprvehol4Hk/HJWdY4glc+uKE2wod/v7D/61vbiiyAxkMFLN9/q14PXja/Z8Vqy1NzIT
GTAXWX2ugzxuN1DhosSFHzy1hWAjNq7MoMzMSZ1K0v4KyGmKS85teGs2izaK2iPx2WIt1CurjWnG
oZ0euksAQPOj3Crr9vfD5h47c8KdbRabrDh0KJm0MrE80rAMOLI1xmh8u9gAbCvwxLoe8PfIJ87r
iDF2UixS/0AwleJfuvAXSkiK5MFOGebZnQb9jOtPKoN/9d+w4eBXB5ZEr5EA47JeHysgfuQtxXA0
rI3I6TYUUDjpWmn4MVV/S2Xa0klHBkGSeUdtm8DZLB5GwltiXD0XHlXHTY3ZSz7JNqpfDJyN8Yok
lOWJeSeTiG4bS0w+dk4c12nu5yoP6LMcHa2aAA9RAoNweGeTmnTAIeIEeTtlcu8Mp1Nnv9SN9aJ8
bYi7NaEX/X0Wvf+r4LZD6Q9wSqa54e5bs8cq2ZP58+mcmVVd3HjEHP5DPXhRMH+aPq7rnwcXJIHB
JqhvmmebpXA1nPsEP4uEbQ9EE4gad84NWGxRSyRUImCtOXlltXvctysVplx46eOTaZF2IM+o6kR2
8gwLFJOTur3TadrZ8hhwm6JAor75AbTSdpw8Miv7mH/L0scmbYJlC93hF+6VT+FB1qv1XLDmoGYw
p1Rusn8c1jvLMIAFuxAvg7slPx8FjHwFFVFZlfziQv9t3WcX+aJUVESXA3PPYrVDW6KvJsa9aZzx
mDFUbXH7IIPf4EEvkjEU3XC3igUDmF8WPCI87I7VBH6g4x4hs9FdMbiYwERkofXo03h0p9q3k+uL
iQWx+7MyLAb4j/nr+tsNXiTMvigt2aL61ZSUfZXa46l9C+gRkho3ha2LXB0kRUHRdqarySbixCp2
DVFXyre9mSomfKLT7FT5plm44tk0HD44FF2c0MLAMLnM7LXWGoj8sV2rjzpQZft9mJ46pUch7cWS
N6IZsB+DKsORLvgOb7cMoYxEe+Rbftdys78DPGjhTyJrjNSb9AU6lOpJvKuVcaeUSfhIPa5wAfoi
I1Xtes/tZ+X9FCQ+gPZaU0aYdd8HJLtvv8u+/vPQhL/UJSaxhoOnGjhjrDvBMeiQjNFZaLevfq8y
a55ODTrdU96CEWOELj7DH/jatA9SO0pj0x6ifcOqfqKGdM+8+qdsxdaKE6X1nP+Abrx+mrXfKX5t
5RNHuitcE4niqAhLFwWT/qt3Hi2U/TpmTnnb/pC6jrCknLAUU69WYjmZgHWF55uBcAeFKwK975H2
JfGC9X1AINKxW51Dm6Xgt9z2g4fSvB0DS+709a1ZOrP5PF4M7KImF1yN0RHy+uKBloywXQJq169D
oUdnLmumbN9Ee4Ru6UuqGkdGNF3rgItb4suN6qFL5fU/Jd070kL2wHaHEbl/TmYqX2OQ7DvXWLE2
5pzS7Dpi/SWPDnyjPt2vpX2Us4Tb07JMPwzNlzQi/8W9odIyqwfmSdxAkMD5IQ245b+5N7YuEw9q
boiJCbI56d8vNASszj+2mNuZz1HpQGg6F90Ovo1kAgOJ2aGjAKV4QrkRvg1bjDL7zoqDbAaDh+7E
1ixDZV3lRuCvetZfDn9DoOzDwdZoMTz3IaydZMJD6Fi4iomxuyKs5eabXCGBE8eoTPDj7P46qRAh
ma6dDEM5rSKdM+zLkP4GEXwF6sVvN5/K7WfCNT2DrHxLc+zATjjcTsNv5cgd79f5dhtmX1RkrO5W
pIlLSdNFE5yNbzzCoGZi40bmmbreDp5OK5k45bssm6NKKf1ZWSrRe/yV4lriYISERQ43noIyqk9r
Kv454hBlwNW33oTp8J5lXnMMYSiEPCPsRSyrec4j+vyUyD2TNis9EHWkLgYj/BOlJKVEvcyWYfZj
pmFWvHg95ayPsrR0fddHArOvjdGk6879b0/r8xLJNx2unrv7wBGAE/dQPZ/EGb7Id5E/GwPDB6Zl
69F+D1RZQOVwB5mxWOErgPL3RLeIojOyhH9BNOngLeqxx5S/enMLO6uYOHdL/UaAh9OOObN5X8Bi
PQQXEvwtKC1mUor+Vp0khdqxriPqXOL0lcJ/1huxSPgcjSP9jjsrENdISBYSFEEfvRSQKt+im3uH
HK/1r7UbaBADP7RW/6ng+pnqidVahOL9syw+H1k6NnQv9hrWD09Tj6e/8z3JYqBu1RkCtR5Me/JH
xzKJh5xRLELxELPDGs7pI9m4qor4qhqxvewzT9DMe5kvYemmpyWkKskr4yRKD317kMvX/L5YrQXY
HzIvLhPr8rXV6VxlWvqxdC81nLbB+d7T94XLXoMOIHnRkTNoMQiJg/dEARwQVgEImZMLFNgMwOtd
yT/bF0BPd6fba5ZLa+tPWtMw6lO8zpo4RIYcJEcugRX84gPqHbYxUWv/WXGAmOJBWsV8lH3wKvEc
g7jwylOwfe0BkfyM0ugNgyEx43WHZba9FxTn91bu6R3Avuj3feTj4lRSxB9Vqidh7kppjjEMoFQA
J7i4ZDr0ze8Ta+YlglBsmDbihWMz8egSWxHXdw4RLYe16nW1JwCuKyH+uMaft47vR+khxnpCuhVb
X6vjC/8UBETWeD+GJuTwxbyDFfKlyOw1q+I16AmNgkKRDS6wV+nPFLyENmDWZnaU7H4bGWE0xsJO
zX81+Gu16uqXDT8aITzkJZfOVf7Qaf09NflQh4i/+wwwp6hq/m23rNj+GRC+b0PBlSCVMgD6MvYK
a7YM7EDbUIsamFqqWeIyn3vpT+mhzuBeLboalBNwfjhM3Sst5L4V5xJua3XJAq2XBqys0DHzrRpA
bx7HOKjdTKHtsQLAG6B07qrOYef0wgOHLwB8K3l5q32+Hm7B+UnOFxzxGqpU9VpUXqlBc9+yJaIj
/pC7/QaKM9O5enQhjPHrJrlKfZhVuK0ir3KX+yuuXwUb6ROWjx9fPtUhsFi2qEnHx+VsJpuvTDrF
PhkcbUbDzE2Q3O0E/HsPkdjebyHXCV0nUYQUidOGnspvMVvlCo2DAqWlYYHr1zwf3wqtuuoGjBiu
Q4etIOjwiEil2srMXM2oqC5mAxUExjZlP9Kc5zK39ZwEbHChKsQy4FTtDDbf07WTs2FaP6xKLxn6
LCZZjz+mLzN2vBq7H3Qu10F2cDvyoL+Azxjq1tq+Jv2LmM4t9q23nBo0LkwqUSxMRoPbL61f1C/W
Atj5EyqpFhno9LPV9vtvJb3wYUTyO/jmffeFPt8+ADC5GMEhp7rn2J4Fg70MHY6d6ZhpHJMD6njd
RDUGLifF6loflZceWJk8ufuIfmpM8eV2Bdzn5a0UhoYj3ouLtXq+Y0dvO+ndke5C7toTbO5ZN7+U
UxFqQccfXJ9uuiOfOWcNfQwlOCAJIf2JJV33lCafptrdIZbPUjeDGZgp/H5WMnAISCQ7mRAkRRAC
fE26brAwqwMOmpDKUdIVOpDxWVIJ4GBvNq4ukhEZOgkZoevwCeyWvzIjCtmV/R8962B7645RX652
H07gINr3/WAvgFnSzcsug7mhQWGlCjaggPGTUyh7M2BYrgp67krN2VCZq4Ar4tbrNT6ODTgQR2OQ
zCeoBBZS9o/Um7JZCB2+/pZ8U5qvlv5KKxpKVad7KqHez3AOok5hUclfXhC5XVu+SsWSTY8OE7o8
N7Ap+uapsLb4hCKyFAzIUlmHhMaZYewJiuAopx5PFQMB4GJqAlPhVNwsvaGYtxpuwoiwmdEdxB1l
o0izkD/rl5FDvC36cFFPcZvThVSw48gXSQMCqB7c+00MPBtOykmqqcXkKXJ2nI5mBxgfdYcrVJqg
XzEdk35bvuLyUCrbLKqL5vEhfcq844ex63kJb7X7qSbU1BNMybPAT1kqlcYtbCFWjtkIf6C8U98s
U4BlHflY11J6r3LlYrSmPu7k2ox38T7f7AXDgevTi0SMOKPsahKzyfAS4+kYJCkgUCfZDdUUwvSJ
TPet9+ajWgRDgOasPg5Tj/qjtjHOwVnbK301E7NtR/e1pNaBTfkTeibcjYXt7n/3Ncz+hv0QCKmi
ievhZFqS4NUXnM853Olxn5KhjJxEc4fL0LagQzzqdGAqr/wAHkEJ4BlIbNt6gnu111AsoGAsjGS4
d5eptQdiuFD+azXc8a24S47qgaGfb23qTsG8pWTyASah949ofpJPkHkDNmvxvCGTqxQI3xredX6+
wEle8opGi8wWn8M4KM7cd9zKI0XQmfxH92h48ohXpLaEw4W5LSvGuLkPTlZhbfoy/MX0zKxtqxDB
SC1lKa2x0mKGSY5LRGrak0KVbnxtKCURY8f0/NjinrpsEQEDUu+iCovEptqNnr8yEfwX9YmnjybP
cLBJw8k5RlvZp7PyYAekrzcNHllufXgrs/kXW+h5Tjvf5/lKfGzy7UMwpR3rSPSZW1U1AISXUbMh
kuAgv3M9BzXvkXq09fVCaDqbh4tJWG0FG0dSnITFnOkEDnvbN4yyE2NEzTWW4IfpxJzNvxQ8aUfW
WYZOkKWpuTUx/qtnD4QvltP/dtntvZff21sy/VrPrZNEfW59CyStJa7xPnAK33LNeFLkZnjTo4jP
v0RZOxFZLhulZPyvoTesZX0CpjbCM/yrvyom16+OlJtPn3Aut4wRC3Swpl1cejyLaY0pVa6p4RcL
LZP1ikNJHUyr/wAGzS2TAJqyddoLPB8Hb7QS8ZmLGJr0co8RKXP6+E2nn/rYdphWuUxHg4Exc3Sl
7AHxl03CHkP5Blb6Q4A1LVPYd5WyjGGC0B5AqbVqCOT0xsVTsL/+W/BvSvfdBk4NomCyI8wUfJtn
2ENqY9GC0rOjZHwCiuZVfDD7HIKluUrb9VE3FxRmyMNF7Bxsba6Lg852Kfta84H++FNmdK6chMqw
WbDOnX5a2DHYhpOE8dwMkRwEp418O6k0cAvo9WMR41DKKxQKBxp5bRJ72bt7PDYOrEiikd7VtyRX
YpdiTQC+D7kJgHZe8AHVWNf2vtV448u6MQ25hR+7k2C0OT8P+F8qkUqHaA0vtTXTCBF+a5ISPU4W
BRH57itxkuTphiT+bl6UwnWVnElwuPtmRP/iX6iz+y2SUaJ0eTbVZdjrpqNmMw4nOuO8JjPtl4c/
zVlGf1HbWMf4sqJHGQimosEjUt3IcskKmGlGFTuEhXpknrZc9uDAE49xPU+153OaLQqWE52wz1e9
vAEJWHWgz6Fj8IM2f6JiKIzEiRviIkMgJcMiOYri/n1HtUjW3/YbYZT4qvSXtgw73hxMvmBTH5vx
pLEyaRPl+vwHCa5+uOkdHtVP+jUyYdhlKPY/3WTJ6pRmw0jgFRp0O9wJH2M9PJUrJDHddlLBq7Tr
IgkssxNnlyUjKN1lfJalipuwgYCNcUEOaW3GAp5aNiftDkeDnUz8tAOxF5xu0PTC06gEtsTDjro4
E7Flp2olnkJm1gg+m0KrPYZE0YvZkk+yECL/p5+j6qWw7+lNTZOwKrsoncaOEXcnF9ugGCMlKAhp
i+BqdJdwT8d92QgJxlrRj+3bw7R75XYx2RXIung61o3Dj10HTUyrhupDtlvt1D1eeHuyYyMyBT1c
l7E6WMQH9GfxuzEw02Q2d/zGpT+FR9afArWsKp5XEb7hnmoH+NWp7ie6sr6cd2M/DlzBzgOi4agt
NTiXxw2Bjes8ZsgC1LlmLVRS31bIGBK9z5GhY1ChnGHKO6m+QBuLH4wta8e9bBnjG77R7tK0XrfH
C4IzoyKZRFAAyaaQFWlzrA9aIQTfYENvUnm5v0brdVQg/faMooQVBFBiujubyIihFOPXFc4D2nFW
MeljwcDYW1YlN8dUZERINlLQmDFjNk22Vf4V+BcEbpZLxowhOzeKzW0iINbK2IFLicP8ZeN5duz7
oKukDlTrJcX2crtoJn6Q1vmXYltpbyl1WPri5JVkfcHUHKouExLQqb4JVoTHUds3aXnHCvBdrRBi
EFASC3HZKvKmUeYNnlPXealGXr8LRLlNy7JbgRPP2U/xT7f9H7BMTvqA6qsvFO+lP7tx84GPswfp
7l8aI8JfgqZj9GWlL4tNuwr5jlRNQqKOGc9at/IoxB+DcASR+3LdJRJWX5XZHRd+sEj5fiSVkh7l
wKqVBl+NjVBt8DPL5qJvGHgvx3/bK5n8UQRMK1AZ1lQ+qRPiq+xAdLdz8tMmD32ldaDZZ+zOxkfk
nyfb5eBWDrEJ7pQZHneS6NubdBuhCduzdeqvJKNT50ToyQ0eva0VxqTBT0C75u8KhyJwbfvf0ur6
9lWIOqwvcfIlkEHoAq2S91zMCN/zv2XALSSHEBwajYwNJ1pqgOVdqSSD6OFQ1/925S096WzBqQLh
9TdxTZLAYEZ30Tw6Iwo4Cm4JjcdAbVITw3CpHN8/ezzsHPXr3jki/msjZolUTwn77XXmtZ2RK+vp
w7iN3YgVO1GVmRfKVHBsi9DHCDQad3vuw4Z80ZmoJfK08Yq5tqiuzQYuRl0kFthBOGkC4nZTcJZ8
kaOOhQVrfNXpBeD5bpEtJg9kbuJLnVyCO1HI+5YWc0nn5Zkj0177razxKK0u6EMw/SX3z0Bv6w7c
qLgpUBWmhM/Mp2q8QJnrXk5Rv4WUNpAYzDwSO+SXijTZoAFq8QEIpmp+thSdeOMtm7GR6Z047Idc
Xur6kxA7Vjr9oMWVSHwYl1qhj5t9ulwmo5BnqO8nI6CP/z11Gjajuc39faMBdvKK7P9cey7ocH6v
8KjAOIg4UtQS2n5SDl2KDK6AyLWP9bXL8nSx4014fk0Rr3+LgLo0ScakSKu7Ychu2QQ39D8ypIHZ
FQfM6hVOdIGp+TDLyFgaPGQBtQQUUAPbEuRE0ABBTnNOWE1HWwDhNevAcbIYQz8d29e1kw2BdngB
1y2Uy2n4iPJAmj6bmxVEv9lAzJp9+apVW9nNC9RwuQjaRQ2U0LNx+grMl/V+Oek4Vc15XutoFTlW
xkjX17U9vHBOBw0fXwW8gKHz64EuoderylhDpIM3CNi7utJDCcZgS24JymSY/6Es/Gy6G6rN0dQs
amgkpX5qEpcK4u9cV8/MVTJIzYTR3rlL0bQTVCfvhxhtsXWlE8U2/9MdPOjqRyBrmVhCG/qL7Ux+
ViTLJC6NOu+KdSGInPqZRoQ1+zJ8aoGvbeuNBEiD79AT3SXaFPAIDRHjItuPOz8TdAfuHTf5qdbZ
ep90XuB8CX62HK9kNBzITjYGN2W8eI0HEtJGVJkq+Lw8TkaEs46OrnnOIjhQ+1H287LUUSy68gVX
Vhm3CQo3Fs5KP+XpuQMebDPaMm4WuJDjpNLX1WtgZ8JFPof4QpIvJd7TQte9Bl4GrpPIowWaOZ2h
g2uNCSfOczdShFliVzTW2Q7bKxh1hZ3LF8BTqM/DFKYrNS179zpuNeM7w7kZva5ui5IjHK0GwSrz
hErg5GKuw6fUvmDOikIYazphj6wL7aGSeeDQwTsd1kBUpGGuTjU2Fpo2vooeAHyxGFIzTk6ABG00
ei47wgiYb1wtT4VMlpDc4MhEBDTVtlhguvxNUWxo1m6qlz5nbHQb79w/nSZd+wDK4XZR+G76kzip
UF9RgFUijubzW25BBVi0JxF51vyPdRo37IZ5qap8LzGh76bBcu6bZnqc4CtWGsrfcbEXLUM50bKf
B0w7IgSXPyef+mFXHWlL+vXNfx2DrJVYEpw1NFqPv3DXWLRKVTRJQn2+oMPIAUohD4wlshDA8blV
xk/97As+l1Jz6ISy+3BBq/+gwtohDm4cWZGXX2YQqm78iqsJwj2j7yC/HhcjO5OH8iF0tvA3IFjs
ynqJHO8cOamLCHWZwP0I2J8kWMN9Ynijf9d/MI+4yeaLzAmCCC3l/hRkGp49QSvoFmUkmZ7w7Adg
g3mHKF8wEVNtQ/w6f/jnufzN/TMgpK2KZFknpa5EIICfSSfJqMYwWx1O+rymq0tfAijNWxuSaH67
k1pt+dKGTV8xiJIZi9HGMuafy8nS9Puy4DzQPAmJsU0R8YZFniFG9FqmL6tSy/lLNFtDyHSBHiVr
4nAVp+HtpXOyNW36FqkzqKDA4n55jgaLho2K6R33wxjkmwZT1lVrLw6JMDgWbJgdWqDtrsQFxzFQ
vFDxl++Q++IvfKBHbziOOKDL99aSGbNIjmQ5ShYsJcYsTJjz9Uu/xRGmT3GEqGoyWX0qrZvfpKnE
7hOvi5qi77Qkqn2wdrh7Mz133/sRGKptPh8xevCrEEsgfsYjegrmygfbHWbxAWi4uBvLqDxrar7l
Feia/08vsKM75D2A5ZcQqjhPgdvcKP7vgLi0rtaivwQ8GBUN6VHr0AIeOEzi5sSu6u0rw1XBCbAx
5O5hMpjQtkoLe70fD2jo6PsQZnuQ8N18v9JObVEzn7eUj07JNCNQ/k+ZVnqEf7yBXdnAVdmxlxlT
IM3iol0qDxFDH42tqvWKH+w0/X1gw2Gv2D/Tg15PrfdLs2ysOG2jr7Loxj/HgYIeG1UQzel7Fk6C
yaCeh5H4gaNh33MQZr0ZZwjWLgrBdfETfXIUb/UtowyFJ0+9W9HYovRWkqaSCMrCUH2KamFMF00A
z3QWvBZb9k9ysmzHBP2oSCQH3NoWAm+hCxWIijOWbH39rK9K1dWSxHHUKqpvx2dd3Qtzz0Xdzx2S
ion75T+2u6yvvcqIlwsg+3umOKsmGAeJt6kVdPQk3ZU39exb5RLI8TC9dbwcyeCe6cNc+NTn68BM
4vadLgg0R+pwynGIK9IyTR23HU0ezpBXU8a19QfGn1KlPgrQLnRHFICRCtQmWrZUA3Edrs8wyzz+
eH92ghLKL5AI5p1nNDeaf+HU483uQyOnlkS6EHl+x/I5bvkzuKeW/S0MnuMrJKFznhc/GXayptcV
v9QqGgvw9dDSJ8uFsShwe1jBQ7Zmmid6PqVf/ApmZpQQ4IQr8owHLqE/JWsp3mkBTHgCmE2QzN4I
LibT/gf6BY9HJzDST+APIFqTkNvEokViiXWEkSgPFPsltbTjQTSzCkbR8lPtHCjOHVAGA2c/u5GC
CIjRTQ7/199ZnIdVhbRlLWla8kK326ZERRXMP9IRXTihX5v5ErXpm0C7gHnIEZ+FotqutdAuEy1Y
q9pKcSQ8BYFIDi82+XZ+vw8anNqhaozaxFGiFKP67YPsDrPoHaj2aC2fnYDA5ydxgRUH0g7ltJns
gt6SIFhS9TbsizsMWF7oUBpdDWlVbXWQULu9bsIoU1Gg6VPszM6d+hHuyQ9lpze9w6HvIGYIl5Xd
m70PMhY6vn5zPKL7vgASNjAwu07SaZkdp2MitCPZnJpVo+ExW4mRsdtzrrqc5Mq6pMFm4KcLkj6n
9y30A2dhwK8jhHh9TNIda9qM++Y58GdtxZ4LCLLCEIKS4qc/FRIoDUp8Yv4zWy5fyKP5ynMbZyWG
P7VARpV7WqNaU9xSzdzwv12Uqo25yzHokSOiVBpRnOsK07DJ83sdIZjxFBe3zL9XOnU/ORCJJ6xW
VjuUjVMdGPES1xcr9Rb7OlW7NWukQ2HDCrj27LWaaounhAXYPX88wHkHmdwRcb3+P4KTrib0N0Vi
FdYp22li4Yi8gyIiOTmdcCAR+VStbYd+Q+qGgWs3BTbu4hdcW8tKgF+SLx5efMdARpyf5vNW7SyA
qWXUfghBN+h94a79K/zLDwOFFmLyeozMiLwq8kJFPwGlqebPmkK9tTqvE/uH9+lky5VsBKLZnFUR
yZyoF4ltIKn7y3EedOGIaG8FrVjngBcnPPNlbyBfOkJU2bx+xX/MInG92jMJzs/eCOjreT2jgKM3
GfmGafTXaT+V82eX1ZED/ejS+J7IpAUcIPU7uTCGPPVFA86u7g1Ipdfo3kGl88ZIFY7VFKYVS2CC
bCtsHYclx3IBQRSSVe9It42dnNpJ86y6g8TifSevcsq5ui5eQbdf5yXv2QvNLm3nIeJ6UO3ZDmmi
rI0AKspkfdIfQVFIrRB9WfaNNSBb+MuKZKW15GENgBLi8pER8oKJh86BHfv4AgemqldhuidgEsCX
XGry75HpSIZZfSI4BlAOkFNhry+WIJZ8wQX7d6euooSx6axGNjd+QLdej1HywcSfEbFYWNaF/V46
ChpaE1RLt2h7dOOWbj8te61EagMOSnY3SIqzZzox/58UM9MCOV/5Po7sP/tVZ81IcDDPwWaKfxda
6J9onlRcLLYojNkVaX6GrotwL4uY0ERzK5q7OFOqKp6Yvs+FICvzjf50xiQ1EyTW9yih92cLVz0s
mNtrIuW3hF1BBkhPjK/ufqXH8B+P6rq2xB34LIrADsQ2xby12N7o/PfwonA6vQrAobf/8O+lTnHu
CSWOQNMs+eETjs5+iGph6+Nxn/c0qr3S8wLcqUuvdPZAiE8ZdYqFgBOpJWHue/DfNADGEBD5wfL8
MXXImRsnErVrMH1MV6ZiPySOAmoeiadcrmA2VVH0CuQH2Z4WGM8Z3QVrl/7HZF1HRY4y/YAIvP/l
bhYqy9sjvr05chLSbGa3iKYHr42xXvq/2PqYbylL+i0Y7Ch/X6L7AgDXwM6pvwKpWC7jS7WEFDCw
mm9NP7GrhxbGKscM2yCchrjO6ISa4D5MGOBnNiH215mjDbTibYbfkdpgYQc/kXuI0TB4t9y/swwU
ZC5F604hBCq5TJYgjeaUOJm2EYpDioIvvGmPYNNdCZHZ9FqjPthoGS7BsLxoFdo/rpewL0x8792D
52WZU73vK2qLfWkccXTsBpKOALyd1O+TOUmWh7Am1GcOEmNKtbU4Z7BHultWMGKhzQ5cXRRlpCRQ
92eLwhbD+5zse61AKI68S9FOxwFNhmNBSUHuRgCPdc0YO8hgCo7CJu77N7+BcVgB+6/APKYY5SJk
eYR1e3DFxxK29YzWqVVDp5CfA+71aVi0fD9caKbY0Iko57mj1L0a+1JylUv4BjlsLBaK/FtjMkyA
zeB8oV9GsjUG360mL/KgGcbrykEsLTRQjI/m9L+LbZpNYHaCaz4wKR3QwQZeMzCAaSAZSs9HoUfS
P89l7BrNIYwm/XL6O3mKvFdLk6jcUXwIRpsxazc6Vu3+cjpPHurjCv+O/aYwm/oh2bTAi5IqXD1w
vf2I7aEp7yuKKbzL/tyrzvRzuKmLSqR4qdFAHcSlN6TxmQpggvYWbHysYXJliolcD6TDmAjQFQ41
pE343cOYt0u6UqW/3HD9D09xHpgRUxXRnSs24FbdyRw+Nb53+7CChI6Npfr79Md6gWdri3cdCXkX
xmrhVOZbBkAa1c6vqD2PGYCRV4jC9aGVD78qmBNpYGpextU+Y4PzQnb746mR6+pZifa6cjA2Tw/W
K7ZrARuNZY/kPKDyqFN7ySrq8mr/m4Mh4mb7qv4cLqvoFWfLsP3JYf5eND3ukcH196ThVyLUoB4O
FtXCNZStPc+Rm4BL6SUmbq7POiCS05UaQoJE6wHy+Jnbpr27Q/T/I1tWL+eVeKn8XMXMwLKObhs3
AF4WtOyYjzKt8szZ/Dq1oMjj5TvbYAcGgw+bjKu7rJIwBnATgMAZbSd01Zp0V+g850Dkh9Abgdbz
1H8Tj7HaCSUr+b99VJcocPGx53aJ4rIkvLetshV32JVOFbDzRxMF/+qK+20IA4gjDL2xQrfImmJC
mfyeg/zDCoOlhn6+GTk8e/50ehdTmDct1tcheG5mxJM/C3R6864Cu8h2vImrU0E9LFYQ9Cne7lCD
4RUXRYaAvBoeNuY4JV4qc11qYp3FljDKeY6GDvV2DL86opuiqcbmer9VSC8v/Vh0Q9wspzNAaKi3
bKndWwk8SueBklVKRkp2tK395wei0R2/YbxJYcJ9NdbYldMS2xNZFMBeOrk6+PyN5lnMVY8ifkWP
nSxTnwErE56Q+TkDN1vRFJUEpXdCeBZZvZPOjKPDQ9yEtnz8OywgkGqtmYA9rJvA9ZA2SuqtCfx0
yDAbyCXG+71SQ37xOicOMHfouzIwo6io9M+Q/gxnsAZxGQGabiPZedRq4ZexenwR82RdX8B9y36t
IJuqOAUzNo6VXiyYlPutP8ko+M4B89vnOakkPRCTOyjqLz8UySge4OEvT8HGr2tll3LLo/0JZPKR
s5NTFuKKV/tNRCe14/6gLsSNuqtk5Y++n/U3JvK4+J/BeElAAY1SHh/NMNiMMVrPPB7e0cmZRjeZ
s1ZTgyRkyPpQBgKPOocWkm5nnoEIdVGU/s+xXEhL50zpjSTUdQ7cirKjX6kQi8ChIHQALG00/weJ
sdpVowS8spmQoEVeURbrUCMrwkuRoA2butgMaOKcvyafrMQiHe4hjTEu0M4Qpj4dl4FjYeJXaS9T
Z9jJTpi+n8vWdR3hf7s6+EGnJXCLqJMRqB5WpjUV7Q6JDwLsUNrbwyRWqv6yehn0lemZWXw8y0aI
+4eklN0ja3tIyF6sncLe2BHEhWaalRgUSoN+lldPv4pRsQPbLj4XIeeu9K+K9cEnysg5p54Ki+kv
pdVeSg5KO/tFRn9TQnMu8/eMYhJ4iW9HEqWhzAOX0SX9pUXLuMMQh4jIeouHCqq3gESDPO6vF821
Vsp8T8wHkCIQnyXf6+0ImdiY5MuQqDP6tuSFFNjHqKECglKeZ4fsNi3ydWJdnv6L6TegwT4U+r2K
3FF+AzbKGiKpHpZbjQ+A6U46uv2pp+X6VbjGq6qUL+xLSVmj4y8ssjbKpggaBl2pLd/8jX7LHWUB
v891PZJ9zbX8+fOm+4PO9G6J6kzb76LREwbvgPCiSlweL+A7/z1fcqEGt9NkNbsp62XaQD08xcRT
iPOWrjXn7jxjn2lUzbJAnUY/WBVOQVaE+sRgMNPivZNSipHJPN0q02lDAxZ0YTmAOAH7TuQOSHE0
KgBdDyVom8RyvsP9pVHWKxEPZQyf6YtBLg447UWbImWoCtoSCT5Yl18CIlTGKMjoUyN0l5PeoZhB
GfGksZ2SV+BznXK1YIJ3zhpZ1/IdJFX7B/eOHnNLZt7KVNwJLQ98zpnQ9N/v2Yg8BqX8HOi0Zf25
0MfQSYXM6DEFuQXXaeCjJ5UUBLW8l+WIbyTgGKtAWYk43FU8WHIeQWknx87n517J5A80GDLnJl34
wcl8XuSqVfrEqedeiCUSFwh2R5kKurIDtpKvuMsYVg3sdR+2C5h8KlpAGZi+Mb8Ad++cy+itxi4y
cPcrkW24GyU3E3xZB8goAbZNPB6iiQfg26QKHpCzQc8OsjOVNuuJLwA/yD7ZlYBeUC7axtYT0GV7
THzGYanuA6qrTa58gfKHF9vyK7fXHwNVmO0X9Ilx8mNBxL8+Mv6n7EDwKQ1PSo9jLiJiclMQF0xF
dQJ1dRkbo+HXxQ84MfMhKC0PnG1phefxl6d4hv+0i0hWROR9YlWjpCbActySRtiWiN8Gk2luzykR
J96CL4FNxCKzbLutUFIemRWGb24Emr0IyT6CIfzDNAC4ZinnWxFGL5M5wNiNRyDYcKIVTfby1Uqu
FeFqRMfruaL70vmZxE4+4fC1i22GS5KnebxOFLQKn4Wg08RvPXO2hMRcG/iiCJngog1U6hghvsrk
hJqzSpuASbVxTlgM0w/tYyOCtoZ2BUkmnCzmLvXSbQfWgcH4ZAoxGOV5urULlTkpuPupzW2wtGdj
E1h52Tf92KHss9/Q0FegG08qhzHaKRHgbf2RPMSAYSVd/3k7+lOIoN7D0d7blg7M5ewyVVMKK3Q7
gbDs5zOa1eetrMVB/fuexU0TFf5KsOeBsiRx7v94/QuyUxa1NpLd7+sWa8pGEdi11XJ9rV0rhwBn
Ge2xb0HKdSlPApytNobQbNe4SCJdVBeku3i3jQhED5fVQL9f1IyNp7OT79m9i7mtFLQbTvR+8VgE
NxjFOlqTPREpeCgqc5nx2IecnNDSZfFkbrfvcdXxsQyE+KvWhRPOiJw59uxEyHC8o85R3r5W2fbt
uBbUVH/cLel85tQo9eJCsz9vpFyo32efTb+iSvcFJGyej6vvcO84IspDbVAjrTpSGH6qxvgyesWV
DRxtuWQ+UrKDX/9/m6P7m3gA1wuqiOxlV9Eu7cW5L2/mD2jphDKoH6lzgVxNJfedDiQ+CCzPt4sE
RTxxAxQYAGUiQgodF6oYptbsnV7sXUw1QvgcCKP/wbCi8UJLUZlTel1Wcxyc62Fsv66uDdvkBmq1
eIoYfHdPPeDfgqihFON/LCGPYeDlLp2xsgphhHRAoqkomNpg89auLYhxc7n8F4m5k4AZ0nhmvBtM
V9EPrdoqDLYEhFy8/DnZHtGGoT0ykrqT6K9aaLwt8GiuimjEBgeULJJua72avKoYYbPUPVKhMA+J
8x0eareyk/F1yyXk/Y56uoxPi3ff0AJX/sv0LQliWiCn4QNk6icBKYTrBNadUmJL3JEcnx9JqYUq
0l3fFjF5UKNeuOrhJiExE0GvBcTtzlMVjQmzUAbLYpBwhwC1EPBd7X4Tf1EwbmZtPE0FkyF4apDd
caLtHGTIIb5VmBk17BCTwKTnJDmC2CRFNMSvCfQ+f4OOwu+R2Q1Ru0Ubl5suT/HUfMr/T4j7L8qS
Iu8ojPConwyZKZo8qiZYszxqN+Ijt8wCZxMsLcQyZJWFLm39kMW2W4qCBOhXqxSMRPbeB7UN7sKN
hkXJBrO9d2j3pat9WEzJQoKCnGuwubYbyrn+sVKhH17svl9pT9Lprl/qsYBPsbKXy9lHo6Rrbdy5
7puzaEeIRlVEMB+OSJEfBJR5tCCPX0+A52jsTiCBVbms7alBZWbb1rv3dOgrh1GUuOslc8BziNra
M+7s91C+xtKAt0xuBlWPM+s4KWSwLGdsd/xHlqppqbpzk/Q6FAPHaZGg5jfhBBEOt3RMNx99vyA/
tmLIZdzmieAHQDUxO6+0arvhne352OXTm8LdoLU0SU1vNXDhUHT8qJAOqPAT5c8JGxnGUnYEr40N
trgg1Q7Ok3NPRCpJfBzRtFZEM00CVgUMuABQ300O/p8Zr56dtAlQV2rSD58SAESkApWuq46JHxbG
9yZ/HRC9t6qBd2LRW+7brPPaX5N9pxIi6wKdw5XMNjisBP3RpSZyjSxWXTnT5z81BAIkSLUkg31V
vij0ZquWYoNvwDG+Hf3EJqUMhjkZGlDVyr1a1ZUMaoCDFCn5Oj3i0FT+Ce0+mud4CndgaEEJSyVM
M+oHoNrvqVXmrOmaySIj4D5OzpfdEK7HuRu6980d13KDdgTonV6X9tTpXkgTwDHIyEBdl8voQQT4
7uvAGRiGgmH6BzqjFhCFwzhX/x6Q/aBqANuIRr7gJx74Mqq7W1qWTMTqqL4iefwglNFfEHi4/r/t
rFid0TEAlGtcHHwd+wUaWU2wiK3rG8272g7CGtMCcPYpJx36sPZKJdTdX7gMWQ31CCVi3c8bqe1k
LCPG/V+1Gi/iRJWexfALGpwe7L6wGb/00iHd1OzEYYFSaeTg4OslBAQu94QKV0oZP0rV5G5n7R0l
NazIcdIsNzKj2ihpg7cGdGyT3R4unipr1O4184eh3LySzornZYoS0ZpvTKPmYLvRLY6ZTWAgIbky
SGOHk1Vuq4TOiHjBwlMJT3BRn2De1IOJJx6VQ5FdbQ1ZwjYjQwP9rPsUn6jtCXOiL2g+ZVQswIu3
Ic/+LE63HzdxrxobWRWbV9fXMJUywtUvpjhYdbCYtaRWCeomlicevFunr47448TuQc5u37pK8wzV
znZdZpRBCQ5UGL26MrKuIm8rxDuZ+Y3MYIn8YTpczOrGf9T+3GVkS/PASg4RsSZdNbTfji9f9oSn
6tXn3NG00qUfmvPBi/oSosDlHtMutgp0A7xo+hq/mohlPZ/Rn7LDES98cQxRDho56TTM47U4yTIK
jaK1UncOfs6VLMs7fSi3nuvxM9II58AxFWReCTGkyAZVRZ+LOvJqOyAuQO4bHR82mZ4rfIC0D3XR
OcfHPYLQM+MltVCbJoozqkAEEX5BrOxmQbBZMPIISJE8ZBDZ5Gqa91oS1evvtmBNXjyilGgHkzlW
+w42wKMRIKdip/Iu6+x5TZJwcIX28Q60ta5tLI27uungmmuOs8H0jBWEaRnhYJZEafC1Pd6BrNXc
M8dy1TdhBz7DOhutX0fWkEKqwtCk1OgmWtS0UZXXC+e96ctTK1TLp+vAUtv4sB91vTxe1UJvwDQC
W1bAkIcmSpCx80ScGXJ+Qf1DLmWk38W8hkf7e1UuWGkHbtyGEMnjhTUdP9bc77WlK5o0nUvDcbjp
1KBoJictN/aYcpWFRgZ0Chk4OuiU6xYbOHVgGHzekeIbAKP3vmmHEGEpbRKZFEK7x9YqJZ+caCW0
/ALOO/PmZXFHskZuB1EN67nyMacNQMbV4IqKx8ivopG0kKzbGDvRI06Dd4aEceJmyuTsXQNZemW/
7EoqLkLN4EdMpns3gB3eoSu6k+JpqGqDgSdyt+J5PtHIJVNTtw7wzwEsFTodA8YIjBy+OMSZWPGG
XZd1l8xzV2LoNLybs5IEFBA2V2jXw2G/IWmt9Nc8puLEm+06yBJCcvQp7SYFYfa55AOc/pihYkZh
t4WeVc8AIobC1+L3/D/w4EsDfeYW/j1C430Wk9++RZwGHCysoOrC069kKChG2a38R68jbZ8uv2rh
8whX4fbQWQKg+derngbiauuTvdqLHopolqGdHn5rM+hqpOwE8zC96gzTe2zyyt8eMLrK2Wj2Uxmr
58KXa3uBTx4kyvhJ9jRQc2mUPl6W1c7fYqJY2ty80fwOpAeiozcmPpqvudvhPuciv21bgUbT7oZ1
409urHumehsj9QDddVCPIjVht0kd8OECVeCKLdPkTbnEgV2pGgdUZ55R6V9IUiowt19NWIWnozY9
vEkGKV0XCoaivAF7eSIOu/c566vfniO7iXedBKugJB+skrsb4ShIQxzx5Vg8WFVDpmbSsw20zSCo
f5qUkg45PUnZgoC7vb5AkBaxs7wnSKtoyekQep6UmCXll+7wc7bmTbBF3bckKlQXyMkDXe8AhQK2
xu/w9KUjjqMZHU6hKnxmFVcjOOk3xwRxUoPNy3sYH6N2ppM8/wyC8JOA52GjTLJ3JDoq6tJ9KYI4
mdV+LdCXwMTIUVaQuHvvprz/CnMN1s54UonAvzeIWYoqwOi2I+MqVDP2+jzyajeb1oJmS74XuZPP
zPKcZqfUYDpvIljBUjcv/TSU6YBWRni1RBKucC8JRJgjE2AN010N+tqZjEHND+N8x5cZx3O9Rp8a
EAM0FvIeSFmv4MOGnfsbFjWAF7NE7yOqH5xuCztAczJ3k/S3vr7TGsIpbIJLyxw3i42zSg+3Y/u/
7S2RiaGfuFU6XO4h3/116uEtyEr2/GAWl/VGdt+juPZM6BcsczLo4l8etaB8zS+PmUrZprwenzF0
oMuzrbj78DsLl63mtIuHnUWljMm4OXeRxLI+WZk4/qZKkmudvaIopqiJp7ylSvVKILY6y8YPzsKf
abZORtsLUbvIB6AowsoxVZhqH+Y0QeP9GNqhVUiR9MfDG4KAMmfp9pCrWbDBb+Li+4Mt0XmjYK2s
QulR7rNWICj9zB4lqI2tdFaboctU7xcY2oV/s9AwsQn2jUlk77/gZWud+UAZUUlZU2apiBYg8pbM
xHE5DkgXmIrSdWmhj7dlD1DtqvwHJCg7UlYWxzhv6H7sy0ckBQ8dQhiKiPlIt4e+mAqAlrl4Pkx/
oS1g0uy9E7NyOsMLJpsjMsBNaBpV7YykWTVArj26P23JZRpwWPvreMiwr1vc01jGjdxiDFrwxGkh
zR5ebEk/H6RoEj4OchP41d26Gwj2bK7MBln/KM4iypTmaHBLZo3qEOIEMSjO2aeAGitJuwZAP4Hr
mgsgTOF0Gs6IBSgsOWAXKyy0C7GI4xNJsz4LgCL8tUPM0TRn/Tr2Zry75TA/w3knuaT/kzl7tUJQ
UpNuZgbd91QkXsHwxoW0sxif6zntgwpzCWeXxO/fzK8OkxifX7qA7tcpDglKSYH87B2+377QjdR4
RSsoQrTztsFWXGzo3/x6Sq2wkvcvpFmXcWJ3VmeHt9sQQmjbirNMScTmc+a2kDJ/ISR60H0IGNWj
cDaR8kmjDhaayrWUWugUBN4gdiU6VeYgOv0VtuZoWJhakjqXdWy+ibVyxEmcyHTWcO46qyU8u6qA
DojJMX49uop3cFZZWKL9+rS7nQ5bkycsmQ/l2VirNpIFWcWuXl/f3+GXvullkBPIJwweni/rGBeb
XRZCwNoQW8ds5wu9t9wyxpzjqVAsV6zZDif42LhqjjhlkAYV4ezqbtB44P43QzXuciyZYPWauRYW
OtE+goS9mJx53qjyJtiFLaGMUpitPrWxBLcoPvXugBtbhELy/UlrquD2Tw2a2edLlu19lvvsaohq
saX+24u5al2BEDd//FRF0eOT4ybWmHOnmwjz0Tp6XmfePwbgeLx88V8joguWczbc6mTj+p9QbHWu
aNGKGEfPBZwlWzXCju2AqvYoea4EUUjPBBWX8l6JEqRZJ/7K3jV59xSDnkCg6ydCKYeP/f6nsyKy
5DJ02zXfKxzfeX9L68lfUg3FBsCLCzWpdl8aKvOyufcmHdtJXOe9VAzR9ZQYOmMF1miUjTLTDtPP
p99Dxj5NSVnTgo2Jrgs+i7xW4SIqxNS0ah3IfASMWyvyWq7oXpZBLaUS63K2A5KUa04M+NwhYBRO
Vx8PnzcB5KvuL9Fduc3Lh8vQmKX6/cW9PO67LDQ0zPQDvocfOAOFT9FGfAMMj7jbnF2OnrtuhOVB
+sdLWjnSO4f9CRJz0aY7GPgmAlsRHmxXRxkg4UK4feRQW3MVCJ7XhyfUagzUKTejqNqjELBnlipV
6m91AaQLEKPGalk3pMc1Ilu3AM5YMmjeWzf8KcLktAZ4Agg4yLYF1QhEL1Eqtt++NCM4AxNknLua
zOZ4QPfeo0jBW/VDNAA4gl0i/wTgWT9IByLSya0h5hdSAofEFy5ug6NYF9bH0widz8sCkp6S2b0v
54PBlka6LQZ+nvr7jLV5Sq4AiBQFGT29HOS179tN9RxdRne/qzJn+mkdHeSSFh46HqUlvVrKrzWu
J8ycIdi07xDi67fFbbKwEwIMjW4epnji+Ev/fpYsRHnYkLFYaouye1m59h8jnpJswGzASj0kUH5r
jMfUcSdnHD4HFW8FUD7SeP0xY1mmzcHd28E6EcHUOOGMcLbx3bLOX+aP1HVyuAp91IlH3yo5OYWo
ZvzO3rsF2AFUf6NcCC8f2FWX7yI4KlnLgp8b0tOOIb//TdXK5Zdi0Hwq1llY/8rkkfNtIFulMGDz
Frue+uvvMR7wTx5jNB2Hq1qeJn5TR6rQyBxBlPrHgZgaLqEwP+XJH+SxwgFX2aPzZclOzzN1NRli
LZ6y1zeqQgb2bezyXd5+WhxGpa8mVnZfO+U5hZ1vcHeydzwn0bpixR5TtsLfsh1A9OKji8QR6ZVI
VUnPKEM8Js3Ud3M45Ie2sOPyDarp07xYo02L9aRzFwK/MPQwIPR4SDBDV/31793W4F1eXMJLO2qb
G3cxIOwwZ13tjxXUpu8QplYlKiC9Sl1wAis40xIiW+LBiYHmWLAKBZVs1PpCWd5YFl04pCL7ftJF
+U8dOQwgyen9rwzQstIq9CnkHieSUhyZSUEPayJeFhzmdvswqVxdEpk2WWfj20cJHWJyTlTvtY65
fridyaf/NL2kcXjOB06RE/rdzIFj7uBL1o7GOuAEbVTYe+KMnLT80V+YvtbSwEy54dpqemLbV+Cd
iYVGtW0RwWHqIVj2Mz//33sQB5vGDEwCCv7751SLyhFBvtpnFJVKMHHI+bo2uJvi7f4cGqAv+040
iONqyily0sVKYW8uSX/PxKN8EvD9TlPaxh7B7n+nuCsK9JhJ0uCCBhjyuj5u14XARklroCb7PcTE
jP9w05Tfe9aEAHdOowLHEjLi4BVxmSP/rb1888bIF5CKzeF30ZXWuYmlLCJy/qSyXtiMvCovRI12
E22TSjKs8q9EJ5sbxELHTjSioMo59lXeAWEsfYXbLHINveqdkNFLp2GXIA+xowNsVzYf22xffmbY
zO6Ctdt+ASyQX1uZKOnb3enRYByN3cJyVkBnPG5vhaAWVdID7cbwvm5Qnnn5NY6dOt4n6MA5fKTT
5Y4xKcw4smyoyGpLpki89MqRDb5HVY92LQlKR9E8vdc+c0/ztaIo4TURkDdQJFGpGu/psEnMSsZ2
zNJ5qoDp1QcCI853kE83Q0XC4gLiUsxXNXCw0buUjF/JQ8tXjZuuADx0IRscdiY4vm3WP23d2xHa
Ms23rTTbOYnSK4psY3I4LYln6+EnZE9UeWfs4SGQwJp5hxaSi+/KPEfk3fSO6hESaKZN0WklLxa/
Vy4nmP1r6+M+6ilZLAR3WRhh+RnF8l9+ZSxx8l2Q8BupDsExPDUZp1S71FUKR1okICGR1iMv668c
IhaTk5lIuNr7cR6w1R7rgzwge6zNPzthjb2dUZKwcHlq9o5kKl82ITOtVwiga6pUWG3qOKDblZby
SrAtnVmygDr8rBqoCraWLoD7e2IwZcOgT529FuAyXrvgP699Lj+1OSy6qoZMroYrgG2rg+s/Gs/A
ryAqpNPP2Oh7s3VgVIHnT4mxSv3lb3oFZtcGvd2w/Q4Uxgt/dbZEIj6Oe2cZQqsM5uh3pE++IaNw
yjJbPaylj4Yh2pzA9rXmMpo+CHR4Tqzwctyh0jQWVXnQmZc2DbDE2lTtoB0BJguALRTG0RVwPJyS
SaKLEJH8OGDUoi6HLZFgxMzomMkjePPWNV68Xb9sVqRv09JI7WsTTR2Ham9MEIel+3BSNMUZTVKj
NrHObTeeiDFgKAAYLzTawqTBT8ASbnT+O4VNnVd8v5TRYt89A12MDsrKQRKzheQFR6hBRHlMlnmG
ku+09kA8ra6eekW6y3eFDfkFMorqd4BWmtfsfGQeZqXbW+lbePSdBUDYuGHgCi/cC3suluWePPD0
B2JNhpvPN+MqYD+ZxA9y/Z8vnbYkJCV5XPbyg2t+c+wok07KnXLOzI00EP7tFh82D4dAdF+LLdKF
zTGn6eckDLzpu6StclQBDOCQbD9bTMBJfWfLcQYjkUcK0otNM+NbenzaNQoAfzRcL5DW1/CE1Ood
BRkTxdAYMV2XTPBCI7gDERSBLP8eMjSpVoJtxnyKOR8RAAVPqPZH5jh/FzInpo4BTXXrdiN8AiYr
F4/dOF5nxMCytm4zSTpQuDwBz0p2fC8y4qa0fBFRur0UtIRSHAazMaFndtSYb7cGz532fW1it715
P7kBdMuF+3Lc8eTIyPIohhO4SwQ/5BzG/bBKnFblQO/uxhO/DIWMrQdbzL6tApRLq1qb3RFFPrcP
Sv3UGq8VKorZcO0WIATVnGcbfM1HBTG8UUNAf/hYV1LXi1DS7VSDQmUB5AxN/PH1gxVBgohXi6cm
xYbeLXCPb4E/JqFCyUi+LL+4/2RbZXQ9hytohnVbaq/c71mW9SPTqeB+2vdfFsRtvwT88+YmA9SC
KegrVzjEmDotJ+jVywImK/DN8F3VwLK4NB8pYOVgSk5b/NAGWHtf2w/bmBwJzjfYs3WOv+iWA2Cn
PKCnw1vwZYN1zix18HFZ1kDoFwFeju13OGDB7t0pv+1nidUhnmgJ+BQrKSRMLgSmYRHIxUXgTFO4
VmGRNdJSHeb7sXYiyuHW/YinbqACdENSOk2NiujEsezWZVTMA+uras/vI4GWog/uR2aNs7Ij4NKH
ziWaqN/+NG204iEZYIyjfuYC0jVkEzJJPvtRIfkoxf8ieweRS17hrWQ7TJPwf6pUhai5Qd0IaFBp
6NECBc3w4Wg9+MMgViP61mIrbCbXtZCvSyCQxzT420zj6IiWcGmxbvtFZ9iJlwyTCcVPvX5wqd8V
q7sByBXq4ua15KPHmqmK4rCdpcIxgfpxAO/cn52YQCdBdUTj2FwZVKnapMEl2Fum9HUk3RSbCdNx
GrCVkpNWwsgRtQo0LOkBCb1Ik4FaGMIgxA56ROXy41YahqVjq5ztMxHagFHhlG+EdiELJ03heEET
Gp6gqAhj2KhpPS0jpXYBdQZBSaFF9EJlxcWNaWe2aOIP5AaTe4fCtSBnFfuc3WaAw7IfM+f0nyg1
NzLJEctr/IYAYxQip6HzE/OIqGqLeyn9TstXZP17WBcCMPQvdxW9tKj72Spb0rpKVeU/9oaCsRqo
+tZAh3mKIEO8fseqU54sA14hEvhiqR8ILCCsOyJsLH52QmOTS84T8F1ryeJI9jQw57mwaLSEix06
BrQT51B+iY1QAfNdPdzuAnZy4FXuIDYeHt8eX5kFsDWzNBAtb91ld9JslBiPm5Yju0gMuZxZOLt3
nIhYP88dqi0bzjGjkFSEB2TY4cwEWZjRwzxxGQhCe5xZJ9tbTLh6EU18pOTCdlROje/Sn+YHbDJf
inF0MOISRJ0CmpDbp6ugX1H9f9tljLE70Ua9kK3bQDWuv/aQJg3H8T/U2PSBPwnHsRJsefKSNBON
nuaCp8eL+VqCezE0AZoCckmeITXe173mKRsX6Hfj3eo4e9A96Kce2FQupokalW8vOV43jeXgFD21
F3LgsC7Ba1HL/yPHxzUmQQA2aLZy3QhZBJN6GK4jNuIaClNWYR6k11FEMdAMoamV18b2M45PWXaN
cVbmkrxJMZ1k8XYHneVHsXo/naCl8vs0FHXNmqp5R2dU1Qrp1nJ6QxvKBt5NCtwWkCyHR0mz/PoN
IYHgdE5qNEahIFmEA1QmXsgSyNtIfWT+v9jBlMJL8Mjp+hQsJDrFdKwrmKB9wnvZ4u2v6ZYwUlvm
NqjOtQImeGulizjuQLBZ0WMYiqUGUKvnCnr79UNCdmtrBVWWrSKmnlTz+VXbhFwN5UekYOBFHjaj
+bTzkOclxAQwychVzqFwJk/mUDtjKBpV8AYV1VzrTCR1/HCwiXqn3/Wxr+12ULvTYfI9WVDVqZkh
L5optyRDtvyOU7UT/Dker65ZfXsBj1BwdYbwvOSweChzke10c52M6vQXKMjY49A7/FtUQ2X3lrQC
NVHagpgjYdTx8MdSXHrpkb5goYMgiHRFUte445QLEdx9y6Zm9RTtRtu97bdpJqrXMiRD2R9d2NVj
Kd9j3yh+J1BbV5VlP9XXwn/LBZ/MLVEnuigmHn+/LHhzu88H/ApML7P9q81TtH6slpT/Co+fwzlB
LL1E2KIeRm5jZcYd9mq2g8ZvGbp93SIig0gM8FmyTMlQ3cvw6cZ9VcmbJ4PPenpOVxIJc0arALRu
mz6GFvYBb92g7TptlTTLIPuWuCPAke/tfjQn/yX2W1JPaIXW9Zuk1qt1HzdjZ/W9Q+58/su86lvW
jZd0TPz1eCtXYHW8J9KwtoDJGvKStQwE59S8ra/nRNBk93757jwUdzLO7c2S2tGWwwL9VDDwujcl
PkAqaOpfcysSu0CXqPLa3407AHjGemnQz7Qj1jhYttC9jR9utVW4BW1yjKp8ddBk/d8sskpw7/N0
B1ZqrJKPQ8ekIHcJulpTiHoc+gUCFZZCnxKTMPISiNv6drb5+rXk+NGYgcBNSrhRAEf2HYpGU/Fm
S4ngyAsZ5sz9M/EolivCuQA08PMVDFyZb2l2yS5X7jYL1TZd45+HrwYrOA8rai9ycBXfKvNYmjFR
2WQrwNcYUh7jj6jJiecges773iETmOluY72a3wiiOW05uVYcgPZDnPXtSZ06P+DwvybeZ9mXd5r7
is3cuiTRwrG9UasiRKO/OeRORC9Teo+RAKt0eyaYUUXGJeGE9U3qE2nxAPWggEL+5CvaVY4r3smw
3rpN6t2bnWI3Hlh+uKiZQiXkfZ5uJUz2Tm374BSbVAGQquTtuwbVmmoeKIDLwmzYu8/kScZ0kSNo
NxVmjbXyROAUCcifZr2m2VV6i9Ao/P4QFlrFC8feMbtOSfzBxxG6vTtS2rD5ED+ZS/nwV+sDzC3S
iu7isv7ff9zuRAqtzH9PpetOd8oD2KUQBqMSUlnK/Smed4oLqMyD1iSVtpTN2MTznQY16gMriQ/r
E+lw4LG7/5tZCc9tM+y1ltuqlPlnGMdRF3jJN2RqySiZyI+RLv2TzNdG31FMsRudmrzhghOpJPRA
tZRQLrTLHSXw5NFlwBPoP1t1ORQiuBIOWlpv90if8VfVX2P0lReh5ESvzwPyIXh7oxNe/yfeMIEf
okCL6L4Kr7DWt5+PZWmYEGcXUK81zCxuWcOtcXntYNMYr0UBg6W5tH0M9esP/XHKSmYqPcD4SVdl
r4C3ruIOju649VXCXSMZEWvbEsT0jiWGfAdlzaf9Y63MB2Q0hbd+LMHOyhhFHEm7vRzzCpYp+bnA
6YfPCtUzZ4GaObhSSGXgRsxOiUGjy5L+v+AHVCZ7cYh9hxMWeCHOcAK1SHQ6o5NzlMgAY3+3D4AX
f/YunW/WpGvUhwBQvFlkKLgO23EEJ5nMo786+a/EbwbfQgBXGZY3oLeNmeQuH4j2QH4goAHDmmfC
muMJSpJ3+yYcWrJTi8O+SHH4phY7ToOdhw08CLiTKs+t8QsEXJyUhg7GcFA1fzC3s0JuvDqY+mqd
l8t8KDuCpoQk88uvCqUZyIdPuHOLMzw0sHjLDs3t6A/Z2D+EiH9CdB5mz2DYQ0R+8jKDsyFsauMH
n+X3mgZFfyYYG4Z2QNy/EZjbsxPZ+UdI9dw71XWJNDMn+QeRtPLWuXmmYH7a0hyQUq8nMdTcGkz0
qnV2tMbulaoXRP+gaw04xea5tiiYsvxwFy5laNxODs2fD+HwIcuhij9lfRSTSx/LYPUe54EP4xmu
+LjbnPtND5R5t/LSodg7s7o/BRvEGbxGk9h7QUny+uV7Wnv3qhtWqeDXaP6kEMStMkSL6Bow5UFw
e0hGniItVZ+LmEds4q4BUEPR7nex6xgj0lIbHymxgtr+nB0Nie8XoKtrhD75cPFoM06s3d5rnCyQ
cD71wnOENEFGlTIOZl78wXACk+rtAcqiNNCr8qfMU3FXXwoyHTdo9WtxCJEVMX6k2iw/z6XEir+4
16PeyGRYfIZgSvb8tIAkOKlEyoZxpaaOFnoAXvwttcNdLC2lD4gldcuNESkUdkwEEWePjbnz0Xku
tryjHK/L8NAVA32uQiNMXUIs7AAREsAwxecGZxN3XDI1Ecx+Ck6nj3kHASevCVnbIA6hgGMkFSQd
E20WaB5Y7QiGK5HgJsKK/ei71JseP3QusDw1WhuQpuaXN5DzOQHwOc7QJ4EKDI2G78GmNbIchFWB
6lCK+0ZvvcSPcbzXCMOW6nSVVrKAYtapvNDsl7O1WaM+SYgPGqqnN8/0M/FDufzq+DM3/6SVZ39u
lWO/vtUrbPPWv5IEW3ZFQQ2OlaDYC/M+ziZOlctwwaq3T8krXTfeGniYEYpooSZ6VBzwrtBO7BBn
AkjxvhOBRFNwXVHUAxqJcl7/xsW3XaniOXM/sV5R8nuzCFh6LbGw9TH9UwCdlzngrX0NRZmKfCGU
iCe4br4oz8e7xRMcT5gLvMK67bNe4cs9cFZLw3cDau3mZiwHY6Owkpj4+twExpzRxBLrQVQWAooS
vGVj6csUl8mQzhwz68S1zsH3YYcGazqXff3b7u1xq3JezJDdmComF0gVGMlTTsLRQwBe48LMVXgG
sJu5OnElSQSi7UGxhi9VJS9mp2JobT8kDDmpJRwqmf7clYKnYKiUzyo9ZruhkJiraTEM9q3SME2H
RlTwDL6nyL/1x1J6ASxi+SWduHk/tlFaEDt2HKmZGRqNUOem22vldRynBY7Dn0K4Gc+Eiw0bAqrW
JDwmo16Z21pNzeVOINMiepbUaVBsItRPmZw5Y4m6bOf3A512OBn79UzC7w5JCHtgy2B1otePV+yG
J4uwFiVR1ueuA9x5+dpQhHh/jGD1jtzYabGeF5XtJc74jYxg2OEW2lCuiT+c7h5P8bSY308pLlm4
dykcaN8qc0+6kc1dNtwyr2astiYIc0rKKixC8zJLvgzEV6JIv9lygLhQcFPzVMxpYd8KSriOBHal
KzthSEscie40Dry+6cnDI29JPU3U2uABGSgnj1HsGs9i2suNMfgBIAUjybAi0O+oTOoi+nLFJ8wK
LUeachuWvpJyOmccPlL5mDY8NfxtDjyxg8Q7BrZsWX7xrMFWiCps5KUm12hE4CFYuC6mr6qjkWk9
Qib+mHFFvUCo/+nDys72AM3PzyeBMLyOBGiT/sp7yLIUhSAr1gxfMDhOussijXAWrGWJLN4179rR
+lpVEd9pcKvrb1hqPwXZliXOjkvsjI2D1k/odqp0NpQy70yZ78gnaezYSZetFX0wF4fa7tH5Rqci
MaPJqFeLkw6nxw3YDP2p62eL+/uLtmtXTFPQcXs2PZwQyno55TAQyWsxtaM16LRjI77McqjXkcTp
acXmg9w8VIwWLGrG4asRR4q7F5UMFNdP6++heQTJi1M8lGlkhw9/dOIynAK3obr038tIs0U0Wmt7
apx8+T/GHbfh2LqBC/8rXbIBrVHiBaBsGjaWbIZwV2h4HCJ552EbL2ckvUz3QXf652LEeuxEiDcf
VJ8y1luLXyU+May+FQVZBh8yjCEjMSt2mo8+jdFnbQ02HoA9J/NmJCbejNWA4fNdTKCeckQrXP7X
RMjGeZlTZaCVanH51vTDrfq8iqry87BIOiuIuiqfencKxfScqfVINveVQO4kOoVvxpnBZyQlNxCX
/xNhjSzrtFpBFe1abqNXe3eTUs9FBAPvMCclzl8tgTY2/yUfzBVEASTcHsCPt0rHYVIUaNG2YiLh
Ts6TpO1H+T0KgUVw7diO/C29t4H36jTI8lFT3F4umoO50RF+bBSESAGR3d7YwbbxZibmdHL5hr+M
Q3ACJkabq8C70nS7yEOM3iRkV1ohsm8xBgnQENGW5mtJYTqaOYFR5swmkr4Fi6VIXoYnf6m9Hep7
HNqWo+N4XUNNJTcOzSRJiA5h0LsXya+mYgE6p/ZGV87PpsJgIrjomb8D+8JbV80lw2OlalFVmLg0
B/8XH1MOW5cnvVJlRTZv9HVKvV1WrQqJ6pmGg+4dbedBledkGaHGXSdVF/xYW/nRazy6PJccFSS3
kZTNSP7pGKfX/GkBdxh8Vz80UE6582wfDikRhJiU38Jg6afsleP/LOUWtb/5vm+PbTtm1wOlIXEz
GZWvsg9aRGaFFqqiyynM4JkCwobjrLsIJTSt/PQpLA+Oe4XH6Ht3kntJr1VBdrktgsXVyIT2S5AN
P0Uv77HrLdpPUgzCEA3+o1ULax+NQo7T1Togl0I/cAE5lKxrpJk45bfDRt/hXpbaIuW65UNSqf6w
MFLSzDo3tXPl+gHu3H19RSXX/m0QQcqCOqVg1ZBPhGM/ttodkbII9EV74nwxl8celAGn2wrUoDcT
1HcigkbQDOl1g6/vBJb8pSwqKzWCWK9SGzWYXSyiq4bOsycs1yE/D1E8r2QowqMkWwDD6TfgtBX4
r6cFDdm54vhkVG1hYn+O0gGDx/qYw/4wEZ453oWlee6DF7jgQJhfC4X3lYEM1KERRMYPz1MIrCKn
HiUAUk+tAY7YMlN01qz30Zj4xWEzxDTlhqUL68TVNDIMQ8J0xEGp1DDaqYi8PpO0KaNDpOfgcLX6
0DaMdub9HmN/1qB02RTgVOC2QjzFewoOjCWCDtFM4T8E+1icizWEOsLsaXU+kTzceZ38qVilsKmO
dYiW8QF+I/MdFKPqUxP1GhWkfN95GlGZkluF8q4Rb+4UoB9yVDszrgn4V9o1yT+9332aHYjOrsar
AFh7ieL66pPhHyWjApF0R+83PlUeuwDCp/g/duZclhHpMBxXdNPNFMqizbbMAT9G7+392EgFSbRf
cJ010CAE8v4K5vftpM59918o+2NYFZRydMorGxxWxpvpONZ/AZ3orqRq6LZppOBgi64L6HYWqAnK
iixMDctvAysj/GeQ0FPGbt6TX7UPxpWzTB06LTaAuQgkjeLmQEvQup4hSSUeLov0YPMWv//nfSiy
S3qHccQHroisbAMN+BnApI8YX9rrr1dpo8bSyiagjgAo8SU2JgtgkBgU1IiRhqi6OxBNIMgg7vf7
0r8KkBf8imOw6G+QSVpZwQ3iAesNzEnbfpcfktKBOOpiwIXe0hcI3rECBXq2fVm/658A2J7AtBdA
EtTtxrYuLLvVbgvxMRZiyf3Jbj0xiXybqhDupvdw/VHVasSJwAgWY9HUyu7OzJQWmZY3RPQniByf
YTaBWO3/qJuaL8q5uH/QEZWWBfcoJGRdaigd5XuzXUPs9ukYF7cG2DktaG0EpVA6vjvW5qS25fp0
ANUsYb67bzQvU7Y7HoLjLx6CR16EI8iZ2XZXFgfX+z8qcbtYk405hxYX0Xw/KNw/5ib5T/nSwkbX
m/1XhmE+sFI/3SSyscwdQfZ4w88hlqt19BlM/zAwUvAGrwNZGNmEd10mWrV3AVrABnjge0Udambk
MsnATSXNdJbVm5D6EgytSboL30lcsYOi9yrlElsv+BN8j46CVJHIqoi82sDffn19aD3JHtSJHXmC
cNy5c9DmWAxK4xKQ38HPNxoPB1yo1bbkkR3mwU324mir6yVfrZ05FgJQET+F827l2CZUURaqB5gN
ytljqhlq3vVI/fwTK7iWvzn6QfbVgit5mFNC/MdzTfEFqbx1BttUBQGerPrFQGUIIpc/BluMKjQo
pqZsCiwFwVeXiGDWog7c5MVGqAu+B2K2kz+IoBQsgwb4pLSj6e2YM3bvREYp8kZ4+VMCu6Hwflyg
gW3uvkVdLtuuO7OeQmnxF13+McPYnHhaiM4rcka8W+04m0/M+2EwVZQO8Uu+EoF8pp/te/bQoOtR
lF7C4FGjJAqtpOwzc2TCdAHwp4JpMWSxqVr96xxnevFfBUJgujxUBvDCYTm7x3Vyrg7bPzMz0B48
8l0Es7qPyOYeCACWCmp3QOz8j24nXsU5+dyAuchi6jaV/HuYj7lEyorYR7bwZzqq9hADhq3yMnor
PnBzUHD8xrbTleboXKwDzboFeNareiuUWDEswFNyIZCMLVJCSU569NNuc9QgK/7BXtSIz2CS2xNB
XujZIi4NVUQsrbW98h1c7ruDcQLVULH11EZPsSEMCgIzapqDILAQRZM3Mc8xqZCnzurE/7Q0abkS
enOtNhHzVCymjJl2dXCFGVrjbqSD+rFZgYSzyes3a3JEb75AEM4FfoeupBvZOA1b57569NAtE2p9
0xXEN58JXzI+j3Q3nSA9NKvWwLrmAA4/64dLChjxwlTB6xbbTkOqfLT73B7tIaHrlmMrhAZUi8XW
MTh3EPeSFWXYqSTGpCoIt/kL2badVycL8mqIwp53FElTaZZ9PU+Qxy3lTGsi3Ecm13Fvt723fOOK
J/+d2bVoKG0BjZfr20EEj9fORmy3dmg82XFzKBFd0BzpfUOCq5rDQ6KqU07GFVuSSt3NseN0vOkO
f/jxMXTtNHpHSyBvQDQHcYc9Ck5m4USgKxcYHHVjdrzjq8iPa+dkoA2zBv40mhDUpnZjvenQeGr6
IpgU7zkFODORik1R4Hx/vOpUf36DcC5hLMULDW5Kloo/eZ0vzgcDkvQzTe+ZM1LUBrBsNaXZ1x/O
9rYyr136G+wmifrocJytk2pXk/iE9ppXHrx5hdQBODmFXZBF0kJhqCgjhBX50b3rl9dhCCQACu/u
QF+xG3vP/Pvo7wLEOOB1YP6kQ5Pyx+C3JyNGTGpLBocp8gE8GnNVrYK3/Y9kZFtAr56zI9Qmojp3
uww7ZBkhRqRxh475l3p9l3q9ALLLfD/quOMUoaDs1YMehLWXXhXrtyMIYHqqtJMybDvPEbhRBt0z
28mWvBQ29eEG/wPlBDLwBbQPMjmAV5mwxlNsqf033JT6WC37I3oSVEmmxpfSps8fni6VnF17yW37
dVPQLUdItmOy3BRSQrJ68O4M0eJgjWX7JI/ty7bIyX3pq9s7OD1zQGMlCKSgtGdBJx2Ys9Q5KiBt
lfwBkhITiaeoY2W1esINPjC6oYxySTMY7gDJ0vfTV2FSVwCf/Su5iLVRqU2QS+6jjDtq2KyBte5A
1/ee+DaX39Tc7mKEoMXdkDsbRlbBvPEpnpiBwRM7r4YhzDeh4qsAcnpgLtN5UZ/wHPV0+iOm6YdI
YT4lOij45+d79ux2m4t8MLX0xH9HB5X4yff6clf3IVMto7bXzmkjmsUN64dfygnmx2SElBNA1CcF
az0tkARmt5YhDalq63DKn8gExw80hwrL09J6DKO7sF6spkOhNdSj5QnMtjFhXIJzfBUb0aQSirxn
9AAwLra1z5dhbtXziiDlOSqauC3f5ZBL58vA4mg3TImrYkd33P0xUmdfAnt29AwUFXY9xOvXFoLU
tS4J44X2mam3cNoW34nqiXfQj1/1yPkg/ntpBlicqD6IiPUXXq7nEgqi/XhkFjfuTPr0GXlbNWsH
uEa47FaEFAxcp+2tqH1zccAAB97uvFIu9b7VbtaSQjCVSHi8/EqwS0YV5oDYTYn07McOZllLxg/r
rvXTA3Vqf0SN85rWzqh8cw+F4vSU6UwGnThojgyPzJBfjOsIPr7TPWDnntLMYTumgBQ7f1h14c4A
uyIaUZcLVCI16YQb9qvyAc8l7E6Uh78+s7UQreuAMhBm+ctzF6ekkJ0Qf82HzUN8LE6mop/0HKAo
XkYK9NiI4zNi7oUuPGoq9dYKYP68tJIHaCH7YZSM9n99SIqycuHnGR6vYBXdQYaxQkaDWpDBS7pa
zpgAl0xfO5Y2XHis88LEzInOELrm+BdOfgVaKoaODjfe3oAkkMVh4l0lEKh3hj2vp+gmW8alDOOF
SPwydPbJYL5Ftgn8Oo1GUG0/XuF4o+uieifP/iFpEkb/9r/o3DtZBrkVWVjsDa9OG3bxdZiQ+NId
9yOxxhLvpJbpElVJdZQzkbReCERVKLMGJB+kRQTyx0UXSqLSi/2hCSVTKa3V6xE2BBXCsr2zSIMD
U7syEG9FfWWSe8yDYm+DzX70/0521QGOoc9/jqWNLWRtScEaMgde1r9Bb7M+CoxPrKl2H72viWQz
dROUKNzMqkSazooiw1eOgVeF1uYopGxPo5jb8QRzAwZmb3Xa7ybvEA3wjVP/ddoTGoMfL9JiYJrK
q05SQ+ESYy2qeEcotvRGo9jkUV+Ccco3YA97ibcKcJ8pn2+ufrCEMN9BDyPmz8AcmRD2rpNZGeeL
AlXPMrdeG/L3T5AG0gTGcq4Yft7qhJxqeRlplEWXs/LFWJYtIcUq1uK+9S4CFLj6giibgh1IW+zV
YJj9J7FtatZ6oXBnJAhalf5h/geHsbONGic5nHcY/zcmkYf3VrJkj2ZvAeMI2cmjWSzX5RxxAkSB
Sp4V5fraHzkUPXTKMz2t2d+Ygu4nZsdRuzb6rJEWFGLGL3zgTuG8ibV0JFWRq6lI9RdrvnPhsiDa
d1L6qDqIWx6qqCXJhxcxCH3HAUyBZYO+TQrFf6M+kq2QpgcomdmC6E8+YuQmsn1ZvmhaZ+EwsK3G
5fwRG17XwKyBjsQp0euI/5PfJbfm1HMuE09a2QvdyUibON69ngVX4jD9/zOo1d0MSZQigJMrSPqK
IvnpTHv9s3m2+UKJAjIfon9oovUG3iOYHJbCdOvhXaOZjc+PQ6m82/xj+F8kBp7U0StNppDIzDVG
+JsRNOst6xXT/P7Zk/Mer4Kpkssbo9DaxAUlbEtmBpZ9F5FCnyzMlTAMrqGM9uqErjIsGR/iNGz6
M+6QGpUI4Qj2PpGCk8z8EWF2FVeuoZRgOnX1m/e2SRh+fvg8O7uO2sS6Pgk7UruUw0MsnDNE7iMW
w+fg1Kqt3VmSbjdBLpnj7BDvJ636uoQPFPBQ8GwwKig6onGKY/EXXkzbB70ycWruYmkAbYoWyYtR
X1FRLmVXYe1JHzs4aBSZuoUBdpVnhCxUDE8WWJcgqW9mPNNyWAMLORYTl4wDi0JpzdXNn51ZdSO6
xXUnGY5/mt89vVrB1I28S9IPwBnwCde8clMkyZOPlLaMMm8J4MHQQwkbnv+S9GgLOSTPr5NT2+Sl
QFifdmYH/AlfTsIiwgdyu2cImIv14+sn8zzcAHLCkeiXQV71yZ4an0RqlDcji7BKIcuFg0/ZwZ7+
DI9F8K96vPtAd3hOf9T4SPZzZ6r2qJXYsJICGoBMZno/iXGTqoxd8g1S6bULkhCTfjHzrHZrooer
o8PYbqG/1X0SEl3NthS68NIGijYke6DxJK+52LbfVjzX+rtblHCCOQjPEhVtMrHIAnl6GpjoEVc9
fMxzI2D6u/wSWeQjcZAY8NWnyQdERd/spb51nB8QqnNLcY7hPm8kloYEHVBnFSTANsVdilso4eDh
QCtNl5Ci5eX9JOQ6XjjJaqoc/wpzpxoll4kTQouPGuSfPMm1Ng7i8xTJZVU12j5WhpTE00X9+bLg
GDQi6XALm/46lTOE3crsBM7VXeUyev9rge7QP/FD3bzJCiU3I5LIG+SuJiiXrp6S683WQ2s3M4hK
zFDghgAsSwgMYths2dSwY6ycrQme3l2n79KbrkZabChmdKPu7Y1ja9Jrdl368PrfuEK7/c3/j6Jx
iPj1rPzSHUkQHBIfzoHEf+YqQqea5BQCVFwUOilexqlqeDenUNPKRse9U5YjdEb4XsSGxlv62wyr
5NqADC/Of70W8lAYm8oioBnE9qTG/Nu7mo482gm8yK6vvye8xWGZ8G3f09n2g4R4jgPXpsrq4/e7
C8Y1B7Q0DsgMtgHxYWgoAdGgvnNfxSi0CTEZyNm98hrI88QG4fgasFW5c0LNB5xKLvYiKATsnlku
N5hd1Ay7cyo7uxXbcSPwVpEaChz3D+0KZZog18c3pCuXfHVODisuHyN5lfdpm2KDQ5o/ZMmqhsi7
0xlQm+TWf6f5AYgdSiqtoclwRHD3wIbZUNaiV7Zcmr9orc6umYA/3Npho/CgnAx5CPqKXkYFPp9b
8j5nib9QFuLz4YJwpzl/MWla5Fo1ZTiR8v8n4gmphb6DHwY6K/h7B1EvoGBUk3uFDGqw8iB9wXSq
Fa2F9Gen/Ykj1eMeVmROrv8QdnvYf3TjiB1Z4Jyn/t2bSA11LO1+SU5mHUF0ZOuE8fbIfzowzxUp
l8Y6C8/pYHJDAJRz8m6yyD0HH6ZYhgeWrgJiWzfC9VM7NFoTFtIWT7h9RC6WpGObOTImhSe5btxT
4ff5xsSdb3j+NOzwPQL2uvq2NE0xFdHDV/Ml3eCaYdTzd5f+eF9sO7ceg3UEMoPDUq1b9+/9GIUK
mBDncmQQMouYipsvWge8MX7CD7mSSfgGiIFPnxUdvUCQ7RdYwvx6lfETwPMOFXxO3dihBlxlM+Ln
Df5MyhXUSuMleOOFXKyQ7IZ5TnbTvs5aQgNTzrBv7syewzhyafCXNpBeIKfM1FZ/5wJV/Cfy5+ys
y6lmTFCTaFb0XB2xhcktx99iLRONfC+Za5evOeEkZQcJy0SYfyQ0RBGZYnXQoz8/0vBimlgi3RBC
lm/5np2qPNueztSf76Glto3Q+tcVsaGk22S40a8eimxqUbRXQjP74yDrTBos4iRMW21TaqUveSoo
l1jUQak53UVrw7qSjXy/J3iX0TYPQlfov61mpROnfiiewnfmz5DJnpndYlw4nBzQ32uGVtY1jh7f
F54vmZ/FHi6qGW647CP+eckxs27q3udWdRKtfXh+F7Kbwd4e5abI3Jm0tzlR5XpXnqwvIGcPef6r
Cls7y4Z/UyuMKWMp5nGscpRwPia1fCoKeEk1c/UJPfrVG/0cSwVENR1XV5a3iouTm2ZoUZ/3SLbe
Nlpths1iPsjzFrTYkaj4zlD5N4PLmxg8XChtm/e/2nEPOlhk5IU8fBSWORV6bszZGiiux0roXpyV
rHbi25ILBFd5FIv8l9BPMhrmkuNC0yBtyPc6/0MGnuYPHOzvE46u3ZAPRjNPLsJKUvSCIBVD5Uth
nrkAxn+Thd+sLLceJBufzWUJN6zj3SlcO0mA3mtfxEzS1OgUk10+jcIEOLtSTT4cyotK8gpq6yhx
4UDollRRlcWu3fM8SMiOHR9/8Lop+64N3azPvL+Pl2mVUOqC17yyGCpzufJJvhzPi4kKa+j4CLVH
8y6vw6OcUk/g/Jx5Zhs3TqU+PbyfWCHUBKxLcrl5WK0rFNDT9xuusm+DGDKHC2lmtvMpbBnBKXcm
wfCNCqZkNfdcwsIPp4bZJnQsvGse29YWMwVbOqWS4Ivbv+7rnzESU+gz7AyfykBrxcuTGuohWH1B
7tQLYaRotUWMhcv3FilHv6GI6DvtJ4osUjRGfjBBuaRMTgbWdzbz/KsOni1u7Az6YSelK565gdCw
GHJZdgmqtj46zEBpGOPjRggAKzj68Jantxazwwf1yOWmu5vIsM9mEAsq+GkIeBGOrboKXjy+HMRB
CVNYFp9faAH9fZDWJdHBX4L7GKzcK2ld4/WC6pej3I8CRI0Em+RSdtvwMzLITZw5p2CZ2qipQWRI
tLisst4G5cu8Gw+qGptaax6y3NlH84322umQxrXrHPZusaUW04EhuJJplHg1zybgtEmaTxFf4Wif
bl/yDUJVTaWEZ5SzTQWzJBcJY6p2urHZrUUMCMmy982yCwSU2VpdMUkVsaoAoZEnzZZmOHTGxyvi
AdU4Mr3IBCM9EBmH12DYndw3wilzB3syG7zU2z+snI54nety/QprHImY+W+2fq70kk0LhIeyi1Sd
Ldn8v/onaa7jBtJX6WqYfRF0DhRwG7wDbbBfp3Cr7czju1OurZsBNlhqG87ChRhferclNja/IqGL
CuJU22dBrZpvhUsAmQdAF62pj2w7xW8ea4kaj0OKu/7hwde6ZU30au5okh/az6M3hl876GWNnZCM
xf47xoqoM0OrA1gezrG1oeBFehuLTd381+PxK788UuWRl56fi2jNpveku5UZr2lXL8ekqDDlbJYp
H34ZkuCtwRrY13quwQLvxBzHpknqBm0X5zk6Be+FtCFYCgrhI1AYx4UcSOb2XppSC2Lgw7ZM1NY9
uIg5Ncl9/A3GKpEJfSs9UiOS9ZfhfK/0gl+Zr6vTbxAFC8lSmbstp0apEJ5s1vw1GtoJyqphiUdI
oZYjBN2iuwtcbhKSPKhiSW2oQrw7NJuqZpnYKnlvYyDAYY+xRagyTgDL5kGLtIQyW6PTsgqJjaWv
9SzeqImO57H/Jf010X7h2BiuLF1ODPFk5rn0+080o6VJx3nVCOw2w525wNZhjdPhBBTv6RaSaHo/
F58dwtuKLB8JtUfa0tuZtncFB8eDkkAPRfUEtxx+D615hkuIpWvNE0IWRSIBEYsdsuSjj2OcoSMV
D0xpPUgZoD6wj2E0lhpGXY5bUE4fD+W83mhZrgx4sF9ZMvM3Ndo7NNZmE49aKxlYJKSNyD29lyvj
XSUn0vtUrk3XfZAakVMy9RTgUxgG36A1Zuo10FXvgeB7IFVRZJsauFzNeeTEq5brpx9TlJaYWNlU
VRJmvlE/ZSpLtnC6OJnnFN8be6dr6824BxurZLid7QMo4uvgEf1CzVkgsUTo3y4uUwXIhHURXjP6
QoFqihqNiWCl62WZdNvZdaiUK5G9qZRcGbXWz2f4xcskEs390BsPaNJhZjIOs/48QuhaEp0vQOBs
w8X/nCtYhBj2d7UZd8KJjKIRPa8/jLPBJykMXIT4s5hDG9Lg2yZdXxwWFlfUNmHtfOuEA0KliPvj
DQBKRXz3ASR5UT2u5uZ4ViOJ8ijozWNxYjoIrMoS6j+S/jO7sMb0me7+4jNZQp6SW3nICcRH3klU
1xfcpFSsQpUlE1WA/Tx9fWB+LOcjOuHzEhZ8+x8VQs0B59ihzLGcH7U8IVl629W0e+cs3pkOKKNs
xNAzqNxFQxdU3BbItlY1nEoZL0yMW4QAVmC5dVglj/UoxjB1soZRfsz3cK8igCQuo812Ni94FsFX
cxezxUCC5938FC4g9B1bdXkONciF3ve6txdvGrS+2eC+rrIG+0jY4oeepoTBkF8qvXj+NcWMgvGx
wtE0c6LcyCYKzyToi0g8x6NQZr1L0sEiT6c8WNR691VU6tz6wsVRxA+E7x48J49y3cJbxazOLoH2
zyArEIhhplLjMMRDmqYCtus086J6K925SuREuJcLHqYxHFPoK6GCZ7/WIk/z09B2VFJUKdp3fk7f
zcXX5baBdz1XsLt9RWlLiR20DlilOwCgI9O5rVHQZT8L6lBdZn89KkTHPiEbYJ/br9VdAe5pKpTP
HVMNBWDlgE8IdnRxFNSmlvfQGI7WR9vtUkC5rfY4sp0gr3DMF2GLqLRHDMlRh8cf50hYer1jzNLt
+/HRtSZRAYoTGqPvnPc3cqZvrFyM91ZWeivn4fzEm7TDDlv0G5rKqtYWCFaJQgSbTDeSae3gS4Rw
VOMWY8/KD+OhKJ6spt96Kbr25+IZORbwKpA/1oC3saRgLm+DHZWaT3miYfAx7iR4kGA4sGysWIH5
p+iynjc8DRDFDcx9wHIhI5en/DSE1Hreum/Wp3aUe/D88/zRaq8RuBFjWQCd+R6mvwy0GEtN03Ue
O/J+pW5J2N9F87KF0xhxALNM6od85ob5uq2PgHiVhArD7BNwVqoPxmNohIa9j0K/Pnnnbvw98QfI
wZ8ey45DQN4KSQ9O72HQcZ6olfeN+SxdyR8z4vbCwEpG+8EgsxmS4N95AchoiRza7ddar2UGo7ne
fxJQBmA77iUrb5ExO06mQHulSMIj7lGLLYchPjfxNkq0JdXOB4M9sdc6mEsrTxpciDEatGUl+Emc
vJct7ywZpekonGnV88bwbBp+XHUJ+QRmxgYiEkq27blibCw8O3gwi2JxEAPz7QeVVrUswC3G7eiJ
7li68C87RMP7E1f6DiwFrpS7S9gMVFmXDkH81EVW41RBW1ghw6r7RK/TWgzOADaHZzoxkCP0sU+y
1krCFSdhCYKjR4mIJ+//vGws4ChfAb4XVLpRiFLAnrxNuTBKFSazC0Xf+JU0sHaGHS0WBcyyZfWX
j/MiHrZ+tt2YFWsxffPERhMYSYEdgte3I7b0GLfvPgTARtR9FazPEX7fR+G7I/ISovwRA4DVYUx7
3JUqdJVmCfIQUy9zw/sQb0yGTWiNfndjP3q6uhn1AGJW6lesB2PNTwKRmMTcD+w3K6OVK4GaG6JD
svCV0Wq4rKuuVaj6mx88ujloSPjgglzuw9pNST9rlFpZSJW0knySfWYziLiNh5QSOsJHd2kOA9/9
YKPAXOwpL9kPMjFcF1WhQaaSLU2qIIfOwdRQvkpbPN36j/cApglLcGJANS015bkXwqqg4i4VROzA
MT4KM2nBriaGq212jWWyqYqWrK1wzGZmtFSyqD7FqCHRy7sExXUV4QZ/CENbWf23te+cP6GI0S3S
Od55tFvw+8cmn+/oLAQNtbmmZdBW0pxQfNlmqFBO4GhRj6UR675wjc6dKdmyPuIdhWADyxF+SON3
smj87ZeCdXjsVnpE4eCdUI0uea/UwdeZD9OWppLNPcx0ZBjjwxwZ07ulXRcBxhC3/S+jOyZQeGW/
8/xopVanvjw1c5fh5BvGpxDw4HmXWLhZTDDNyBe5peA0t3nJkqsCCjkixmetPZXLVWE5Lv3vjj3q
Ro2UFCyuu66n339oX/Qy4CeCw+RUnu5uax9vUuZtBxLMKqY3hMJ3icAr7NUfuPeAztzVju5yfeQ3
Ty+FEU7d1u90iYjrmx/gAYYD2geP9Anef2+7O6Pttua17HLDTzAwrfz8Yum8gOdLZLBTpxQqmt8/
Ul1rQ9+G8BhwB32Oqs+maFAZmi/4fDqQbRctv99fYC/17mZEmxEcpKe7QvlahKfjuzLE5AkSA/Da
/Tth7trGdZ88fthgki8JXCTVz3Sf34JA9a3m8bfQuOrfdm3cp6kR31zg45O7KUS3OhvSXBjUKshc
oH61LJwfD2hcZa9L080Lp7CkEqTEaVIWz13ijAtZnqtu/ss2CLqud8Gpf4xelkJApuhImdbSyQKt
/iJnC/InU79f/y57qyCUlFLmSmFPm5eStVKy5HK03KrkO5Nz8gl4/VqhSy00QqGQhiuax+mPs5zM
hgAwgR5WagCP4W2DXhRIB0Q6gvslDqS6wq13zchHxnUvlpQempoteQ2n5RXT9DsSFSEmsCWFnwJF
pVo40KfcMlVMI4Tl28ibrY/CmjqSOvQwAC6G376yiyDI7V3jRrWVjPRp8G4CGLNOk/Ho20LZEWrd
S58OV4eG2k7A+iHDuP9MLiAh2un3ApIXKjsVahF75YsUnB5bw7Rt4RYn6qYyQeEXoGd8uTDUpYHd
n4/mMMhPglFrtrxVORmzkhtNPY6ZlKKOr01pqePDe8UDP/1vIaimqYqeXOUVwSM4AsoyRlGSyGjr
A0kkqVacNnaQUbsAdvDkA13Nu0jpZ50xbCioRmbc2imDtgcmqT7poDt0OaWbgWegWJiYPBfd8rkd
/QZpbvyQh1h9LIoXY06RaDe2D0IfSVpq1ss/E9iMQBRgr7aBYbtgsh4QspNodENq8uBdOlZkACZr
cgznrR/hwjOFjfarn9+uLXke/JVNNg10ILwOVYRaItVg1duvmSoM4cHk+ii4wysHB8bBES2kLic3
Xtl3HNfkFLHwBrgGgp3l+G4u7bQZCqxKl5NNRp8JVfka3SDRu0V/zVKv/EeLL9JdGwv5FXMDroPn
k4L9Qm0OB8r1TjDa4v44nnBSTjFoxPjCrkLiQCgIa4SaijsboFVq2RVzZIk0ZYEbNrar5OSjG5Of
iguUJJDOvoz4j8dcsnIij9PCbcWBlZShBBykXu1U5uGgrGndNHwm67Q3Pzqp6+NjgQBHkkkYgA+6
GIrF/BnuSKfB6kBiBxrosW0CKpZydtOT6DN8XmHZ3KSWEPMsVeIFVwbhPeQOjHdxJr8PLR34neCx
mQUD8FHLKJ3XQoHVBgJSQnknWPmTKfdm3dqrJV9Ul+3TE3PLYV57+3dmUEFyhiVolN1qJQgj+1cN
+Ix8+IVgBu13DQkLRsrfILhjMoVm3PGpSlwltRemHzzdk27lUArhBfs6KuIoUTZptY4aUZJxFVEK
ryRx4+VgG4BwSYcYB5Pj5c8Bosn/GIPc3oEI9Wf18+VLSkshHZMxmRa+VyGEvOrDHOlfyEZV/Bbp
NHquzAEOHn6TaC5wFOUtzlI83pyemd01EwSThwZYTvwPazVHkyI4IRNc+QSWXNvARLvea+84MrMf
bcSnAfHIdraqJwEZXaprFsD2eoxJAq40MVJIm0WdSeNnm+zSsTjYbRDv5svzc3C++dqL/txHO/nT
DPxzqRHNU9U74dZJL2IRJoZjx9NEoHYHIppbfCVcTC5TFBAi3QyDiCFzHw8vRNPEsWWn/JGJOD15
QMJfE95tjOhR/E1ApiXHk+rHtW17OlcpHSbivD3A1Fao2I1HvWWaNmKXlO7uYgVRgzfc/LtXuSod
sDBwPhSSmsBsiTpAkV4x+TRrhrlEpjFQBVGWgS+T6+cACJNOzajE6l/gd1xQrOxr4WzAc65j63NB
i5848hE8bLBrJ1gibB8MP2tkbpmnviBbJI9swjk9hbdmU1kIH2BZdrBwaGjS3CzZE4woObnz9mmB
MPvPytpHrRDQKtNxV44N22jOVaf6nT5fP9yV5xzrdfuEHK4Sj0DediN0eVDmXCY7mtXUOeIrg+4e
d5Pqagyi/y07lPmxylbJ3WujW8m2JBZcYExUbhR4WPNb/YLVU95ZgTZImc4OHY0GGJhl8vh102Fy
4DColT+FnT1Z7HeRgxL8h/CiYs8C1TGhvTrY0G2pvsKRy8n9TlbORu2XQwcK5cZNqCwtDvR8h8PK
mYUNWYVMLej5wHE88vTyCNp+XdTDVHmtGyMIoIS6+VdwPBULXWpbui2uT4cSO4tswnicLReX7DFO
R5ntXfvkA8+JSjo1dsknGO9eWcit4aGPlQjuxa87eGp39O4c8FQcVEHyL7ar1rysGhV/TBLhBff2
K8pMh5sB/drG1UItRGDDwdCbDLSbjQnQHZXKDY4XdQBO8OllNZ+k0249VgOgr5fhmq4sWw1dXOes
dTKX6pFvXnV1B1T3IgaDBMX4JDQngmR7sTCgAp9gwzhpNXz9LoeWFadUt288/5hq0RtgJNlKPQZN
/b1dm9vOx5UeyISCBqaimXimzSF3DfRgQtPonpCLz+gain4E4LbHHQy6tJ73CNSvpvo6d2Vl20fP
Lhb54FPjf2ZhXGNOjAyoDGhe+B3symMBfh0MpHHLXu9MkTj2uG+g6rNlsOOwZXn0fUYhvV9MYzBO
4aHI0Wk6smcTr7RUPYooxDkM9r2D1v7JYpXEbZ6TzjB8HaKc4N2svWVaUpK4Zn4p3SFZalLdjfk6
w6dQCzPc9FzdXKKiiEVwn6Gc8jCNgZtPkTdqMGsaQNP3+x1nDvmrRTjTBRLFciKZELjrMQdkJFQI
RKXDhL4HqGJ9vHcdtynm8TUnrjGWIl9ZsdqrzK9dobXIhNt8mXoRkwGMbf5Iy9ZTLVSqCkrCF0Ji
UYsNTYJrTFNcJRQ1t+6QpZE54OdkhKWZbV5AvcKN2QKm+kgAQ4kfyYXu5P9Ju7117QG9NEtdwU7/
Sw6/XrQrAOmbZvns5CzrcNJNy1cOQHAsYCITmHhRkZEW67dD6uv9nEifomNbPdUQRgta0hbYWV2k
RO1eq3boZ8IYYxIOpB1Kl3QIOwToYvVNLyahFcq+8uUPbFdoketQwRP1/WlCjZJu34wzRgtBFCy/
/xgWpX3BAF+Ey8w5v3ApttYlYZ5ioI01oyYCTLqkCrAKe4rQ7/A6Hoh9HWVZr6yZp4PbSppwIbI4
q3xRoWVqKyzRLVQLCpbNkEISg8FCv5emGiVh4rbDGCGr5H1yslJOmz8gBZNtV2Y1md/BemCF4Z7/
Tn9UcxeRIq1Wabs1hmmlt4DvvVAcgyqb2Z1wM9nv1JyBltB5Yc1XTNcksEyUvz3Rb5g8zBQZItvE
+9Kg4J6iQ/XCYwAKORk61E/o4JnIUjfRM3OOaEHCLQcRnU7U63T7L0YFf6bGq2giNYSEUNXEkkgt
4L4TJeYiCN0+qFqfBZD2+0mJkakzubgqP5Y34uUrk3RyodVkHdKN6+5d+qa5EGGJ6xNtGabsN9re
5eHwfyB2QmEy4N33ynfTdbp3fjpLLIVETXa23//NbsU3yheyE6GCZ5Hs7Nn2h6lVC4vHucdYjvCi
s2UQ0RsBsvMY0uHGIIDnRl9tyaKVhGsLCwv1D9FX7Mlpk+rEEZrgP0E9HUY8M5adnrtjzrqsVHoW
8s6FsLevuyISXF+OKqmyjRpNJUy/3j1Qvg4+4Iu16t13PPyAX22eeoLsulq/6XXavC+b7YIFj5vY
ZHXbmwkQFTiVpbCpVt6RK1+VZ7T4DS09ijLCfxPxJYAEwa47P+jA7HzceS8C9zO+CexkLFTBfnQ1
wgwYK8eiqH2f1MPm4PagIyTxGXmq0Yhg6G929/D4DmheB4CZKhNv642lsWddlGR/RBSfOoJiOT7v
nA8iAjYAT5ivPKVWxJnYCa1FvVT179VmIY2jfqAsYZhwBQshkPs9VXlGFRvLlxd1QAuDYvpX616e
J0wvSYosgG6ttAY2XTnaUTIiRylrwgmTkSMOTBVDpDucyZWci4BZj/xBvRryZsQI4IFSMVenSYL0
6ANdS99blfTY7Gjo14Mm0vGZ1gzHOduG6/6oblJL043y9xdUUP5RYaG8+szL03XZtQQhyvwBpmZL
0ytg/tHIPgN2ZJJ/jvISr1s1UDlN5tvyte/N/aqmrQ3qRnT8fk8b4nyBNy8mbC9Ai8POKL1eKMR+
2ELWgqgsHFDmKrXOFk0Jk7RPzr83b+MTgWOP0W1bZpcFkxvvW0Cq62qvzSbyCB1Dab4KPjobKbds
3UdAOtle7XJrdfgxlIhrSgE5lRWUF2NxB3dh+vWNGuVg9guAZjhIzgIUAGD6xPYTVnqnzG0ooYIs
z7BapOyofIbcmGW+AlTLYxtfP2dixwcBLgRT2WNV6mzCL920R+WMfgvfnIyGj1zrRm02hbAA/A3i
Wmr3fXUcW3opqpGdiC5ebRKTzBaU4vrOHNFojhFw1g+wktWG24Tjl0ykb1lL4kfuotAi3scpi1YT
IfCshlL0BS1Ue1m1eNu7Z5+ZpE/rBdXqVN6VtTypdWYZjqI4oOvQj/8p/4CnXOhKGo4p+AA1Pk1p
YhrQk0te9LGXTs4FRxCoXQxZfqLJu/L3MNygpZQmBokAMZ51zLGtH20U0Y/R7hTlMqHR/lsfkWaj
o6Eiq6x2g+ff86mXB5iYDtw1MshEB20IsCQwLlhATb4wh0UMaJOB5vcBia30QS0Vy82lxtKE3NQE
bMJjhXDL81mHm3M59Pxhw19SIuPYpYvTw3cxkF7Whhf1Hc4VPRYWG45ieUGTXhvNY1Y3Um47hKL6
fkgZNGWSQlzfCSr1hdPuRTPruUQB+9fkdhQ25sj77xUByOqUoFzNpCop9gkQgoTKX6st4Hzh3Q8i
3hyKrpQeXMbwLCu3MJIE0A8q0bH3K/1QUOzRr0m3NARbPSP2TkfMlxCNLMq5iZ9+sdMcsxE41Pii
jdnv4UA5SHg9aVMN3r26630ii6yB76YUOaG3x9epjF0ti2zEeOt92BaR4UzfCWx8sBMOXSB+dDJA
dQ7hMMLbawJ2dGmzffSyacOm8QnryRn1cx6ljch5OImFXDWCDwyFo17u4CpSqo3Besko9Ljs0wzO
FS/cvJ4u/Xw4GbxHstlRqp3YNzG6tBL83oWEfYnOPz5tgz4E0E9363NACDMn/5vXO3EycR9is1Pm
C24rRtlOXid5Ij/Fn2eRgUcwa1+vw3V5nqeQT8g4a07hVcgJqQmH8PRR1KIzeims6QsIPqLoXkQy
cdyeIKz81bkqn78RDR2DPUOPK90w2AmjMq4puVBWMNxrgAOWdteQ6fqwd442J0WHJbxKvRO8e5fM
dCXX2tbndAedP6E/qtcU7z/ELDn5h9FazsVxyexzV4bK4YndMFEMnaxdA1HPQYzlRJDuHdc0oigo
/MRXCspg+x4zn+Vn6AepKrai2G0Ha4thW3Y6Wa5VQ97jjvv+IEIY+ey1ssRHC7X0EBcUjQVfMGi/
SP6ipfV396f7H/TYmVhdg1O4debqI8Ayk+8cCW9+R2mK8JwmrsVzX+Pfan5WRhubZwBwi4FMzfEJ
sscCb40fOmQvtnKpWDk3cRBzYCxrAGxRv3YNNsIUIcy7FQLIju2PI5POR+9rxRlexI0wKN8OW+rZ
pRFPPwbRO7bmicyWkuTcVPsWOvh3l2vGMSS7ddkKpL6F3vk8wyU+T1dupMlDBkt6BE9vkRPtrpp1
npg4scxb2YGLfmicLAAEIwOhm7jsJd9+OAzNxhOeR9LlYL0YNozU+Z6G3kmSNUp0c1nGFqUR7c6p
xKNSoCZgA9pe6cr8rJRE7aN8y9Hs439rnID2dr7QwlViiqBBUTcH0e0DpmdAkEfFVhBFzGMIrimZ
F4/A8JU5QkLm1F87KgK97QuUjt2aWK/cDQdZsAzFzgv5OV9WfUyGkml5luOHut7gQfyJFndR0eys
HkPu1KRXVO9ydLbqF3+EnEzHfH58osDpwY8ubruK9F42BKh6L1/xSBoAksebhE0n/gmyymUcRHhL
ES61b1XkXmRoLb1R2/tvGae6m3/RVF6wavzosuUFgr+wM7GnMx1dCw3k9X73z3fFY5oGlsAi1tRe
pbV/rRotmiVFQOpiXcp4VnjJyz/3RwH/JK/YWoH8xr0dLvwlQta0Z0LPptOvQ/Ppl2wg1sVL3cOG
AdgomCI53jngt4piXcrpXSy49/sBkg+8aO0WEdqbBx8eyvvAl6XCJT99X5oykiUHF1cTLXTFCycP
DX14dr0URPi8QXdQ/9gQY7BEuv1yB2VshPzHr9rtU5nfFUQz6moj6bEiSsFkmjGd70xTDy+V/3Tr
z5d/VP22Y8tZCqeQwK/tdXCyxPswkYo7fsvDiG9QHAlsjih9Uhfori+vOmvoyoJ6Kscvk2AnITkP
yJesGogfiznwiZe92Af+5i9JzWisRk2D8C2/sVX7ECAwe49CsI6opvFC1/rv9ACR4Ntj7g6o5XBQ
CPH0cnzZA4PToMsdGUm/x6GlWCwqezrH6WV/s9HvTKBGqqqACcihPn88N2Cil5PG9s6Q9kkLFNJU
1XLIbkpOzy4+PL4ZXe5UUl3bhRxa0ay9auYTdag/2IRnSfl5V+vbSuDNrLPcKqd1UcCogRDbhuwa
MClXAgZn/aDor0yKQwt+atzaTlWav6Q7dcTn455F5Wy1cp0vB8mHkLyQElEaCXY9spI5VZvY0knJ
TZij0pYloGG8gpU2xZeC9QTgVpdcn9ZKOhwk/R4nAwjRN4o57poEZ1Iue/nnh43pmWRJHOHo3pXq
lxp+25T7wEhjHGPBaa6Fb3F37ylwpPpAroPJnHWIRlE75zfGjDESQjVLIo+CemgkLZYmIDzXb0EW
cbAj5gLW04oWwOQub2Rxx2oiaACRVDqG128xDCHtNX1K5rMTFccUcBmGMge/3tmSWb93bzIhlCg9
RX1MhytD0r9QJiYps5iyELJW5hGHF3aeujIA072LfdvUJo7V9cJWQxn+4Brj9smmHiA2oZc6W4ss
1WKwgt/RQtt0bVrGBKOtz3UJKH7E3CfMEG0i/ADN1YdGtXAkMJMR4oOiznXK0P53aulymJ1AucTc
dktPbLqbsKHVHD9ENOUKrkZhm85aR4ThZwjt0kT/NdjfScST20ymxVGCZ6O72R8YgF8+9TFKqijl
iyWdN3ABAu4MtP3KlYWgw82GDdsb+wRiyQQXZeB/H7dKb+owkNXXYUSh1LiiytXnurvgmzbta5K5
l8pPKkRrPg5aBx5wR970K+hp4smRXgZK10BzfVdsRpHfXM04/aR+xDB/7j+630kvaK2L5mf7pK9P
CJ3W8zKfHOSHr/ikXiEY6+yTXbeHgTAdFEkqAJ/mqwluExDtr/yEtaFYDd+ty9J3+sGxnRmrUYHf
y70w7rBLUZ2OUjMBJSUDqnMjTa46xLnnxcLn/UyAput7Uqt5cT8vqeJWtHn3NrrmSW3i3Qxw6zqt
Ple7T2rGWXZcqvu4BV7fYmooXHVx7BScBUbkhRoV9gX4a72LhH/j84neSbZ/pfi6BX33Zbz9zFIH
HW0RNRZ4eTleKhBLW2ujkyMCb4EQPwuv0v0z4r4um6T6Hbz04Rzwkfoh7xFCFHEkmcoiMFpiP03l
EV3rnU5r1abfQTcYfOnWC6NnCZREAd/O+4Aq8Q6lNpBwZUKUwIAZBTc7UZwPhcvVZdfkkf4ausGD
vq3zZ+vuMq/kYqYV4r2NFTrMweUduZCKkBVDxEyo7p07AUcuzqOzJW/eeoB6XfTHopeVYnlOrLNT
E01zxAjzP+L1Le5l8IHr1sQy4+KSwk94PVsGj1Vi7YMHtji0Tawd2yX+Jhj3V4M64RQNHP9EYjyK
1uZ6SNAU4yqTPPk90nQQ5DfdUx9EhvEDyUqPfY9DYPGypq+PTO04oYibR+r4rbkbeGIwwm8vbjWc
yO4qWn0PHgauRYpf7ojonOuJzr/c9zRhoeRU6t67wS95zA5QL5uAggobO+9OF7qV7cHCSD+AENkf
vZU1USFndRq56gEC4XTx5u0UA6tX8szjOPA35dsphzzL8UBq6jswiYzDV5t+rB2/RSD9TfR75L4b
NltX5fu7s6avLMoIxb39HO2TmCBEZCnAD02qMXWtz7NazpM5JSsK3ooUA+AmZdHb9Ep8W/h04fWz
8tfk/z+bHu8QMPnyGBSodtZnMukKUjoodaUz3/uGdRzk+BugoVJio5nHFyBH6f5nC0vEEqhav9k/
lqZUL/bIhUNIP/37gOwho1Mi/vsBwjunHYqKIT8bfOdyKNIU35VrRCVytRmV+QDs7xN9KjG36Dsd
tQIVXqkYofX96Sm8wqRVWzhTgChZC1LSJipKm9gQsVH0A2UFMrP/eAcY3aM5whiUcNHYU6VxTIvA
ItE2mZKusyxFojBQ69cQBe2DdPM+DvJYlwstyCHir01Zgup8p0seZdya55mw/lZIYDcpzUmlfg8a
INUwRQbITDrhuY179IIzsr9VluMgVnZzruqrYB8eS7GSXEVF6WqDcfop1uggnLLiD8x76jxwtWQn
gJnDK9JSha5NlBf/dmVuZBERlATMQP9jB5I1Ore27kI7MxUJ34CffU5TzOzP3Hsn0sR5atfJeaxa
3Hgp2gWe4XkZlcLJiNy9DgFV0zEgsJ1394kYAdfcQQExH1hdG4Gt6sbNwXWPzc1OJPyr7fGnhZFT
df0EFvWULtwAYOusn+ZuVnG5SbBdBGc3uC/bSN3fvtuu9CeQcEbovftgTASIkQR0/f2kLTdguZHU
5+g1V0nL1xbHFLSJg3EXMFUe/IBEDA0xAer8yCBQhGKFvcROJH0Y9BpNspdvLuCxAh4ejudifKJJ
mcrDaNdVvrUAf/pZJ8T9Rb49rmHJlDFF+uHhriMebOe9FazDwz0XxMGVizkgFXCNtyEpyl2wBMaJ
DJDyCNHfv5JCzhV4wwFmsh5I2n75HID+DfUu1QcxA+e6nPr1QasKRtFdxMTAK3mwLoJf6w9mKfJo
a64y7U8TOTs20oU0iTNaeBbc8zjx4gXG8CJz0XKjSHqYtSJxRRo1WXpKHW+K759LZ3cVlO8qm6lt
ijtMAsHPCaupJ88LtmAOGzq7RFb/oGSalxoDQXMdD/xHB7wW/KQuQxlogTAAKCCibFhxTpH8ASf+
KmWhvIqL84AqYVpJcIV/ClmwM/s7ge2VYEoNAW2M8/VlNPEvRR5NXgacB/TmC+X1lMvkzqwW3/Lv
jx7pPbpYGhdH6uqyHczqqjGiG1qap3GBBzJY3q8hLk4DkFjwQguQRPdcQZMZCO86OhFAsWsmBH35
2wiKtbXosG0O1t+g4Nun7lOlV4uPaY7UVC3alFsfkIaiYCPiv8dzLmvQBNbdzl7KF+2K7PdF+VQK
SxkmzEzecw+sj35lJhT425snCNpWQ5qmxyya2zLau10OMO2PxKWF6ZZQujKkTe7bbQJhUr6PdgO8
6rSrwOvqQabEDHLZ9vB+Tytoep287VrnlBasGZJDUVzlWQi1kBTyLoIjSYgA003Z1UmXcb5B4QHT
npCo82nZMx6JpGKzsnhn+yKKNITUAcXxn+R0XWquUhlvWk9qS+BM3RuKZ1XkktzlNo8aZT8+CGTG
iw9SzxlJWq9PHK4DGWuj5nCDjz6NbVbrd+UbTfnqILf20iCPK9IYI1dim6XqfPj934uMFwxaFi3J
ndDujlOWp/NMqjQzoU3SjZs5O/61pzWXT6xFGDj6t4tB2L9iWdAFaXZTzOMQTdu91kgRicj2ncOY
CBKlfSYOfY6W/vRMaH4ARH1qJ1vKFvRN77OwJX3DOPEgTC290CSxCoNsbH7NC8KqN2Jsm4TZ07RV
Y9DfUXmqutiVEcWBhOVwW1gBHbg7kQHDqQ4CJ9FXk3X0VQ3aSbLIA1C4oiwMt7WQrgymKKGYJs9H
utck7HC9ED38BybWqBNbp1N0oDmu2nZLm37NqEUoXBd6jf0xNg/Hs2xYaBHr+46wyoYRWuzhn9nF
PSZA2Fqi+jWxMoo4RQoK95N0aUxvR1307lWsMipJ+QJslTtzROatglESR4hJ1cJbssPHqjrU+OHv
o4z75AO0jKIvjTcSE/pDRCZYatfnwAU9T9Cg6VbqCY/Khx2UjnAfxQKzotssKiLVGmTzGE2MkBNl
moLkb5MBQ/Ms4qc+wm7K5nHVZgrYmEB9dzMNmtaa3lAxD8t/St4Jb8QMcoL1uSICahzc+UX5E3G5
T9AKxh/C5+64xp9u8O2j4KMYXxe5WVWST7Q8toEyOQUwdABPSrsz/pd7YeLk/uMdPRHb8VnlnN0d
2I/1x1L2zgYEH4+KV2Xp7yXqA5Xw2Cd0dMOZeMBa/ri1agTmezm/DcXeki6mRSpVfPjJ7y/gAEXh
fEJOKRTeC0lOxRz1xQOA/E2cY7DXkfoNR83ac2GgsZIgfQX0pGqHMxJdcvVSsWwqSsUGagtDgeIf
oowR3K4PNid9j4awRUNc9Qm6JdDGgrAsDwErED9SSnLlR44pyECAiYNni65EsAyjhNKPgNJTYjYT
B6BcKi9aMvaVs8J4CThBdEU1wQfkRj8GQPOM1AllvvmCSpZGbLEbCXvfMPEfaM048BS1oVmA6tnA
rAfyMlO41Dj5O2RR8EbbEow9BkZv57sK0+5xQDlobYd2ry3lyIrI9idP+sodrqYG7IkWOO5BLxoq
0tHQ+gTPCnOHryuJ1aertU7r8g04Xvptwbv/Gg8Bq/dN9Lrer1ZFNrM4A3fBMZKmvo4FvsSHtDIJ
8hUR9Nke2Wk8sAcYmaE08MEYW81GbNdpa9UEKiBN1luu2mrpDFTZDo/r0FdQXfxIEp5Fm8KjOaG0
3mO0xq21OFKE8uNskAgUl09Wg5QFORPpPpVdQvva1l3FVzyCMriU7nIGSIhwiSlDcusKAMOGuk9/
DZ7LHsnjSt0Qsu7dgjge3rTfbWBh4sdvC0hlggwpdkD1/K5E8Z/lDFqTXItZ4/ng6boQBldpP9WB
RzCagLZgBwHTgXv8/nz1m96BqAsBuM9WfBliBJp2PpMA9KiC4EUOPCJktO91wP2vIig7hcpmihuz
lH0k3nbgstOJFFEotKMspBexUMSxuTlA3Fmd+AoEhEWsfmaKIvR88XDkrPLLDAI35x/66r9QI3rl
kvIdKrxqmdefWX6qeO/AOi1iS1zpe2HokdwbmEIdJlMn8FVMt8860ozdyk9ijkiyzo7Mo4kco7wv
3g9g/+QjJzaUimQVsHkBILnCG0fFATnzm0dl5qlYBUR2o91F02JH+j+RIu7UerVehd34I5EyPnnv
sFUvDL4sCsitnJDdaxhSYYoe07SaJapxApf7l0QghIkK58iengBndCD01Vnvug1FcFZUoAwZusrx
YfI3BzBy+szOAeO3IkidC6BsujPcCBwL4AHt/g+T69+dwdWYFle6i//FPC1gAl6DVcYuTogqkLih
YckLvmTdyzoWWl/Yrfw42p3AFbQE7ZqN9UydleV9oOi61LjcPjTh5INsnARgZdgIecn2XLTIvntM
grkpY11BeesXkJuyPEIQMrKaJIJDnrootXbVMdETUiFxAxPVdhbADTtGYpmsrGpHpL3kvc3yayM0
qUViMWH72c1++3Osyn/PGWhNMyeBx/FyQmgwEst34tDrjDIT/re+bQsEkkxV+SOKC1KHXPon++Fz
acm5hCB082ygPKwsz4mz4yyUeLxVDYRQmo4DVLXLuBcIXtwxl1x719OZBj+Z0WhkAm5FalB59el2
YdnEL5wyKasFOWEqijD9RaqHOWKI3Sn06w2DLDs0JlL39MICITuN4SrtpNjNOMTXIgNUa52yiPBd
/CLyie0EhFYFWjrte4NQHl6Chy+PX7htKle8Kac5Zncs9vS8Jjfz3hMrqxtKLxqhc5Vk2rPvggg2
R8mr8TAPGmnBDJ9zo0oJMoHoh6OpXpoET630x0t+OtOjIIXEZnEBiW+p2/LspXP9vujlrY5gjiVo
fQq8rawdS7FNrr2xpCXX0Cz4UVJqucZf44ySKbjmOdIf0hxYPK9xCr4SD4gcz9bL7uDo9p0uvnTy
lMhWbByiuEfdcUe8oWIzfPPCaA7RpPg0zZemeuGGa8FPb9WmAYO2IR6g66zM2fXKzCwEf+jsYYhP
NS/fZPN3t4uPSnLRPbbMF2xaHEsbPDz7cOic+SnYWQrD3N9LWTV5nRy9CKXT7n2KT/FmZX11QlRm
u+gBqdkWrhUjbfhdodCIcIhGYOrVtxiD6UOxfeWpLxtKoUGA+GZPdChy1AuynHJuB3s+wfDnEZY5
EJEuilmpoluAITaCo4La+CG8apJDKUi8MjhVwD9btO6FOyvbPyyRZSVXVvNui1aNIWRONLbwL7rT
4xeSuJ1MeRxchf5nkbwOt0NiYMbqV6NJNWkqJXVHlzaAoi/hemGeFaPpBMW+B0olVIvxtwipZudB
HU8BACTHPN/iK5EsQ1G7l5+27qdKYt/xWb+fNY14Kt21GhcSICrMZtRxzHSyuPEhm8fMKeX+nmO5
IZPX3wlPtWG9/J8JtffhDgO4FvW+BLxiuS141yhsWZOeqdsOzbmW9Tg2iAUqdkSCFyTb8PqgA/cd
n4yae01K4kXk4Qfzzz/ii3Mx0Y9p6K41aJ5njO/akE/u7E00syq+Is6BWEdpfhA+yU4F/VbTH5hK
g/5Mv2mMkudlZ4Em0X/dHj0b38Tf6Kg5iQ2X6VJx1ArrhF/3qw7+FQIU6UW9NvnYBj+lxqFkLW+p
nVUteZQbkVTx1dUDH8XwvmQkIziM0a41EExW79GXjbCccJpHs17RUMHRwuWRYkuyPM7TB+u/Bgmh
zvCCLAx95b/YGNGceyTSWPCSb31NY+JNSDHEHoUjeHC7tK06y8mhKXgE1wZ/pT+MXBhUn4EW2M4F
g0fUa6eCAbmnS+XnAtIyeoi5ZVNJa8XUMymeAwvFChIDTBUU/TiRAnrp9uHZlG+jUkMRnqTrHNKA
TIOuFBxsXrJ0kHiLD4EJcrrcOhAZI+tBRNjjmRNkvk85back6S46cDCBTFLQ5uVoH2QPDRK+zaiu
wq61fUOi+84lDwIL0LYNu/oJs9zkzQW+VbDUcZ3d4aoUlmIVYKNByOuJTsHs1tUX/52lfRDUSKvb
PCXST+T+7aOJ61o3kkLhmOLnDF6KjGNBv7TLJyGEU6ImgRehJo14MfPYht1G0wmsBat0BWFCOC92
BgQE5QCc/3EFz8cvp9CFmWfpd8R82yXIPCtzoeh28DUd+udPfYK4YZa1hVRIhBalW+Bp+T3QV2ze
9VpQ5glrXLATDgePxbO/GrSVUasEwTFMewictneuDN46zpNZLiol6jfr45Bo8nuwvrrAEP1ptefw
0WjIEqO5kI7jx9llixhKz4jDqQLdQL3g6x00Dgn/qOT6d235EbcVHBN+4F87HWLxK7r/PHu3xsoa
hRpYpp0VqtNsarap1N3Fsw/rmgjyT1VTgPjlPGXp1DEkNt7CpfMIVAnpRfySEEkJ+7MlurjGFcF8
q0CGeF7PeJPetNB8Oz9E0rkcI6E4HFNKVwmT94BJBKOgIRlgLL87UJVQgL2ovt1Uga3ZY9SpJHeD
VCjvJhUK410ZLU/SzvCKhbzO2ModI0zect6Ax9NUN0L6jbsVOBShCxZCujyvJmfEhQOtHlfge/Cu
/CLICVpjKVRLdYa10w/aw7qmHL4ZQYyxM0ZAtQrISWxHr0jMUaquucZJY8nNOWit1O/dbrddZ4Av
nM7nK+eZUGRh5abehjxNMvKW5yv9OMUDp43EUgrhTgrYVY/bsS7rzifBGMizip5AQlhFcJE8/dhf
WI8Ca/WkMZscJ1hf1Wv1OjXaRJLPivPDpZa3M/iRZJTPNEkCzgoNAs3HP3HoDX9DFA/UcCsFgnIJ
BPgQkvOCUAycSq9mBJ03UbINpHGA9R0yZBClcGCVWEM0UdYe6PdYjpGP+zKheSLPyrqsPb2kZClp
NPnbGFtJBa7GI8D9haqAKBYMeBNvzmiuV6h8dClEPWosifB/fMLUaIWpJK1W7as4Q0oqRaUxUL6B
9U0XtRJD7uouKU9TEjQBesuijNexykRjNdRbvB/0MmnM+fUmO7lpvzP615JgACZisbKYzlgQOKZB
M+6oKU6dWzgWNlhcHZo+poy2zAQRpVtsP3aAlfXri30f6qOXsynQOg1/FcGGvS3L4EePtw2/dS8S
Jxg+ndTiFSac6u5gdh4JHyOg9PtjHImRICr/vb/Cx3MvNkfhLoRD8H1bBsYyEVcipIs7kZ4PUzzH
M1GIcFZQkTkwSuZQRwW6wp38kWX/CKfOd1vfJd/XsIqBQt/ay4Vh3BU8sOOmhittVetqE5RoFBxE
y1IbpIaQRxje+pfdlOAEt0j6p7DSs4Dk+7Ki8KHchktctDzzJG+isKuneO0o5cwMjSSJoTZQhn+7
TpLWfrhDdchG7KYzkRDA4CXBkBPZu1+tAByfPKtAdIsTnW9vcALshHhNZ01rsv74o/BhrfsPfsvf
5iJx55LHsWj0K1xjQQVKux8IQ9apPjJ6BAPyeM+8ty0j9rRlWRHyXkheeSdrGX4PxulbKXndqHMd
phjJh5YvkLKTKrIQc1KL59h0WcD1oW83aYcNc33ZhEsFIAMNf8tkiNGc4/fqWKEz1e1TkQOZRiSb
QNO3teKHomPJKz6zQ1A4B0NNNxnsC4iR858LL+Zm6mc0zNHCSz713Bh48rdmIPemM5+JsuX6SK+M
sPqGdMECzoaRC/lGGgMiCt4gEE3bkhaDDWYX6mqKGLGW3xTYAEk5a/8l9I5WDommp9hcBSnwh1Sg
3AiF8smhznBGZan/4k8raj0TTsCe2ctgq2NSyV+PLEabu0IBn0cfsc3Q00HZE29ibCaOn22RpD1m
eLZ9j1GqhvPQqIaUSoiW0qUABIoQsdeuIioZ6eeMfh1R2BYNnhQ0rm2O6H3duj/WN5q0iZU/cMqi
oRDVuvUEnnvl4APC6zea9HKlvnh9Z+v5T0XK3ggXb7hNWNC/YZMBKFcqdmD9Up4/nD8Cru+cRoBQ
BbAPz7osZs5jfEUvK8rnFYHOl5mLsaSdbjKoZoW4WfqSmTI17WdFweBr7MYARTR5eIsF/Mfg0Ixf
iMGHATIVMzvyGPto/0p4z4WyQH8nP7k3SPEPHh3n85XDwwcBg/no+j/4j7zF2ZFntaqTEkfxUwti
GvBbvOUIWaIdZ6h2WAaYPWmC+ZpaehPLUU3BnJpv2dbwRdaH8b7kpo1wZFWoFpCnCqwWDgnd9Y6z
oTc4AbzS6P9rzY2rMntnYuDgZ/AkKxGF5u+NcSdkSkr6G1i50YFKxjyPz7Wc6N1BRpoMU/kiiJCj
ezscIP3gk1bquJKYQXIm0hKsgGWIF/bfIgjloAPQ6o2dX/seGd51VRLPdHrzaFY7GLeiT1gTF7+1
hClAmjnnqawI93dRP98lo79f+nCljP3+xWJ4WLGtVMG5D8jFptQPw56d46pofEtopw50WxBvttWc
7WrkzTJUYA4czZDm1LTmJWe83ZtoBUPTVUNTJkDf4T2a28JlbrYWrUQf2KlIVw24xjPrk/R/lRfu
JJYemCUZ6usXdOqI7X/dLH51Zr/puC/orFX3xARwOEo9MSSUt5H4jogPcoKabFRuOeJFTWccJl9f
XjvI6NifEPpXHAMxBHNdy8HEdkcuMQOIs3qYo6bKpOjbhxaaapual0O0aCkBwkj9JDsKNkiSyqp4
NMIODxC5+zHxheBN74hzgYh41TsV6XM6hRVpvPGfUuL7YOOu0qg2n2Ez6I+oFOrHolDgFYpeAPeK
iD3afPlCo2pDQEE51EYzmiXR58B7n+SHl+vKhuS+RQ2o63iCJg54w6XouXbjpfS5a47Zv+Vd1sIE
NcUKqMU7Mlldq7CWq9AnZSAi8TMqjJ4UM2DAELa5KabfduDEkZVCfPur/5XdPFnAdh+wh7O/JHUC
+tJkDhno5pUer4HP1GSeLjW76PgbX9QH6UcUFD/0w24aRWw+IBTiByZbi758beLFEGhke+0t8Lzt
9xMNADg9Klv6+HKfx3HJUNhAcgmFJFf9KWNbfZwDY5jcbM6jee6GpKoot3lu1U8IcxcPadtO3nW2
tIubUzW5PIdViO1+HnlthIziw421vEo9e7KH3iAPc1AEBAG+zYpF9O3+phmxCQTOQ4OwALMUTvRi
txlj7Ir3fqpQpmVUCtZokqeN9QgLPkn8wXjUailkm//JydBU/nlBFb8S4mhNLCfHI5s/K0R6qdHH
Z+DSInCdYMC/pQBlXxNHwVLDCbt+HyHyyicrovDKa0RtRVnZwPKKw0VkhXgwZ+jdy64cZM2lLDmC
ujG8/7a1e2WELhH78FOXPmjHEmwpX51GmyqLkMPszpgkGOsafuKnvFeymSLypGPHpf+zdokZYa6B
WjMPlxbNIRhB99LsD3/Lip70IaZwIGMe9ir/XcZNFjhOXO7HDGNy3KnsuCy2aB5fFllF6nD6HNWi
2FqEabnvQf2wsVEWGQZUjtp3CKklmCszd3yANBWvXfRY6A5zHmUJblff2Zwg/cesJwCsJet7mjRE
QZa6pQy2QgSH80L99HZtzxH5mo7wPR3TnY6t5jHw2DrlgPoU/8x0ECX6QAqWWo4MADzWsRfSVR/D
4SA+eHTGqM004sVTeTWSlS7q9bWokoblaW9NQNT6pW9lepvzRt5gUOniScEIHLzv4R0Pp/ZRcZ7P
yNwLQ0R6Wkr4oDxXMyzL4DssJlAg14JT4A1EhpXzFWFMo/gOOeVHJKQ4Wr1fDS4+znQKfUlIHYVV
Qf5yubYYhYVH4hyUs0NQGIApWgBpmryIafv6xWzvDoMmuerIAZ+hG6PQyWXVZqRFzgm8bdzVsP6s
GYVnAIfLvyxw2+WwmM9oGbNwPJWIP5n1x9xhMYAhkyDYrtoLfrsRD0e+UylfaIqgIjd4nz5jr2eD
oLROjHdqzs9yb5UgeNIysYZN7llQ8j8m/gUY6qPoJgybsxRUqHL5YJd7tdXRGKVd9j3Yr2ZXs0d9
6aS49nx29PArOqiEQ0ERuuMRMM53SrtDchxwYri4VpRg1LhBruPrHutuwNHXvzThwcbxjSeYTwWT
QhHCg03NsEao3IEUcT0iP3x5pLr7bBShAXEtgUpAVjyydoG3uI7CPNxVjacPZxuUGtJgaPgGn7e+
aw0pIDRGtBBTGQ82Rug7mxiwURmqlYamslQ8ze/yCAi3GIoqWzVm8eOrGrrZBuCFw98+EQEBArAr
Idr0/bk0FC4if5YlFjFmYR3LsnTM+MyJOZAYge96p0Z6/n/k2gG+uOySyH2XeqGy3WxdgEP8q7lf
5JByxqgGsoqKBZU4lhy6IPi7IcIXwoNN2jbKdWGLLw4t5Ymem1BFYeaMtuMBSjlwtdWtrqr7rUbT
Xyi3L1iT+QuM6r/KbVdyTOSIdQfIW08tVox/GsdSYwpfQ16umiN3dSGyjGVFbTS5EWiVjQsUr7xA
3QuXBDibZzhpIQ6+mZRbBrJ+dWIvtXvCB4D4ttAu3Jf/JGcE5gAl7mwpcShqGS8Ntnyjco+wsGUm
6uU2wzHB51poq3Xbqht+g8A32D8l73Gn73ReeJO/mUSU1RndXBpzOoMFuSnijTCOIri7bNu1AiBY
IQd4xWI42GfmHm3at/xTJVvZPNwqDpLUATUBuMVFJBM2ZcqRE7ekg+9Qf44N6XcvFZ5NJGpAsS9z
Y/If2TLnFdW1YFRrF6jg+I5rg8uMy2EKTB9bpxnyziamPFQfo+nYdxbD+3AkylzprYEaG1Dr5AmG
qrkrzpl1qfDyoJ4QgEHDGhABDhC72mXVB43GuHN+WYG8cWQWRbMx98sM5mk/n75FSGEDWP9go9CR
FI19fCg+OMU+DpwNAUaL+7wUz2bXAPoi8lIwYcKHWJxkLWkc8KW9Ep2Kj0Hosq+Xg57Qex1X49f2
CWLRK10zKxyzvKN8W7fcn1NUE1ZeoI6KBWWYe1MxRZ5pWeq99DW4BmKLsw7PO80LJrBrv8g8a1Pe
7T2EOeMs0ubUgweb/HWxnYQv5TZvzRnyffxn8dJKudpXyQc0AtqicroUDC58cwpQNRzYSmXd3AJc
fZ8gpNatRhpEfFtUeuqbXhpMp072wjwzee0D6J4dVfhol2+urlcyEpfLz/IadHAnCMI8XOVpcc9T
Ep+iiS0sfVdLEay7ACzvQBcEzjAL6GceOvEQ6gbkcV5rbGXI+i9vW8iHyIuPYlXkxXD1Q1wIoFP2
Xn0suGH06hbb/Pm/ok2oroK3LXlOcUrPcA60qJw2/jw6kRvXLjE6IVUjYfbMQEE5a9WEwlJPnCe3
LcgwgsWWbE9I+Vu7Go8p/x7/Fo/Tv7qHg/6pU84USNEalfQBnowd8ZvcHoKUWYs8c8mqJgJ4Z6Ae
rKAgFmxmVgok0jB3XTaRFXw1zhIdo//NF1SnrxjsyRs8m3owBljwsdSl+igZTjKydrKgj+ku8Er6
ioghZeF+9vGZH/XFbtIkg2s7vaTydgDd3YCsr1YbPuE61x+XDOUPK5nMEI5Kmp2kzM3JoxqDvpQu
MKMmmAS+8MEELce3Pl6KLroON8C5Hy0qbQo4pVV+yoXXR8nG5AOI6mfMAbzQs9VxRZ+U/kjxm06Q
uJlxEs1r02miNJOJj2uf622Xny+cuiB98n26ttyCuO4omuA+WQtkPV5m3X8MJCp7vSYbdsdqqeuS
nKJS4zx7FGDrgUEcdQqyc2PSgB5B8sjO5lL1gXp+HPuRKyMk9HRDe/s4P/2OeMKEPc+vLj/fGx+7
woJHRTToCwpd/tlyCNF+GMirhhtn1Mo+K977YXpCARcRXYpuizQvOutsxEvreUxgNWvhw+2gvdHD
/isgXCKXrTfm/qOHPt0CEcHUUolt6PKF3e6qFjyRmpuzu1wnofmo/SyLOzEKyymOMMPdBSyp9Lgg
OXDP6ol+H9BljmSUJW/5vCGN3GlXAFFdTJqU4IshuCzDsSVJLcjhj6R/MDoRxqkIDVnpWRgXa19u
ZrX++M27zmXB14JHV9SXUoSvEurVl2MA2QxQuNLWoG8Xr8x0SOGtEz3QTIiTsTXUUsTirXv5kTr2
NmEZAfljZtZnG1BdOUQtMEJ5EN9Y1cnrmjpsd45elp4wMtmNdyHvpz0+8nPihrjQJEd1hL7KP9r+
IA0g5mZsSRQEdzO1kP/gk0IyzOUwNhqCk1vU11xgTm6ekgbJRibhOeVkdBM4k12Jpe9ASVBA35mf
W/FK26I99NtAGqpXu0Jm0M05RO4WiU7VLHMEszoqrB1081asudox3yu1ZY6V3w34yqbIUs8rhVsN
N/QJI0OVThfsstqMoxdLUmn/TWHLPHpMy0jxA/ur2h6Jh//5dPmp0mVGWBy4BeY3S5psUFEwufUS
/8B9emb91rKe6aWXiLMek6/85zG4B6SJ67jHoWbwXp0K+//nUV9BNvNcXozsxpTINR1oMswyxOCy
C47TEw9RypyVkmJEjeEEsTluuWM62hg03R9kMBSj/ug+ghy2pWS41fXxxcXNzAXmwBBjSGoP9X76
UUSGLVkepDREDxJ6wSGh3DBamlzCL3TTarJiDolHwUe11WkqOxQkkyM/P85q6uJ0a8t+iOOWkeCa
GhdUqO73cuqi93F7CqJzOQ3gBg0JlUr2rOsznRq2eyiBx9eR7uZSURpxhzXLjs3d/nvEXBaI0skH
AUjllGOeAopk6J9z7/AwcB1IRZ2L5LpIrmakxmMCSVtUlMia+cdzyG/KC5+H/Gb5qTcqtR4aYKkp
szNsPbMXnO2jDYIjkjL88Zbb7cvy3Wt4y5p7wQwhPrX7MACngJv97AxdqZbtzpbEoVLmJKI2bUKd
M69OsCqSV+m+U7dA7nhEcqklxGF7SkupyTjG0hMp+H+Lii5VFDshE/XcKx3MymdaPuca5nVOusq7
6IDlJt37ZN7EhsMhp9wfHT3rlNEGpNWoewKS7VNsP9xFO/uartjx1Vy54atBEqkc2acdL1flIZ0w
v3jr3qs6agrLpB1DqwBZeTK6rnNZflypA/DOnVZ9JqqolipTgBAcEB3vDAexoiuCdGX5GQkI+O6R
royvFfR2T/Xo/eJHbHbes2P3BpWndZ2oG9lfJp4V9FNCdGyIEQnF+T5bwHcwwV5g7bqGd03hE2lM
xrKLOk+Ft/z+O6OkQzSz6Tzcx0p/XhoByG09ilqlgYS9uVwG41acrqc4PU/kRA70Jr3bMlcY+l92
PB2xyue645Bgs/u3HB5tHa/X7rnuYWjle8JgbQV0kZY4ivoAvyQdGHLh3ZGeYImY+2waruJa5OMS
M2+ZnSd1VpnvpuDD9J9To7GdjPNqV/SQvWlFZ62+XLyIoMqn2al0E8V4KH3GsmI0d/6i/GmuH4XG
IToYM0Uo6a+tYC26Fob8fva644dGaSe1fbVErhdBCT8DkYRErOeNwExgo2p6713LDS9HIbmI5LTv
3uli8T/TRuhWDWqZkqcjsH6XbPKN3+2yWOD7dws/g8JaXywEb4qzvZRRNJ5IeT9A6K6jmCc5KVjI
EhRgCvgc9l0tjs4aSU2RiScw2dzmHrmM17ds69vsT0O2NqbLHdANaPMUH7YaJ11UKvgniLnw4Tbd
dlKE/GsK49q8iR8R4WKxyucckZY0998ZdUZGpxKF+p+UP5reBf3nFiaeoUr4WbODnbuMG/PnwKPU
16fcyKDqdtgVlwuuEe+JbQRBBTi1kS+6O6NJOpedaI4bg//QJLm0a9BK8y7cVGMWg0N4zMpB5jaw
z6UQGjOySJlCKPHnUsedOjP1qFNRb6mFV6siNBdtYwE11rei4H453yZjYQPcvgMOkZMzwYbkkOKS
lG5wf6moJfWBNSDLsfdh+Pe8nxpX2kJR/e4+KraIcGSww3Jy4YLU2Hg2R07jRy6I3ED+Z5Lns9mN
zAUKl9t7GqbGXSBuL+bgwNDw3u3LZgSwLCi1NmIo7uKGSobSe0VcxAiWSIPhMc+X/pBiK8YhIGPI
z3UvH1ct9riPnWmzFnyhs7ZQQye+pOdu/WHk8xaMNx4Jl/pD5VHRpXPgoCh+v0BHza9jYdQ0kYVj
M28rzSQIfcS1tBAUxssHY4j7NIlN0WewgmMx3j8U+Ke9Biij5RTBbtxrgTT12q4kH8DSEcNIrhmI
p/+pnQV5Ioz5u7j3XGwsawrMI35M6BJQtb+w8JkHRAaosXwcZaYMShgUdudUZsEtN0lOIB9zDljD
mUXI9ZopqHwXLm24N6TDIxkxWb3nmBKGdt4qRR7OZqaDlambpH6SsoQRt4JwHOo5bqe4+bxW3JdD
b6c4k1vjQTL15S8VX2n2snsPZSQ7jwvDUGPBB7q/5IPjnVTyoxKQwkD5DYCuYQBcFTgY9G4v4Ei5
Uo3peMH+ZyUtxNnEBI9qNT6fRDbPAMy0a6DPww8EuWXMG1Xg21HOIXCJiRLf40tZO3JQF2eGl4sk
AoqvlxX2hnVvKl2SDdr7aylP4LR5500OQWxnc/ZWPbyiYFCRdBfvFmTSHb/spmlQHwrunuHJSxz8
A1dDlmOV8nrcTIscQuzCpCy5bnscjlqFdv7JJOU0pJixSkUyPmzgngJmb9Xo73W0UYZlmE4qzg21
Ok6GgzXlPc7KzCA4m/J1CJnWwB7rGa4wrfBi6C07Er0/5/AhPaW85l/v7AeKOoWfRaqFEg9TPzzN
hPCIasDf/IX9pg74rwlP0VL0mbmVv87ShdlwVtMeQDLlyyBQZR58xBaU2nbZBR9z2fI/0LjfxI6U
MC57w5sCd5Ys/6sTKx2Xj77RNyjnNOxXOMnSBSzTn3N5P7lM7wa7+4vODJGRJmrlM82u4HOoeWSN
JQPg+rx9BBxfKuUR8OINvwpTToYfjbhWBXG1bTnE8xUxS6FX3yt89lMbfQWKY8UnHxwlxEIE3Dw+
kTT5S1XW8crDC7MVMq2SDr7SAUi4yH1Xz9IC12D2h/qygoIaNprnUaK6Tm8u88mNtgIzYlaxSb77
4bnB/XTbGRajhuvJf/poDNFaIGmmkNsCEMqKFBIouMc8xR/bcctoXAi7pNGMkdkcZD+KWHhI8Kop
FolB9ZTs44uxHqTxQJFuYvxkEM/NyNdil55KeBp0XS6+FRyRhz7wcoS6Ex8j+Qxm+5MeDRFqne3S
u19zCyFTHvZGmaPBjOGITk5iy0k78EDNlJwUJ6T8niVumqirB9K3R8r2xMubZP/Eqm0hyc3h/iRu
/KX3Xv0HFr3Gx5jctrjMZnSJLKE/tGP4A6b+LBDEf0flzJ77/dm94d4inkQIs9idQoPVuONyhE+k
9nuiOLlmxuawlRQU5m2ZyF4hnIsGHzhRZ4kYr381qnXb/S76SZcUmV6gfXjmGzmfk3OyTAJkj/TU
KeM5z7QYwmDwJRLUh0vSaQK+1jb6cjATtakwRk/X1tJmOn+eGihFqJfSKEeBeQ7YpIxiRiKITT8R
eVD+mtq+74GwBvGb85BQ/jw+HeQk0wlQekS77JBd4+0dgZQ1YSAaSkqRBgFcmpBNrVL+aOizUTN+
po1/zFGwEl+x9Df/DVm59x3jw9BGU9WCu4usJMc/PuMKYXc+navrAE9hR/U7fUk0Th16XEhNohXD
JRFc2oU+fRDOPaPzy8nmkZ4fxaD0KBBrRiKltXXcOEF1DDctkYoudLWzJUWtYrfXj+PzM4JWJJM3
6EigUNl97LWWpPad5hDt6SWe29dvQ0zACP9Qt8zt12DfrdD2GEsfHu7WxRm4b/+zQH3QvGTqrSA1
gmtLZymkZ3xqbklapMaYbvIYTPq3p1eGoNSLxAPKC0i33JyaVtwTVT41rzyLJXnRPPBoe2oxTzM8
MmGfVdrk0L3wE4vn49H2tz/okt8Y+8n90bRaeOTFN779n8KhihdOoh98oRGHVJjghgUQh/LuSIJs
95hhU+GU4Ut+Az67aKBx50WhCA6SSOjlhAFbGLUp5GiUUi1F2JyZhs5K3fyMQ44bDHkeZSv+0F3t
7qDSeM9VyqTveuJfx3G3vgtzLuqjM5QHDS+W2KBW9s2bPJPAwH+Q0GrfSbFMlw/PlTCq0d1sgV8Y
WBBbakvb3qTR7h6anhzkjcTiY3stBCyUomkAGd1uD2eRn9zVe2NLV6viFAQ3JGLaAifE8biHIXCi
6iX8n4pdan9hrkzpJID+LzoBX4FUie/4hLKl3wZbGzcTMjk3ZCPNLIe+BrXvR6/6EMeCJGT0RWgA
vuQ/ot0Q9UmQaK3Im9m41bpUrQBT3nzk1zFvOYNx9RykiKKbH2Qssw1G9p4Je8deR28MufQkRunA
Az7lOYRcUSDhnFeaaexSgsWsXBdAWd+x+gFrClxc7lt8S391vstgGauqiYrSA0agddnmSeNF9C1M
rDXNWzLnNaiPhhXh9yUjhYIazLzH48PLTUKP1J9XeFVqUSepXK9xIdF3i7bNg5WXbDMgNKrCyVuG
BvjDf1luLYpsQFXOADgBcN3Mr0e6gFghMu5cAhTzpXberkqToFdUb2uItwJcf1tdLh3fJAYy/amf
sNkQPMk1RIMHRwYrrwKUoV9899VH5HIPUTK7+D1qUs6MBVfnI6U4iblhDXJ35pYqni3zcq5kyTRM
TNdkaS0NNDGGg1LuC6juEP458lrsmsQv02LAtJKoy8jXttf5ktlLQbyYCg90y1bvslTqIpwNsOIU
VkuhC+wGX1AIffADf8fKpcwiLavOQ0Bca+h1OTnmAy+dpDMlsWA8Ne2FgbhQaVKOLlRVov0ceOJj
obMfK9l7Ip5t0fMGlzKNXZHaj0/wFyl/BfKa5B0HNgeZ+Yxdjo+swIIsjyUIoy6PmA79Yq7cUWHb
pO9So8WmqNm89gogC2G3LdsPXy2Pcx+3Eu6+yCET5P5/aD/NRdLY0G1JnjLQQ+F0xMgNlldraNO1
uTmqk+vegOosnEajPmrUOg5aoi06HXnnGeHMN2HdZHCFSX/r6QXHBuW2g2tZPm9ZE/ZtSw01J839
MPsMUC6rrkO8oKrH5k5b/WXoTu1z1WlkZHkyaYA5D/zzPp1oQaCo4SIQtfJJJAPTX9RUshAF9Qxa
e4reeD6uKhR591UQJCdn3kM8j25/h18mTATIFfSowW3dDT48pLgOvnuB+5oHX8GFliuPnsX7vu1+
gmTZm3EoyHmYRC/sne7H0W+oPftNwLfcbOtLGdKvBRHLKwQfspvUiTJb+BbFWn7iZVvEQxDeq7aK
E91BmagQfvBEtFveyIPXyJdFuFDWq1TQpy9wV7qUnUC3M54489ZonBYgaC42ZEyXspJQQBcR7ymU
Gl0mQPpZmqfY2BYMRa45T6DNVOv4cNIjcgWZAWTkhyvSoJxtPGgHALcsmDFjOPTsOZKK7GXoI3t2
k3OZScqztySFV3M6ZG9AoPa5LY24QzEJGFpXOi4O8NMXAgooAOrTReWkZ0/UdxO5puIGBOIdpwl+
527t0uNm2buWyrXTYAbuh8ZI642wljOA/5Sq7nmdLjQqqoCXwKqJIJyIIkzTzgQsDWgZ4DLivFEH
0hap+tCWDls5hESHisei+6GVXG818D5IovtZRAv9HkjF8I7TFVgJhGNdpN0M/CmDaM4J338dqR49
BZ0np+pB8gjYP5NluMA8HLNs1aStqP/6kssTwIHSLqWFrQSu6matFnk+W+YZxrNEQ246GRzHsUuH
Jz6bsz9EG88XOrUS4c64K4NwO9HlcWaiYCqlDoJPZRJw4+puYXn8K5ou1vdtkiTkdI50CadT7RTp
5UgxLVcRqZ5QSqJYMRHNDwn1dLhaZc5FkVZcDQjt+ZAKT3O4OSGT3vPrz2PZTc2iSLsjITAQjq7q
RbB5m7+rPGjAXBhR43HU0M0qDBL2ogcYl51+C7oFtsU33AKJgg6mb3F3eh1RV6u/21k1oHXIp/pg
SA76Qg49kV7kI23PY8YW+1LUz5z2sJT+tukn4thPoevRwX2jtr6LUBLEWXISgtEW9AlcsEbjQyOk
RyYahXtMYldQVDDnP4gNbPSssHoKnGnfnkdXyJb8B59pX0Na2Li8PwTzDzE38WqHwTH1V1t6fUGB
dxPDUd7pjSU/FsrlmD7Tq5XXpvl3/yc6OO4RKSpB+Xmj6h0iXt+jfVQRhHevUy9qYD53I5BVv4WV
JXFsDjoMlvuzOkhhthMv0/eAyCFXoMiKQkRA+xxcV9yU1GjrwWX+JcDt/SibyHhHuxoaO5UQO8Rd
HsvntnKamceMioV8J/BGa4f363qN/9b7Ucc/+/hfjasqUIt2WoVZcBXMlQP2tWNiHa9MY0ndAAi0
zsPBfOtEtrXBz8lvfmX3BsIt4lW+4QX9YEJyfh4Z+o6JxQR09u2hi8PGYv4K/ftSex/iTdPUsm/c
3KA7Y12qVG2Qg1mvu7RvEySoAiBms4T2YvhOwrgA5pK7znMpZs/kf/RoSZAxd9ya/zPbDSNjqU7q
liP4CClGoEsy6PgYq10Im02+QRyj/0iiSXxrrqcl/KHCMA3DzL4Xoj1S2rcA8KNyXtSee858ISk7
cYz4keTzAiw0SpZZrk0dJrV8GQUfYew7zqNucpaRjqI/tY8hNxGSntGd+WHPVVoYmx6CJ3joVkKD
K3RwcOSYymBuUowqSgp4mxvpZVLtaFKvqFQ06oJtfymne7lxegT3FZIq23nsFym8HqfresJ+tfNS
Og5b6PlpPGpSjobwhq7NQMEhFr0o7qlBDim7ZmxJipAxFu+kMjPopDolxa7iCONAALK0d7KAtknG
ABUW1MFa1EcrtRBWbB/533KBqR9MeMSO4++wWXYh1+wMLCcBveOael+hfHVj1xy3W9PPMFdAbhM9
EvnF+hBVZJdKXuiFVbmcNlKV7pp+hXU2I6Ce4c4lXeYjEXJB0yxUHMz/ZK4eKNH+bIcEIpHyoIEV
ve24A8COOADnmD/htURjgaUq9+h4SNE+zoGG4aC8pX+EkHaONS76ea6RZBwQ3fkxiGa+62oXruWf
G0724grypArKpr6ZMUEMqp8p02fTrnXpBqDygX1MkvXnjQm26Pv7c02UD/D/UglWOPhcpbWM9gib
MBy3gQTYlvCqX+OEAZLDlM86fPckhocc2Ov6MhOmu+coUm2qC9r2FKGzO4TO/wWgobm//QYhGzu2
7KjUwEMPvIfzywgQpqFSMuHN3D2Bm17QisenT5ltFPbhUtrBZ18QAfNj8bgEfmH7JUw5CE2Vu5YO
qX+TEngEvg7Qa1U7gcKaElDmX60WjP+2X0BjQzPzwEsXDEXxXUtItZJ19TMesU6uO8Mhq+8fmqR5
E/u0LxktVdq+SAWP6Zm5qMBfk3zOyNNtS9x4ATD6gu/l8lkrHb/3qYxyy/jndcQT4U54814Ch+nX
HKeuHG9fdvb4aSwuMCAP90lPeXofjALJPZ49m+11g6q5d790N8r7JZtGO3l/uJn9QEcZG8f8hUyZ
0uP8aDma8Kitqgrm1oLKrjj8lNiNpPuOw3PVX1p9qqah0/mLZvJKaMk0fli5OMnJk+VTOAq8jiQU
m/XzMre3N6mBvHHzO1kTAhEnO5DQzbzeQy373YRpI2MA+XAWA8NNJxCbsEwSfOILglsoKfs6n/fH
2nKbGW+dmD1aIE2or1bZPQELOlz3E8Af1kehjFn+/c19hbO2kGoTBG987qCiaJFD2utcd2NYzzxj
/ZHH1m+f2y+3Degk56/clai0XmNHXTxlrLqWtx5Wp++v11fvy+ZlCWXwlJQdTvB7Z0cQyBpJvt1P
gc/eBH4q0Uj8SPpV5OMIfQVbknWg0lK3TPToAvvJs+DSZaVpgoH6c0q+Pv9fhAbj4AJ8QKLCtufk
Ghdw0z2F1KhGFPV3QO/DhOoVycSkJ/F0dRjk0NMiXL58OAbTgYJf+0OsTcL0IQ6z4n6rULTqVZMI
jVSzmVEpTttzsCP6BCdf3I/LI5hfzGWd/55A+PKltsdh+aqJ4DBYDe073fDDb2sksQM3qH/T/LOb
K48i+WqULTA4KtJ6dEUNPiaOHxxaCJVEhgN3LRLb7FiVaB3DqcNZkRv8zYpZk/T1xPiyPZSmV+gs
tELCeHoRyrbmV0c3DzKw67pvFhXq7JaSwG8TUKAZZQFlSg9fIA4Yc1FLn0cvfNi7VCZKZ0U+j2us
1+svZX89KOK4SsvLYVThddVqzCcbLQsIfj/blT8KSgu9tOPMIKoiMj3NITVciRsNKrNl9mwJok6n
Ee6SfZmW49qo6riVYetxsikwTABqLJag99N24oak7Qb3d2XD5BncX+QOa7bowwyYAt99rTVmNaO2
wOz4ptuKXftgMs+x12egPvmEhtaXKuEKlwoO0rmwgGeukRk4l1uRYQHQ1z1x/w/xQmQxj10Ydn2N
zYd/ocflpAGR/LqdqRH4t1nWnBjxbZpdj1sAHSEfq0LXdD0rzt7awLgh0FTPm9tvjda0QtXBb5IM
rweEL2xoMe7bn76dfSCabIfXqbK5xHdfIO67zhmINsNQo7KjSzpMwmXoZQGW7gam8IFW3o4SVf/b
ccnuvRIW55XfK7wf3mAhh81mlOO+Ses2HpgfHaybB2VooiRCc+mcGbjLHFHzcqSgiIAH+pAYnix0
WfVaz8TLbca4I27Q00BuAGfvYozbwe/nSFnMq4gqQy5oLqXBm+KNO33zFzA1hN6Q1EEaRiFzrSVr
Mh1K/8CWyu68W6unQu45RvkamMgEGBXk5WLBTjFJiiF0UlbC3WOVWgSQAVTEiL+xzteNWPtEfNua
Ulv1JXZEKGySuIxOqPni4vdbdjYH2vH6QGyJZ/rWOjbnsrEHEwAorpLssC4GrcHO65U95AxxX005
QViE7wvyfIHhbS6ucK0UuzOwZv/OjIFsujZOzNvw7/8CGZX5xOW6DyRF0kH8ExYia2TjX9ThpaFA
5aKcXnnEKYy3ySbtPD/gpukFqUn7IVpC+xyVGgx9IFi0uv4WWmuMNUBNgioRo04apovf5SE+YhRT
NZiZ/WtpmZ9KfL2qrYXcdQcq+prllFQm1GFRcN1AAPF2ch0YVT0q6nWZKp+93p0LVeJHES+eXHhL
4NIiTxx7ShmNmDkQTuz6HKpyxttfDwCQ9tgSxUDMWtxrQjsENI+Vv9QUyk8HnqSwNj+/Z12uiEz5
sA63MJ2IwiBvrAZJzZeT75j7Qsi41GCNxAN7thJRvwlYreDF2tZApBvWHAE9qcrvQDzQzYYICEwh
AQYV4zarA8YK8BnvfESZatIc2UBZceJ1laXZaSO38VE9uNHBP7WwNryeSAxu2Xh6sBWpB17s5T+n
JthVxMXXIZhK1LQeusSVKejVAI0mtkjO7ziIizAOu+xiuG/b4jrBKHjpfdXFhJtin3rSJfqOMNji
vXm+iBehz3ZUHtP/2Qo/TMTJLodez6k1oOHYoZQ9H/UBwP24NSxdpi6xIVkvm9SoaSS+AjwIt/ex
xv/JDLcpXiiE8O99b2OYpQEFMpJNfUe/lWwt5oV2NcG820ApSfq0KwcmE/tA9GVj3ZvEid1VR03+
tsGItoRSL32rTFo8qR/u1qpdNkaCxVQ3d3LjlZ+JUtskkGSt3sInZBbT8qM7Pw3IyCg1tMQs0+Gf
gs06PQgXWPNrzIh7kgjavHxiOMHFzXSndGeERnB2GOdA1BE6PieFbLOnFJf/k/Iw7PNgc8eAgLHU
NTtTODqSq3uOxpDQkMWxshBZQ0MKwgEfu3uDGuhOs2HUAANGQEgrIpMRhs0iMZ7XeAE96/n+OifK
yHoe6fslhajyRFZk6+0ggc4IA5HdH2AFoC+S8rG03Br9SCzSp1kJfr9K5jH3td70xZmG0oUOYrVt
g78mS7kyY9m5T+GPFYIz0lgffsBL1Co6ys4NreuUZz8nEldhxhd6KhGf/OL8lO68MsmxWV6Sorc3
rMvqkZ83DNK+2bDvSVa+vW1qJlzo4sgQeX7YcPIJiWEv3fmtGmc3DCOs9cUPlGm9KVQ4AVzOO5Zt
4arQlJBSZOYO3Zz3fUg/JNy02NKXnaVc0POrBE3KN0GSLQrLCLspWxHgCmJhgMyUizyfDcRM/0Xf
kPl4Am/HY248H2Tkh/P5QfIfZuLfqgHzKTBICV2TJZDHvC6aEdtcrFkJWSJ2/CAjRTxkWFddqva/
YboKmbCs1qCSJEvuw0BekbK7hkHifinppTF2FCIjr5UKc5SaDN+CkUBSxZQyov9eIPOZmO2SLBIh
V/bfjXPKZftCe5KU1m/dVGkmnQOId+xxrakxFGWIPmmgW54Bn6s2sLu8MXwi1R4+rWxpGV9jjAit
CLhhMwu5MPzhTxZ7Tyr11Gw4oKqle4e8fwvEgcls0RTcn/WJRrfLNp4iWdFq2c2QQPxY/bSlXCsf
RFxJgxC4CZDg2HPhst3c8n+458Ua1vnlIqWyV1sBwn93OpfWcuRiPtpU3qvWZ2jr0vZQ5cBqF4qK
9Q9rwFCllFx1ROe/Q168tN6riy9yVQYm4xIJJIKhV5viA7Y26GhgXJbW2ymrlGV/RcuLy1XJEdU+
tUxfVdyuuVgYf5yDVy6YJOOqWwwpuQ8GJNYrCK7+xc381msAwKPk66R4qxpU6Izg0GZdjSuw06oJ
eBcBlHKkU61kK8ro/uhZWKx63i8Z9OY9VjzTsIK3oUDIqjMt3wQYQohL7ni8BPgXqo7O2/UEQUSm
I3DEOt6UxvJf/3n63gNXupR55RGOrkVrDIERNVl3jT//sU2vA5/A6/gyfZ2l2CtgaBNwyzEx859Q
kFvMDYHXOLm47B5edEKFw2X51fbGAXB8dYD9hYMa2l/sWR00lO0aLwsdsQKGj8E52eOV42jicZVO
N/yroXsF23sbMbPZSlmvD+cPuzJs9hsyCiPZTF4A8oT/yTwbmNC9WP8i1d5332+2BhrJI+7ORBl+
EuOFGamGTH85v9LT60/hn5lixzLnMXE9Cuu3/jyES5LNbWyO6tdu9GYloRv3XJuS8M0nrwvpK21T
3rpIHIQ4hozLcYrfBxJWpz8LdwO3/2tqBaSvRuFt+hS65JE8y7dzCRBFCKJ4HPRrAUdPMAApaGcG
OTUKyXM27obh/+u0w8UrAo/3UE3vowdqwWElBeVoYM+8B0upSxUyelUHpY3nNKZphT9Gx6ntDSCp
CgL5v4pjoYNW4mKi7NLPbJvuYQtaQRB69qgmJvcvF/Z6QfmVFZNiOZsqi3VoF2WanbtaoW0TtK2Z
cI8rIYdXh+WfWzZWBlKQjBB4j0jOV2Eyc0+ypFxOruTa/GZdeFq6i6C7bl/Y+nNHNiFUYiMMtAEu
A16UXp+oCqE4G+aholgW4fZm5fKD2rWvdvxgSSQVwLkD+umlFqzgwbuV41vZKQGxgrhHG/GQGJVS
0DUS54zMUsYOwAvx1xW0dgelWJXQqifakdjNpXqcHkF9BF/178vIgz/4pcadp3o6Vx8ZCGZzEg/J
hF0Y8Ytoxln0ZrmnsZ6fF+lbRl/WpUWREQ5jFN5fN1o02GDZ2k2UKDC7scbU3UIR3qFXEATPXsKE
9FWCUM+4FCTWiGCW2+bF6aNtLMp3yaQIFDK3wBDf8l3IgdNjfX0+8UVsviIP6TMVXvvH0rrAEzQz
VtHnUZW7gCthWg5I9hT8BBt4z1usZu59A18cp5lqTkqVUek5K4npr1mcD2RvZsQi5nrF+8bognu/
4teqiSRYYF4hvizlXZ1NAB4HhK9kBD+v2z7RBSikfurHOXVZd2h0kNW1XeUH0Lv2ONMLLCDa5Vdt
GYwR70qROWYTWiKxVhTmrOw+aejrZYWyrR6fd8pq0ER46KMitdEwrYqHzc0f2eIswQ+XusRdiXn6
q/zH79nOwcRD0lwoQ/GdAnm7T0pcWEwDDQf8RYb8PQfdrlCp7sJzUFMzq8MJ6/6bSbKXVmSoQixx
0JypnwRiufkzjlY85138xaZw05n7cM7jfDaj/x6Co+ftyurg6L3JUSxcPOL8h2FEJt/yNABniQlt
C33BeNfayRyGEocUICM+tbPPHRjBzAoaozHptBfRtw6tdbiNP0k7DTQYmyt1cmfn2qFRHcoPO9vs
JQe4hlqpchOg3tw6NEBAFBY06aZoLomjCmlceTD29l+3IciJKs6mQFNQrWfI9+RrHHDJm/CBdnsA
yVizKKSrfDl/w1UHkbjdhb6saoRsTEZg0f+nEKf+WmevCkEythBVY0m+JnYaFmZ/VKd1ki/I6JQU
mRYE5X6Z6DE4b2ZRgBWthubZ7vrx0pB6KnKVfGELjVEarkCexS4hJgsNpDdeiFEYXffFKegsYH1m
qb+oNzO64A2XEZCHsc7ckLv07Qd1lfKZMSuOHapDGFvZNsmBdjZarszaVuk5GRexGgWCVk3XXuvY
qLAlbN96zjelHH1DKNqNrPId+D9IyqRr4ePPyBh2LWC427gr48+A2psgwOwldybS/Tb5TWN6O8e1
umpQDKvbk0JhsTNFz/S6MQeRdx2HcCVCh0dBv/wyGMOBoUL3NNbAdHTNQcg0PNxj4fQ2qy3fmLyd
X5kpQyaDOYqh5tt4b3k0OMO+g2YuLuxLVO/+MzmHa0YlQypwr8aq3eo0+bhigdipvmEy03URHx0B
rxtKSU+e/jO5IuVTAaqdVVziGQAqguBnjCHaw4eoGmx2Jc86dKMKTiEwJb2H6oG8ENV01HA28xxy
K1OyxmFEeBbUJMW7klEUM16Eez0IF5us6i6owENe5z/EGwxQXvWwAJgv0r0aVORriqkpraRY1CQl
+guF++TmYTH0V9QJqHcoHEZLqqiLykWUVdfS+9yRJQBmcGv9lxxqejA9ZKwYnSytriV/H7Bc3hII
ujN8nW89vb3QfxYcMeWEPxEfqpC24ea1DvCBC8dr93AQg/H/elREL6vpIagAjges0IL0HtzshLI1
SpU2ed6ZoZxKB2munSavScqrPtw0NN2iGxhD1n1nJ7B/8OJxG8JLwe/jNKUh9w+kzMWVhJTVEGYY
yVe2e/ripBc5L+KVUabDN6NpEIxggIBvbWLdx/l8Mx5kTaKMfILZEjFPJFVSuP2jQRHQFkTDY9Cf
+sfKNq3Ftp5Cjcg7qj4QBzegE8oMP1/7/nFfqewzXAw4D9ZgZwuH/TXpavCzeSxWEjOhanzd2xYW
W+fe7yZNfo8CjtKjynve1IyzVngKC/Tg4M2h/FRkO7g3G/OsRIZ9/9xxUeGI0RFaXOZjUaBmvCS1
sNJhLLPL4Iqaz3+ldZ8N/RtWcCBr7ryDYfO4f/vq556WqmPLVKAFIGrm5EO7WgyZomUv8m84BrZ+
qlEaXwhR/ROe0pcYwAnGr3Ef3aw2PN6N0ndFek8+UYNv+ueihYKGh+ic2LS4lKgk5bOHGuJoc0z7
1zmugN4GGve1CbyDhQA5uA4Z7tcv8R1JAREeByc6/hJ4ywIHmCc4PWyYyqnlwUtv4WFlOa5tgMzt
bFuoqmJr6Uiu8wPYHDNhI/cYfQ+uX4B9qhakI+5gehVi2JUr+leMAfvkxj8SVRwUgnvBGT+8XRCC
A5aJZO0/nZTmYkKmUvHFBrT0edb9QYIHFLKlz4gyamCj65QDvde9CHd9Luev11tY+IEeNvv3CWYI
o1tBBZTpfyf0BcRAjkPCtMXckvBcTCesYa0OBfVeu/cMkYT+EcjDYM+kYzRDvuHieuzlOz+d3Qd9
6KgXOL4of5yKp9x3jQwfSd7lfR5DDCkpw7btHzqnOl2c4SvqS5KTDByJ4mRUqO9hpSy8sI3HDWn3
n5btbHiJhXbDz9c3Ly59r8WWMFyO8i6vzM/tbbk9bccEluN8J5qrTVfCPFdhbmIweS1TXRuN3yyP
OFfv5iISoResgQfZ8/AOnDfNzHB47YOJ7Wbon1oogk0sHwBIxEullhNGcMLobMQhkYA33HoSQ2ta
d+Ff2sN9bhw0SDZG9q+lhL16A7TsvIfpxAbm6w/3S7G3UPhU+sihSG+dwTh7zy0/6rTgFGErFGKJ
hYCryhh9X17cY8qBmzIgCN8bwoUSBCemXhmsdh+HYlkBTjQy0MBRqBPHXJah8ZKHb5SsaI3f+SPC
buXQl2UkTaDWjSwb9DGRByliJ3iNKqSLOMtYqnxlonYYqQ4zfcRhmEZ70iYarr6FvabHNynJZg7c
0y3Xcfz+y4mUp+d3Efztiaka5m78oZI9X++ZiK5OEi+eCSd2Unc7yeat9b4EQQNbLGFVg6SgTxSB
hFguDDN0AgTVj9P+2HiIl05MhBwqOTnLMLRbxmTSCrkxmh7qWbIZuqpSD//h62SirW4EcNVhobSC
WEhcd8f1BelinbFuxD0V84VbuXFJMK1R1TmGbfcb5P4UtHjjX2vy0rBb6ZhKACcouXYZI14Dphjb
NHXif+s0nOf+YwBKFFJYO5ehO2VW289PDk7iOklNn7FCFE7qT73R32f+hZxr+a7o1XW2M+hT/kwY
ZQRarhkHfWd5Wxhbofu734i50t6D8eLrqumerBBY3Gna4yz/Wh8Rp/EXSUPSScAXwpsHIkj3mAu8
beaL5ykvrJRqF/jeVvDdewa9qeFXp5rv+RbWKg3q/QjCNlsbZVVJ/jXl1oTRn8dyeIJNZb3DBA5Z
aDepYMPKcPK3HuZJEWSl+K1wQBFYzzMDD/LOWx0wu0wZ1Qu7Ah+YxCTSaGnuz0xuMbGRevaDtfG5
g29mxQD1EgA3/lAhk8f+afnieXTN3M9Ox+HmV3oimhwo3VVlY50+RMhZP0s1Y6xufRJY1HDzBPdX
mXEPAZaOUMHm9YassjlV2o2D/3FpV61vaIvog+sJxV86m9iz5ZZnaaL4Ujy2gPEL5ojiak2xK1qw
si0aQlt9kc+dIsi5NvLb7sMRyA+jvyMfTL9v+l66ZGe+XRg3O0A0bGWaIGEWHSJY7DY8NnUUTSi+
xeXOCeHG12LhHynnd/VUHeqMsuisRTh31L8eaEX3n7PW8V5v5Z+peTCYFtD1CPjuDIqMlkMvZllo
N1rFDIO6BKUPXjzWyL0iSQeHpYJpnLn3AJEJPtgE5QyASEKGLiqKCQB1JsvXtarDdyKoIyHBEFuf
+Ur6YNOzmC50KQfhAkC/5TXHuy5Nw416t8jXTerbUSVD3/5jEbIqY5/AfyUj2uorgd0PdBu6+vHn
mRYPMZAsTdn8VkU+Kqesyc64CcjCIaNZGeU3e0H1M+7wbtSNUKT3oGj+y+xB9zrTnb5NqPTEkw5K
AmY8NBgHSxgJFYVKQvBBcPZlQ4wuuCUb4bP2BHxNS5bdQai3mBbTYwHrFagZFF/PhjwjDF4eTkCU
38YU6THZM/dy+YZlCKJ85ng8JKrTS/IfKI0cfyT3BcuDCRp8dC0B5qfwhF2xzqsGowa/AUF0BSXh
WL84xzyOAO5NriekA1hqyalsQssKSjueeSxqKPgyudvkHQsDE58pMflTe1Mh66NKqNi5zQA4ohrC
Smp406tWaYO4AF7KbP1O/GdtVQjkctBPXv6Idb32dsMS/TkSGZUKppMjbw+5EyFr9s/edaMEcMCy
cchD3QK6DGkM2+ledVcSev9X2SIfa2U3V0w8Rmo+eNEKsV+xVSfRlisFcubBrHqusGtspuzYZLRC
9XEctBOBGMKKDY0IueOwzs99Vh47gy2JPDyclYo7kxTftv+azlVrwJmXDQcKR85eE+/cD/BeHSlD
jKPXbh8+7Uf7A/cud2DnIJ6Iu0D14G9UHfGBbMyfwYfM+zkW84DXVDIso5n25wP/J+GeRiUGdY9V
P2iGyIVv0A3Q6U6OtKEIHwu6tr5ljJGNal1eyRFbiWthgC+Guty9d/D8ajgay/wh+1eQSQN6uwdM
452UsDOERCEI8HUTPZeOVeXx3ZnwZmcJ4e57OeAOuFjwx6jb5lymX6fYxDQa1nnmy+tafftGsdNt
ajUeEjlKn7sEhSBRMwE/FLflGzVsHJkhg2wCfDechih6pCxeG7kFsl2WErGJIAJgI741Ufuz80w1
PAvNPlFslT3ougScO9ZbYRRL/xOFHvHp461X5IgEO6iTDVeBYfihdTkHkisW+V717DZsDrVpQ0p+
gDV0Jm1QqonaY5T+zhyM7LEVgw8iOOTI+diZOXYIKd2NdS4Rm6id8rmp2TwNA35ACmUm02bWtFCd
QTYOBcX52ubw0ok4M3dzXGjfz0PNQK+Myg0ksfXVURDpXxJU4H1A/ulznyk1FZ4MOvRAICEPh/9n
EIm4SQ5Dkhjl/tSN79wS3Ceyq4FplqKJ0YazrF6ENjUwdKWIe07eS19Y5Aba7NQt+gxFU3cvYtrt
RTzdaFzsL04Az8BSlGqatNJGd4IPXpZO+kGSyhn7c3F3WrONFoMv+ARwjWvnQ8MynXROvc6AIIPc
Wgh/vMat/nSsTA8wovOkO+cUljiYuYNuBn5+rFUmLatduhK5jDwe85sjJcVTpWO9dWlcrUHRRpyU
ATnstgyXdq7tfPxbArp5ynlKI0P+HOCInAOcSJwc7reSvg/+xK+GGfQeDnuLi+IayvVCejvNAtWk
DY1mvO369vj/2MupcbmRjIxSmw5FgiPU5p1Tk/42K//ZI+D0ZGj6zv4oBB8vdCCZkn8OUDSjI3nl
9KBHr1ZvvQ48DAxbcyI9UvgwNqxHgef3kuXJwxMV5IcTW/a0W/BYx47giaYhK4BfvgYzoI8GBe+Q
Itm1STEGw+uBBPM7zZ/aMGWpLHZ5mVlbfQphgrCbkuEonBuouxuEnEpp6bfDbxK10cTXzCi0Lx3+
OwrpnZCBhHDAtconh5RKRhlkhopuDoF/OpXgtCMhfaH/SzOlmwCzLPaI0Hsc5lfbU2ZaDtTtPCEG
Kg4AiEyASY6Ou1LJ97lSSVDI2L2o4g56v1/sd+5UncjRAUqJnGjxpEyqL8qYd+mjHBg1suSwHzAJ
ID6dfltB0BsVnbs9jkC3opmPiA7UCY9pmezr2I4Zhb59+zeEgNvPHTqsxV6KP4c44/Vzflf1jo05
KR7KQQQES3r+l93ZjTLpQuMihVOrDiQukReHvupZcyKnPGI3t35qAZet5gfC1KpIlga7ug+2ZS2t
Y9tbjHd3Yk0vcx/vxXm9zOxUtTyIWlHLmqgeWy06oiiywDxhIpLVA1Nol30jb6myiLffLzn73Bml
wGPcsIMxLm2SiHxDLabM1fPasjlybkqbYLmew3TjoJaWSaBMlzw9gYuGfzzJDILpGIt8dQUrtsT4
9Zm9UAWS9kpBbek8R4siqG/6UHeLL5Fe2TN9Ky96DIVKF03VaAHbo3RiLlTSaudfGgqASFPiZ14Z
S9BEfiT2PIdvkpdR4nFASxJmwzTLOv86SEGuiwgdZrkyb3qCSP1Jv5eyCZwP/rLX+wHfPVg7z1Rg
lKmi8dSlIlEKqHy86xkTenFvAIqMvvnY7qc8v73Ha8b8Zql9QOFQp7JuuTw/MawwDvwLAEZ7BhMD
kqFa/yepkE9o6QZSqBYsYWtDQtnmijHAGvioN1z3BgP+6bnk8KcCaie67bkGxAJ0+UGAxIPT9h9N
E0YK/Vnio1lXJD+la02u7tkl+ipywJVhSbxy6u3QWiM4Ui690HGSEa5fSi5UaMEyWIzjJ4mZWSVM
9jeU7MPvCxjeixtcul/APr+Fua5hE7IANiV4uhRHoJeRRQwz+epc/Q/nmXHqHAnAQTaRDwJcq4CH
7oUQeOWNw+8IXGSstiNfLuwJfqbA0c/32j4rpkGsLZbfvM/Zni0Oy/wqQLFE2/a8kfKYXfZlNysT
LeyV6fvdniFrCxnduH3/qriIFl4UCi2JVsNkHgXjxJ/XAJN0YHrB352ftUhBaCr1ISpAn79mWQ0h
SqygU8wp/pGHC9Tk7LaljV3f5CECbMx6ylCwKQPy8TGxn0bMywkR7yEEtCt7uY5nZo4Of9lA6Bq6
uj5FRJL1qZQRSQ6W5GLTPhYGMlkyb2dtKRFAXU7TCnKBBErsLLPD3FEVTVeMe24qkDB5b5BIAuI/
I0INFxZlLx41oCwBWpOL9Ct1NW6jPRyi6Uc6c/D+sUZ07j2++8jgiwrTfRUyFbwtvpXbnJ+ELKjY
1lFxycK3O6dLRcLr75/8TYPKEFuxByqQShkPfXwxkmaaBpvNuUYahBKkAZHdeh3uGNz0gkN9K7G2
GI5Lx16pldOeN319hMttcS714d9vQ9m2q6Mrxi4fziP9cddPK3GKVYw/7UKOQnvJNYAdGPT5rGph
L49T1Mlqt7ayUfTwdwf9UvUI2o9sP3kL+NgyxQXc5tP0MGhRgDJY258VQTqviOHd1N3GgHy6runU
14DzXRfuh3fEmgU1I5LMgo7WbxDKX75oad7mOfmCrc4ojAclqHkn2T35DgkBwYcNbWYXFNwjRmH4
5bXM6VJhXlxViddPAEwJ7Mxz0ax0IoMods6b4KPBgm/0a/RqOdbcbAlxk5/2ZUoLYrG+AcdC3Z6L
GqvogApFRF5RK1N0UE7zNLjXRGEk7zHTQEyikLIrT7Y23kOSmcmyHom+BwbHW20cOVPMhmXaXqS9
4oZQQFw2uyUaXHer8V/B8Dz4hg7O6uJ4TlT4MzH4j0WOS6B7/LjUDzdXuCgNwF4BXrfeBnGJjmup
fvNSASAEU/Vw1rI2osR6c4xCD3/DgIyE+jmCpKDYDTCmz8DwXjp8tOIJs0VSgX/TJZrGW5OROc62
rgNwsDBGOEMsDqjAc+3wM3qywV08YFje/IywxGuP7MJkgBnP+9Lwa6YFvEyDuRxS6j/KJkWnxwtp
6KNWmSEuD/wZPUd75NBSPtkD3cOPkw3NhzQwKblm55dSI+SdNTrFQNTdNeomTJ4iKFFs3jIVG+Q+
UGIrASAz1DBCs8/+1cV41fnry2bF4n/Qk17H1Ld2wt9HJoLCN+nwfC5lbAvTpqfqeELzXc7FZH6A
kLrk0cbyt2J9a2QzSE3LDf3DznU2zcSxCzQn7pwTiPGiDVaBXHMxB5/kblPIP1hhUQL7jk74rm42
JDy3xvmXpbJaDkQ9Vut4fGbWqVRK2+S6dcjhmcTiuDBiBpL5MdaycBwyEY3ffmTzr8I3pdY18+j8
RcgoJPnjWPrD5cs/QcRiqZ+AbhVKD1vC7nYqeK/fFu8GqbMfqXTOMnIGdkI42OkB8WTOBC111H9r
E4dFZKkP3TMIdQIWo8/nlQiywfTJW+idu9uxDcCBK+/p80X8LT2pKgfWS5yGoqftln4mwRmfzfg9
uKPSXxoCvqUVi9HphC6+IVQ/Bg+s/J0u3aZ1iKC/Z+Ro1LtUKtv4LFfHnca6NJTCra5GGLMYghmX
3sytKdglneQf8kjb9AZohV63MxXH4vXrQ8n4VoBdHSWU+3Evblgtbg1/Hcnc8U9U/ZT0mgSnDFVS
TrhKy8bDJqlaPkUHHtsXGYOQGkMx6fFxLBqOpKPMFbUnfUhwtN9zgJmr8GM+X3Xlc7nEHjyf02oP
LJ03CvvJN93OwddEZ61eEObjpni/U09p7hzz/w8JFg2J1sBcfWTk3Ynn8fnRXpd57ZTJ0bM+2LPB
Y/4f9MJYhyyAIw3S2R2eK/t/ENFoZ/yp9z3IEp08Bx5DUxBKnVSuUHhPQaHDw77zy7qlsX4hRKy6
Y6MGbextW6977qdmiG5abYrUkO6AFwOd062d++3X9nZzEFQ6tRr5Tpz56oOVY+dv0A8s0/RJcC19
uMjPSuD0jQ8jxlJ43OD7cyZlETlTTiGBir7MuVLKK3B/APynaSFeqtLPxxbFFivVr0xCivis7Qps
0Y9sCaJS9FyUGq1r04L2C9fZhilvwBZyJHq00otmek0OU214mu9+dpUUNdYPE+HFpgvHDSIvptcM
K9YIGFRqfBWsPAAdDSl2W79uj/ySYn/0569wmc5RdQUSS5CtroRdJZJQRgiUxnLdiSxju9Pzo1t2
wpgQWkhlSnS2balrZuhtADrxlin264z0X8hQLXJ3uS0bvNut3pVdcMgJQVtzU8FLL4LMm5LED/13
kG3r1WBj4ttI7ukSNJltcV/SBL8wk25RxyWkzCai+FG1Pg6Yq3sWbvGWWJhfxueyZOwEhSgyhqIi
rLLKAZFi9LYdVs7xNRYV7bLuAiJ9S+YMf3qN6kz8LatkVsxD7+KePJwOKbdJvzMbIyH7RvleXXD/
F2aHhYJWSePIuHf/1ynWB0REIx8U+fVfPhNNQUGequpbQ3KLcqZors7MmmYc2mpODMpp/y3wqpJL
pZe4bzahHUuhZLZw2MsgskuTYfiX3SFhxN7YTWnLntse6zs41IkIL2yPnczBPhGLbfoNKBXGcr49
TCbHlIzcR/WH/bVfUyPbnARFZ/9XN1c6pon2eIEKINnFYytgj4JY/wwF0AGHNnu7EWfWZmH/AYJB
OiAcDGQNy48kB/jFQelRDHZCcrkujJhGyUNsHuXomN8LzqCTuA6/arip2OjfhD2Zmh3IWgE9zumj
Jl3oli2HezH+uz3I+glHvMqn4WmC4M6O+VOLIP1Y1k82D6pSvz5ZkcWevaDMfWUYBp+bBZ6P3Aw2
IFPeNwGfuQxxRJ0CRcoVsAc2XjhklJXPz9a2Jlcwq1RZ4pIal7pqro2x7qCc7QFy0AEanDNUfsm+
N3YwcMHiepVioEEPdqESLdto0+YJPwWg4Mn93K5hKES97QbKIm2MnlqjnpVGxkCoFX/zvmQs2DTa
5h27ZPXBGNiwm8w4RmcWnuNQ8Gd1Vm0nqVU4GoxDOmGT7g7xH9crKBF7LroI8HVzFWwT/7o9r1Sd
nfRjEvZz5pBduX+T79vsOWmOJDQtj8YwHiF7bs0UgMVbbTy4pyFc9Bwkpm+ayeX2iOacps6fCuZn
KIdvtjHUY8UqhuVzKQ/lQXNN2Bq3EMC4RhKHojgGh5NuneE95ANaZsgCYXpHKHfMMQhEwCJYU2Kf
16qEb1y2eMdiZuKzO7Uebzk4QMfHLVsb+sJAoe+HubwZNrk6Zd+aiezwc5ftMeE4rsfL+I9pI2I+
RoWyj1op6SVtw36jTMq6xxcaZPeFf5oyMUxslb8SbaH90W0eHva1a5qi1JDqg0ggSWJeaIuELVRI
xa9/cKrzMZSqRCfxCey2eEi2tvYD5f+th2zwQR3D+ysJFay65RtfV+0qlmyuW2RL66UwAda0HzR9
Xps5X3wnbTn8soD3mlppxOWdoM07GBBgBetQP+tE4jW8oD2K+K50J+DS8UJ6pncb8DjXAXFKW8YR
cJTqgpTvejWxqM0zwEuqC8+xsuMqeG6EE7ad/aKByoP/7cnHe/lOsK62t9QNlSm6u1tmqowdcfGB
NhqWV84fLRvzRpnfXNzbyCFHIM9jYJetyQcAlv1zMUqi/rDAZ3JJJsl3wKBgZsePYiw4a4r+P50r
EGsCgBAqNSUarL/zzz30Cg1ROIF8e6UnSGfbtNVpB6pjyXgeTXNX0Z30dZXnDcgpeNSsWeFkD3hx
vsslCxoHjhzu9NduHMkC+8MP78Q3mekguzMvNmPB/vxAWvd8LSim6BzeNVxXjCe3qX8rksxirIIz
IMPz2GaXUCGPhVuw1DBm+BTtvbh8+J4cT/AUcypowvqjx4sqOy+5U20rpeVzQxvj5+nacyovSQDq
JnKWHImn1p3gOyBQvreF0Aw16zitQMbqLbIPEumJTgy2krIQgI2BY7ZfZsNz5rrIPsAG+DkKanpt
vCTMD4EjdDjwh/8H63f8q6ARgUULRO/Fat6ce3dhsBdGWnMzFjl/nbgPvCXbtSqXJxFcNz2Vz8gA
V+yXP4DPWE0D4/VNTu6p7HcFG1NL+4Jojsaqs/8RzWcPvq8aEupQpERXDrSQIBBaHiiDiHIoJrho
/LlG46ifXLgUxsayTPnAr5oLMy25xPcFr+7Hznulrt2Q0j/9DGc15t/TRPCorhOdCPAGDFkisx9a
O+oFSC27JK0WLzVHVkv0uwSYJgfoC3yi7W3Xo9ShEi1A23Msn1XzQNKctLH3M23aNcWrvWMHszpW
jA8PokPKlFJiXpHVmtAaAEoiw8wcI/HbE3Ymo4RU4GAIt9H1Vq43TXCfdzAkF1zVFMB+hR1x13a7
V3Qlr6D7eWNjYRxGfI013oDpGQTg4tIqtkSQKzIwo4AAVqoZc0Nb6al1RLrECDAlBZhRo0N4DtLe
/1qIpSuO5urR8gj38VAk7nXEEWsnJ4iEQ6xMgccfpHtkS2hhAKIkfvYEZw2mvIXHtezvntPgngSI
GH1p0d53QpsdjloiFS33+HRE1pcY36/qc8UsL4ydOdCdYafPRqntJb4VkrbG/N2RH/D4lK9awpCH
HHHIUs2pFNsUG/n38SffPXTuVtB1hdQ7lmb+iwpdz5dOvGnFHKu9cy6XhFCJiA9g9jVfCR0/h0Mk
1OWGOOgUAYVceVo4R6DqMo1f7se/y2/Iyk2wCXw6+w3HUHIxgVU93O25VExbGxQBHDWzBXCQrIZO
5Cbi+XRVAXC0HliEXb5m//aDgCs+fZM6//XpDFmRr+Bt0bOs8pOEfziwHSu6LqMpbv2pvfK6KeVT
4bpS/C0a6RG4pcCOMg69lobgK/Wwyoz+3zVKptuDYC9avScs+qpqGGY2WVPQywFCsfjKKA06TS6O
S2FBDcZaIVA8sW4NfD5v8nbEI+aJTl3cMSOljTf1fNsKxs2qFSp/GA8Oas5CCkM718wuVqKKe788
woAMRx4PWGhhaOM9ZI8naFJCMy2xPeqMbWusJwgtgpBRIf/iyuc2SXQ9nvAEwZ88NDdAxFQ8P+HD
b2ft5bbz8z2zI8xykC+iho64CgoXd+2C5u9HA2TQUM4SqOXB+YOnFSLv0IfWHdFlYUMLSl+ImEII
Cg9pYJjC7Tuz68Ej3Xrafnyg4WQe0+dSJJBtGTdGOrh5r85kVE3EdM4DQQfO17L22CB3BiSslSAG
AkUEJGVnf8fscG0gYVtYGOmCrxcg+1JnvSb7vMjJQWLJ5KO9hOf8jNGVgEsIHlbS8OE/b2OzjbXV
B7s+9zjDcWsGkEcL/D76ReydxLjMXgSd7OFwJ18RkKGvppXRAhjZb6BkgCo/zgpixAGmNs+/ETn3
Barz5JXQfvPWom51kjLYXlMZgjYbPUxrUW+i6wRHCcrUQTe316Ivred6VwWLkVPXfDpcKAScm+hr
03Gxw6WJnaFvez5sPUndj57Odf6W0m/cA3tPvha/LqvWGGkaW4P+hLFeZw5LBflwMUyR2fZD1mgy
souxLZ5BbyASyLGEU5cl4lq2zUUPBz318ApwHYSR8GZV3NzYix7TwH98Hg/W/lXTttcfvqw95RHw
KVM3KoayIh7jG2t04o8CAkjvM+o5/9QeISb3BPhe5hI0xaXxdR7tRYTa0vqdTn6b7Cn43dKUkmwA
qJAqlzVkeijVQ0qknwyjiqsu6ZBKUOP5b1GxoHxuEJV9pEiOy9TTj8pRGzaelXnHBZdKMj2YvC8d
5Mr/SAjIVcBr7Quuuc31CXueoAq1+qAOrnFuIB41+2y7WEXAqtnmmsij0BGrVYXO1Mkm+NBqL8Bt
hnmHpCucyKDgl1Fl2P9Obkl8Je/SCtgH1oVKKQXgY0prrfrKCV/lluEzLkmAwTNNYY7Lc7C1KKNR
YdQ7N+nPuJTxsYpuM3GQYayX2rwIf3FEae1ncdIINQlFTBSEEGPdPF30cQjuShQYlIsMp/fIC4HL
MDsHhYHQpy51kxk+y8XWz0K0n1gKsUPRFGI7KhATxi4TRrcT8+KcUTSBENPGOMC2RV+ypBedu4pZ
jAQxRf9ABpR+Xs80bjar+iuH84QKrRhoEAYqW0j94/3PyBRjBpBvCk2rTjtZsGURzGc8DtZHzGGP
S7cHtb9SrxY9ef9zVPPYSBmgx0NSAA2UUDLgcr3Y3sSCIS8c3qH/YtGOTTsDGgELjc2rV7csU4ut
G1gzR06a4KKyBl5EcfoQ/7OBXJzZnSGGP6a1hNO8pbn8SNTxgxkUtkOhsrRbDCVeleJr2M8UUw2I
83mi92eDc6+GjNYrTUaFzqW9pJ+YIKQm3U00sns3vMjYSNi2tBOb5ry0E8UaA5sSFyjOyN+7MR7u
HgDmB1JsjIjLAd3jnEsK4/YcMkdfiVPZBSx/L6UPLwjMjfGd0GNe/dQT826RQmRRg6GeIBkqm61X
Pyea+Y44EQ5eO95xycfhqykpfXnaRnHV9KjjP7Tgps5WhRyOaKX0JtUq4HPe/m/MQAFxxhnx2/Nc
T3Q/3xx7mtXfYRrA/XVAXjs1oy15c7+Sbonv9hrQ5NOh2dHwHIGF53Hr2fbvrgzDM+K0CjL4bOM2
Sey3cvU0XJhFzVBRvmIScwAXCVS54MHd06MZINYQBP/Y+bQFJRW8dviGSe2wiTVhEXNpV/Nuccnp
C3nnpfhgnM1FeOa/w1n+aLZzw16dkF87tvH7mrA95+bCq1C/awBN/iusUOAyLBF2B55q8O4DnKTb
rPfhV3AE8jfwjKizsESUzS858xDH8Ug0Cpg5FFaWYAoUN22E9jdIiENZ5I9Fwns7ElmSsKaYyeE7
eMdF9nrpF8iXBtPrVcpN7hGEtILzrwBxAAlX8vDCvJP0YdPBShc72vyjAIV5GbyXeyO9auAX+JKc
iRcpI/r8GmG3E+vSK8igW+7EYREnmM78G82Zj9fW1/J/5GVZSL3bRLhYPdzhocUGwKBD2CKE9x0w
5TTGKlrnSAvUWlB/vytsohHsA2cgWM01JQXQjbfkMVUpMf4O//+tni3Ghp+tjNnfxjDUuiO6TIXV
svGM3fLr2kUCphvMoHXFi4ueuJRDndnk8bjDE8+1TsmiFx2kP1qJPlHJc1E4UrLf5D/yaV34HR6c
gK1mf7jjGMb0LQ3HSG/xweoA3VxkGD1ggEsxnZGCsrO3tCs0xbSM1l7miZ8GGUPN/SbJK4c/4ajD
6f43bbfTTyYNLJtP03/SuwXc/z2MFMwxW01NsrAqLReALI9D7p0bIB0x5WC7zIRhDJv4HbNoNP07
w8szU1M4WNegRoaPp65/whIJVbPNCHsVjaYJHlM5OFfc45bTOkvVunXpPjTZH6Z1TO1iit0ZHd9Z
FfDRnq6wi8Ve3pb7AtnaImon/E/nt/bGHB9HPWN7NJTS5e6/ywsCkkGUy32ziYlmIUgQ/fHbdskd
RgvN9aEaaR/dV2/lcWIGaq1LvHMRY3mNKhYHI7uoBmgfxUWsSpLT9EFckoe7Cp24mO2fapOSUdim
Xv8wajDC77eC1da7WQpt3ZeYkG7inBCzOnG6njxGAChmYe83AOV38DXlWmKVqzDoMwLafZOl/2No
aRJl26yTcoi06vEJen5uqbbP87SZHSbCl95EVBeUVAxeePu8TV4d0E8+EewuvpIQ25p5pfjXneAh
sVYV1trzBVvip5Psw++DnJP5p17lIimwcf5nK5ZcmtXgH6LnuFq9KVVwWueg2sAcILYTPIdjr6Ah
h3rpMp74HTgxPl0YsYI9U/+xzkwH10uHi00QhLL031nMNATz4+FbpLVXEyyhLc5lD580XZbIWBi4
ZuzFz2418Di036i7cQyQzA07Er/Af9E8YgB8kRdXxEmsAA8XLPtxUXgkxjJcla4ueHdiTRJuiD5z
4ZI6HJmnuL6dc5D6ONxexUt0fbPfSu8rAEjMqaLgr2aNiwLsNVciECCnfOeWqIIn9CmUn830lyaD
ubCpW59hEeW5+p0HBcR6L/PeuLThK+r9NQBtgA5f8fz++yubWoVaf60NEj3jBDuwP1I4Xb106txb
7I1lQxJch4DdForHMioTUPYOXOGNYUp0nMCTOXrvsizWQ4hBJVBLN67JAc+FvRNpCPSd2FspD0o7
zHUBNl20IgD+gyPUAxdRvP6EeNF8eDIGu9qPe3m/eNtmVI6qng9viV5R9E334AB+2Iez72D9qaTr
8Ds1Ft41jemnBZLBp2IWD8viLjBbcTvkrdFXB5CFFBswWwA2oJNJA+OIq5B/BdjRUS+gaiqCPw4w
lYsBlTuECTO5X/VKPRSny+QZP5mFWKr+0dr1OY3Ueakh5bOo702osfHfdzGV5EU39JkQJrOHQtN8
HUzkPquKmxEojRtqmnPIEJqIg+FZ1yqxhHrivzmYPt0FZMHLDvwB0gb7ZcSB4m85ZkVIU/wGzb73
0JsEYAeTxKA49j1uTHez7LIZWWH0P716VqS3aUCPc7QES6z90rBQNxRxgYrqK/5nkg7bSiZmYYgn
RCjB+rlMWChdBNKUbTLqLJ1nFSLWejBsMNIi43GLhQQOTdla77Js4qxilMNXZoO4wq1bVr1dP0bw
/bguRrz3aoxFjOcajrLXTzCl4SH2jy0KIydt6xVtr9RCDBDzx5jhrslHUjqRM2Z9IjbHgkL65QDg
SA6ABTCypyJfCsb7j30Mr1iHzBfHZTs5TbRw/adwp61MqPYFDQI4SI197HapT5tJeJNeWAMfQR8O
E3MHmSfTiH71aHDRD1awvOVNwN0tzCuNAGxHdfoo6KO2HM+IozeHnaJayw/5I6mcLy09Y82pPAJe
vsD00BdsFyb1aSln+59M5g6l/udX9jRA6wKT6I4tP4bVAPaADt30N9ZU36f8P1ZAWoWMhd9mTay2
MmbOfnze8PO5FuwEXPx+3EBvqhBy06EdkFPjgu8MTUkhxm/qpdA9qZ9ppnRJbFEQgZx+jxAubtd/
pkT2NgbnV+aW6+aQINH6G4M1uylnI+yWSdN2WfV7RIqp62XTlKFredRUc+wmpQgQwa38hN04mHUw
88IbguBWV1Hb0cEQLiP9Eljb4Xc1qDuy0EdV3MYsgKqVFP5vSP+Zw9+KvZx4fN4k2N4ubPqImJl1
ohXT8ekW8Qp3/19LBsmZgOznZzrtLrdpoueWH1KRItjSP8ZRmIRKDo0j82mrEm4KiFp0tt5MHamM
aWh3hncU1owDiu7X1KjuSJY1ym8527Av5dGTobB3Z2tvsspi2ISD5DUaJvlmHbhT7loFz/lsLPqn
I0yGc3DQ649VS5p+EIaKNbKOOcxb4T+FJeI5k8sw7/J/CD6LdG0T/MisQf3iYUlqEZ3tBJ4U0Epd
PSvnKaDj+NSS9sJmfqRMol+xCDYooON+u2ZHmb074gdbn5A/3UWz3yJWN2EcXunR9coJZDls0sWk
qcto+ee8kPux3REu4qcZdu0dU524Cp9ZLIUmnFVlAe0uTbZabJqClygizSRjtKxpv65qoCxZcfZi
99st+pvRHEq9iPLU9v0k6sWWBgDO4T+CQhq5RB+L2/nl/wriPMn7JGLlOc7CEaavToYKRiGKU4vW
eIqRELp9KpvnclpHVCecc5dbipDRGkz+w+7m6xBblbOobIMEDKRsP2EjnSqPQugTACTKMfEcXML0
gze0b/5fLmBBN/5E45l9y0fem2Yz5Om6IybubeKPJwAc3E/8djU2ulr0ty1lHImRjknGibPntyxB
h5isZZluwPvCjhtuKDEWbXpYwlf+qTgVRjbMyHRxmjDhyfMnuypkso/xXDBvO5OabVeVk2Kd0XjK
+QlavxfONgMjVmbMxMqQr3wWPViKjztFvBn3pzd4kaX3RO368+WXYjVjQKT9t1dollbI0EfIoekn
ocC+5Uyzl5GXiJf4alpY+1qOv+euyfEKKJ0Otj7THhEdiCcy8uqroqP3NFtk+I2YOD/5tmolWNAB
PSlr4z8ggKRep+yp+/9GheLTObDgUH2omC4oajHxPIe1v8MAIHggAyl8URkXPzu6jADtMUS+wmPF
i+tR1rMRpuubw1Z1gbzy6sITmJYd0bIZnOpy3uOvBm1MvWLGpZurpbkIHlGfVBnUBLm8QMUBnJ89
raygk4ZRo36p7loIVMMfNw536IHGK6+8PryJ4UEXVmGTTDyTRE3T46yPyX5AQamXiq1SijDBfavx
ar4XQYYdtwm3KZeYLw4to31EkOujB3bW7QrMqglP8uLWX7vtWUzgWFfkPhQZ6ZbMKs5hbzNacGFg
vKB1nglk0voHo+LAqRPBsYcWWtbor0Cj1s3w2rFUbZYhOAYo5QnqcT3ssAsmEJz0choE1vWs2+4y
DFrPnnViqOh245QJYOHHqjDppykPttn5X/caQkrVO8c/S+eB+UbPvD4mqMnH2Vw3TIUFl0GwRllb
jPIqpQH0og71Ws0k/RTHdTvqbpiZdbMXOWW5/LpvKcpCME4IzDIyBzu308mTFYrf17We8E0bpO/H
4AoRGlbK0cEgddh2AP+9/onN7YqHfduM+fGLaUpox+AgurwdufO2dY7IOTjCkO8RL/TsTWDYcTBc
6rqOPQrKJpqdgK8f3o6I37aQqjpf2EKEv9h+x2UPl+vV4BFyUeIOeIInEEwd/SVFki4KT09XBJeu
RAyu+3N6yx0RvKTQIiUgqwbT8XV8OlIaUtr1WvzyOl8MdRbup5DlRVcSnB5GkKtsK1palbM/4ZgA
RA7/XQdTyig5SobBNdK8CvjONNDkO+hzrWnIBCXGkvT4zm9DW1nmEaL0qV9QU4LpNgQBiGw7r6wv
qtqLGW+TaFyBMMwRfZ5VUaqZuRn3Sj4XPRmT2foYVCD7HlKnMiZ1I9CSjNvrJTawkTjIWLONa1Hq
lvxCKhr4XjWOd3uyrbSEKD1HNohfLkLUJNB5750JWwmIFu6eDktkWmwuGS8oyy1DfQkuAzeT1wj4
9TIkKjC+7a3LCujG7/3TeQ35YLeYRDd2KR/ovbGUQAZPXYNcrhB2x+xZPopUfb8MuvmE3oCkF6e1
ITFfmv7i0w+0LrIpaDh3Wv5M8dICXSeuCSMt5NmY5dWyhdoCIPl39gI8vWd1qUPlAV8CobpwRZzj
tkHCr0bb6rAgOnpzbOKnKhTcjbLzNp+ksHYEjM6AsAxQkVMl6duKs1PtT9ZuCKSZFXJ2rNAlOdGL
Vx919aTCYc6HnEV45edExaQgT246SAFvYuyeb7jeDS11Gl7e8r3eHCQ1KzZG3zlzz8nSi6HoBzZj
qwaWOAln9mo5gOWlOEx9VnnKvSLWYD5XqBNe4Ggcazk6Qb/t7xJba3licwMfvXoiV6cq/5TDqyBB
xDo792ljkbmFvdYzWawgoMsuW1UMm4sa/eHgZHxF7CQ6ZuLmBAlmzTC+v2fJWQ5hRQU6AGfwoFmc
5H2sqB2aQG3qoPCkUBg2llau3L4kTnm4rF29DpL71qJrjsEfu4iArkNdpkLY7ANV5eyGu+/5oqfu
x6Q+4dInfWJKBOqdM6fuaFzQ9re9/6v57AfknkM2XIcfwkvtVqjJXHrovIlCLJhq1jWEnbCQuZIM
P76YJrwnMVlNhTfSNALB06+1/VDrDG9pwGH0jDkMHt9oE+oH7HQtL48Yjge0hza5MWrGTEx0wTVs
+ui8YVP0Licd31aEeA+9qnEI6m6hv+e85fk/YVPrnWFXyGYCKBb9Hj1R2kj9/NBahXnlL7FviSLd
KxEEJLGWpAMy6+7vvc7HmN4lGcQis4qC37QpI7TqXQ2rF0b+R7kh9w3UkSajRLKwXbhB1nbxoLsv
nGyWSoM6l1EmHLWhNG96TjQDNocq6KA4PoQ9QVibK/WOoaxwsAJGnjWfI+bSHl1TXBDMVpQdgUGJ
GH5KKNNghAH7N+IxteU5zvJwV249qFJJ/CgAZRdOnCXqOly8wJ4bRAx2gFc/wJpvtJ22VFTDw1yO
NgAeRDxSaWqKhFUnecb+zDUPMAbAarJhB5Zw4qY8TBykY072O6P5dJJYB4LPawaWdKlu+YRxFGPC
QBTWWtw8xm2fWvftiBZb7lotuo2xdOyER8G8ra7ynM5Mo3TvOOEpHHWz71Rnr95L6+3GL5tskqJj
GEjRHG/DtPr7hfqYlcpp+RHJEifBcYvytw79Xp5cfyHtuzoqaFNsPQDupGfetYENLD0WEYMcVXVD
dMlDG4FK8sQNFW3SnETXozPZ8H76GrrzZb1V5LpVPs4Nblx1dzHtPuhjU0rFJesfB/cdWLN9K174
b9Erx8wdeoRln97DzT1gvfSrAJUuCr1KMCNET2Gk8fe77qj/AgfO+s7RFI1OK6zz70+y0PMQPlq7
8RijOXKLIwdwHTo4oF879Yd8cLQn9KSTiss5GK4gIQ/yiNEjx9FWruWlyVR414qhz8VSTxBkNtDj
RWNc+ElqODtsZlWUVoSCuI/Sl6rO/ZYDrunp1LV9nn1PLvpWN54JtPTcdYEuFOw2FspLoX0OLGQA
24C0964JU1sgp3rBMRdqB7Vz5UrdfsbPcuI+4Qw6BrsPPBz2lPcQYVP24odyS1m87bS+DStpj+df
tgDPTXvsbRPSuej+Z5N0G25zjiQ/1IXzoturgcVD9JzGhkJjNI7g5N21t87ZWmaQ8+k2qvx9BtA1
jSrM+XrusRuG6lyOudAsfoJ8fiP4YCB6DaJw6PT/RS3B4B9UUh+EznIOe3zyo91F2nyH5O2POugJ
VPzbuXxN/DtW4S/QatjAdEPCBs6I65DFDGZIzzxzUJ9LWCnvy9Ump/139WZ19cBDOMNVHVlK1YjW
6CJt0nTV1p1ojOpAAOg9the3oZ9LWLLBy+EpIgMG5CCKw0xdx0sb0L6qH7FeTLPIJKVa/fRf0rty
o/yxRbn1FZGB5+C5KoOfIrD6kQNijKRSR8KwtaLPRzSAIqDYKuNr7GhdwkqnNsT1WkpX044PNHjb
LzuBGdk7rYSvz+3F2MD9ZeSSsmgdQ6x9jrphmfUbEUEyhgLEK6ipPcR9q6+FAbuQEPPqp/XMUQMF
oz1VslKZ1FxM6BZBLO6c63r0rseCr6M+Ih0XE7MZFcnIuuRxLfnZrMimNqvoKpL4Em2VdwisfpC6
XfazhAFFiZdJwdMtlp20MEf6KL4h70SsgGxj/Lk3Yx3K7rC6MD1vxdArNI4AquD8//2Tp/lXlbex
5xHLB1jrKA4UsA5Wk7MD74nuGapf+m0mqPuIxfQUcMMPJ4kc8KP4eUEOqu7EBIGAuMlu+plLv3dt
Zs+4Lbqifn07BPcx3CTlFi9EIoQRh1G1nUQ5/OKCLKnBx9uw1uXX/mQLKrUnwvEWIJaj8N6UL9aq
KFW+9Jr12hCgzXcx+b272123Cj+33VqgjkKVvoXQjB2dntrtudBg4Pe616uJ25TYdSJkSy4DDIf0
buvspSQrbeKG7iPX6GgZ4vattwXZqULZvhV7yES+SroMtORZ0/fPEVWqaw/+DBdRGg/NzyZmcH4z
dDrWeKcaFd36fU6lvHq+62GhwwhlpiJ6K5Fsncx0GrC1LtGgtVQA0W8Lyh0Cy0vPFvtAXWqmy7Ec
sTlfozusM4pAPGed0i2gXuG/ZzFSiefQOcvkGKKdTWhoWsLWIkNSOKImxXZTpoz3/rz58pAKCCkl
6Bsy9DXtCyrUSnuGqvf44QHylgAfgj6AqTymFmJpFZM5BRKQFxNdjnCKLFnx5OrOSij/oUJJxSom
JeaNfmFIdvLfRof+SYkKZVKTLw8mK7kFG9zms/glVV5m7FXHZ7VJJkKw7iJOcnyfDjRUbix50atR
7FT3rJDd7/S4ZeaA8mSf15H36JhD/ybeWAaE2TbtnR8EbbM1aDTq7S5fjwXvbZilJOkK7Z2q2cnn
ubvoJ5u2MJNTFRgtRKFMhFDjRi2tLyh3x6iJuPnRVUvvrSi1Li5IWyb9QZhWMcyueUEeudy2sSEx
nvlmHVvNaO34ClfiZX+7e4y8oInKRQOJe8QlP/421ThMqFbk0obpvgCV5/+OsWaHLJDyAHOUHoUF
xDBs3JOiNsXwJKdYUfOKmwSlrt/QpkN3xJn/5ytpBNUFcf1kVteZr3R6wEN5JICwn/B8ZtA1dep2
39Iy0tEkkawgLlqRmq5Vb3azG2hsfRpwCtgUqWmP2nZGJSupFHoCjeR9PeRo2/ipVONVAMcoxEt+
u6TB1am1DT9siVrgJOKn9DrmvRzT16ahtcz6677MtFs6/02S/Hkq146iRS3S3eP6ynSuNhziWw4N
/qZOYguTzM+kvgdRVFZilHbnCd7AjQG9BoQbCbpUcbZN4AEoUWLiYhP/KF6NwlOdI8OC+i4L4ekf
eqftwqDrjpjkKn6t6gXhn+v4MM9TJYGnJBsYxt/wSP6txc3Io2yDxsv1ucF885k7RbyvjECSMu4I
Vg/h8s4VrEbZySf8WvsAWRBKcOL74oZImcnf3XpXg8jphTdrU3Qt65QYLYGjMQ6CBU3ZPER9c1Ts
elgMP9hTnMzfUHSoMIlqz517++ItaZyOZ5THjef7DiQ/p78lxJIwGoMMnPR8G9gyV1Ie0uCgK9un
Nr7MpMSEdh1u745y6V4fByLWIlLqJwypWOcbH1u4/eAxJoiIs/4ceMypDYzwFoPvYmKuQTQURdbq
QA+ijKL5iDN0/KZWlZbPmT/1f0MsFLpi0oHHEIV8yDaiv6cmfq3Bi+QwU/aH/1T59ZI6qznQSCe0
E1LKr+kfddtrqAlAvR6Aez8em016hO/kiKPgv3e5aLF4GbCpibu2naja5ylROyJy01qxJbpiINvh
hGfeLCJwJs24Z2M7kFWPG0sLP6U9OYAROIEEqvSx4pJI6W2GDFjlk2O9fsK92LLe+SJEEi7+U3QM
uiubLqtBEogHKgtAGNLXZ/oFxSmL97WUJTDxEWrxNlybZWRteUEvg1ckIH7O/1uMinFJnhFusGXP
0nxv0UF2FmkErNrshNFm+G6G0/lm9a2rFZlnBW5hduT788ge0OtmuZlceH7kaEjSlivy3hz1Qznd
YHN5bt8wG+DTzhoI3ok848fBeD1EpNV0Zf5mN2BBSOQGT6NkOrDyXOLc2qKLeBYHJ35qVZc3rCjX
B189O7acgj02BzfGMH6JD/mmA6lWs1tExN3xIHxDZUA25w5Xc8/VtGfpRHHKKqpYYl0689V1sSex
HiBSdE1f4CauILYyyBN6zppOMTvIs4dpy2HEqN6cws9I2PYMt0eLSocItQ/xjNnbnQe7vIJlQMyI
Jrm/6ubNd6628n3FZzMxFpXLZedYk4dW9LPDwqJwoaqLXcBNHQW9iNcpeFWzd3b/5c5zcBADMvN5
4ULfhrDCCV5ImF8xHezH1k0ewDVpuIfP/cKAtzjk9x8JRs9YNVVFAAm5JNQTE3E56OAAzzlTZfMY
gRovnlVBGzIvsps9mHqUkis3ch3AtJ86n8urhlq/vq41TWPqVHbQMXgXJ6G/fSZj9/q7UTIx9oEq
eZprQlmpWxQ0jT6hZq4YGint8VKqP8QagbM7lDANbEqIRxbAGS9rPtkNEQeGooaigOlZc+/knvtQ
1pCNOm9t6Op0iHRwjhkK0RNXZmSOOS2uThEIqdvaCl9IOLIcvSiXpaeWO/uXzIjnLGSYeaSRddqw
4Rk2KU84SD6GtYmI8nyXov0PBqRpE9nf6H6sA0gxGA6LZ2wHPz7SMXRZrRyCP9wGjyMqvcy4XKjt
CfdpKrDVAPzbyPv4nMd6Gh+I32Mel3lS90KzWNf9jBIqJkxHmRNT9kPs+CcUVKOHUKGQqzqTxv1t
ca/gHDMmqaLLIoMDPzD/mILG2upjFxhKh7Bkb8id85uXKgucCeZM3Xs9PIQ7+jUCGItbnaVnLMGV
ggp9rY2DTBqC/nY09AjMptgKOUe64WliCaf4tLHm7Phq03oW6FpaKceuj+fgIrFsN1OOM4GKMS8v
32dpyBdvcEEYSk5/iQll49JeH0Iimfkp9ZYjl51bNEIHwmeb+1b88UaFQjzpPkd/WTjBM1BpTD7E
3XoO3AtwEEDzwKOeAV32T4GW8EL/hGfEZLpiDAazXr6/1PqE8oNS77VmbwimrHWlk5LuJR4d8Lmz
kO7IbBVFnRjsp/H28bYWciHp71XSxYyXMshtHtra2W9s+hGnpzje14bxjBfX/NJ9I88+zg/Zd2cg
akPS+6fuVNbGomFi1CMA8mxBKh1ijVOxyWyjMOoQCdtdA1RpC6hGDD67z/t+0DLrnrGb29ZESrrb
rue+0LlknIQLI8+QlmPyJXNYclH3aUmmxTpjl8EfA4GG+02GwMyrVmRnmp9mBgq8ykbK0HcoFiik
J7GnqM/QVtfsqS7kDZkElIvGnRbDG+qJkJ361LXj5HF5RNtnXestCnjDCo+MZGzW06R69f8Sz8hN
gWEwGiCh3BVVPbFtI8V4sIT/Mn+6r9QSfdcU67kqNvFB6su1WUVLB4Oc34Xh8ro27YPSMlECqSc0
MrGS6aQ3pJovD1fwrK1X75jhpdFSZmyakTaGb4xKhQ/IaLF2wHi7CGkKzBClti0tpfB4RId6L6/L
/INxyXC3gP2uccuqRPgxCLuy9ECs91RHdVPDSv/4E9WsMulwczTF5aSU6sVpc2RXD9i75F/meEp5
hFvcu3HwYs721L2G072Tj0AY8ppae8gq3Vlhhy5m46zjLIrwCZfUIGk9WEDPP5Q/37g6E5hsgiiv
1kXHVqGwdElsxdGnk4Wf3rrzXnUMzF6G0BmpFd0ODoZXaO+aR/H/k+2mv5K/ak8MhJatus/yt7RW
mpEUspEQzs+pXJ/b9ZBB6qoUk5iHB+RE9nxX1n1J0T3ujEAGG91xgxpzExWTvvjJJLc/bhNED0+8
ndlmPJh57wvwF8NHnikMR29B8CGElfb6Up0nVEFZLG/w8VhYlXm9uikv1AJfl9UqUaQQPR0v5072
838oLzAbgHx7Y/2FokhbO7o5KJNoCAFFFxWfDANNC6gNyG8wmK4jHDoWuujobZZC1YwMmPirUGH2
3hIkYJz0FHNtLXDTq03DMceY84jQcxiZFtuA16olap5qlBjKLgIvBQtOkShokmJhr2YWNN++0lZP
m4lkx3zUH0tTTLiQzTK/rWenO81HVv9+auHi6CAQHiGKr3FcpIk9dDgSmyVfuVUexrlaPiRMHpH8
WHoNZsg7Ybk3xFOofLdw5E7lsI5oYXC30iD+Zagp/18gJ2//xN//NQfD6+2B/SR2FUVWw65yoTmH
97M1zNmZv2///jE7lubAXm2Slt8uiOp5v0zWH9NoDk89/xLpe5vvsNcXTVQKAvZ7Hlc2A0brp3Iw
wzEWxYMrFy814+Pq5PqVYBiLxCh+os27r0kjvU5KKWGfuW9EJDOafWlaJ0rliYR7vxvIxYb7iBRy
vwkTKMPfq+Qr3sKclAOYK1WLhaYzE3cDcQH3vfWa/Hlr5XF39769bGWQB3B3WAgHhzfMieLqGEI3
Ldi7DGOWIA3pvQrElzJ3hNsYoDRj4yngjgt6WdSfhLuMgDZy4JhOeYuuosCl+5H7f1z2RDAqpMHS
rWvzqH87ZhHH3dzBqIPwjPDKW2NfnxlbqrVa6dYR939QLio4Knr/0lkcRm967WcJCdya/PVCZeor
YloNnKnXS/5BRosCoh4EnoNwTZNNIEzFIX6vVm9ID2mvWAu1BODwZon46at52t9EbGNdqESuW8wp
jKE6WwaGKmJHe/wu05h584HvZjxvyVxR+lvhVOedMX7sWsK+xPYt3Lgy3Drc7cowAQXxqT6MoZFb
uF4J0OipRCS64SpAiy2Bi6WBzayxqg+J3CLlIM1RgVoEGt/C099YhjRJOPZ8EJtjxq6J8LM0ejsm
U4T7JMdzXNqTcvbhuqUoPgaUrFbCW/ck4OdOb0ZfBqXqCp6yLtdSexq+BQ63WPfORq98PlCvAAoy
L6Zk84CuTLj7/KeRqdkutxfAr9eAaYD+bOpnGbsPastgyU6lg53ZKIZSJayxpqy7hedJaS4PKNZH
zOB0B5A2mJC9XJwTBiL2XXTCwblyJcscig9iyX7GPByDOoQ4ARy9pJrQqDIpgKS+rV2LgnNkhrx8
mvng1tSy15e0C0At6ia3mfvYlsBB8Va58eO5CLJ2J6IBg6JUBU+lRCApByGtrMhXi63TMIuYRD+z
HjfupJ/YV8bSdCnXR5Uo29s/zZC0b+vNqDJZnerd2bio+DQY32FCU8LNWA2iVsotI4SeY4oPEruZ
VhaiuFzjaM7yhPles05ER5mN1l74Fh1P2R6T6RglCVK36ghloHMGAY2hcn3jCb0dHNIXg3gjtWT0
C/z+LLu1pJDSf5H3HwKfYBs5+2APPUJrFOCoPlUuvua73s2ke664zdxyAIx9FFr9n4UxXH4Iskv8
SaVc0R3ZbkPJz0t8eX++l5+c7I/Rms6gqApZNMm3+nQxf0Uuc35s179G1oGOPpYs5JjRJL8aCfup
emZa8vdEZqDr8MHIFfpHZCI6Rr5taxKMjq8inUO9KzNEeapGBHFafkxWlfJUo55XIsAwVHO3NUN4
QXuDbZXrDF0RptzQigIGvMuqkKIn62NFFnZ+UL6RqH7HayELFLJ7RMeLSRwWfGh+qaBHeJlMnm9e
6+2gsI/GmSSUMZKUXuBc1cBVxHqDCtVSlNYwEBeGZEMuRsdUzEyswy4MMN2S937/yBykm7Iw7/4+
jFUkpHdfF4uL6K8d5UXmNKt41wTmiM/G4TLQMi3ggS1T2GXi2vWrsNNK8W8OztkQn+WrBCi8Vijy
//XIVqTyPYgsVAfOJcw4DX1uUsa+xtSsDtf832w/eODY/2xEvxlqIpPCijTL24oCTYEQXoo8Jz6b
rTxASYJC19Q6LTUEM66TBJ1eLaQhyvJ1wiXx4Bb0QaczwJtiD4GLYwYikMkoC0IeiFvpCsfC3PpR
joSrAf2eQmh6ZKekkZAmO5R9xs9SDWHnY7cvUmfAN+LijFd5ez3t5/SHzIZlPNJ+2m8rGp3/nhFI
N8poXGhce/i9sNG0HFMXER592NcH6wiq+u3lhH4r3y5eaFQ9U6q6hrx6lhWY/SX9ofE+IJ4gjGS3
+gHMV1kgrYnBgqDN4xfAVor9xQAfkcqH2eg6ShmaBJBVM+5r+H39acz19asKu3NZxp+Mw+tQae7C
ZwnQRlQrwsMcXU52swNDZwUTL0KRy4wOBLI9RahYUDu7I/mnhdTOXN7/JrbrcTLzwEPB4JlT2Eif
3192e4seQiFwXS/2fe/T5yaIh3fy6+qOPGG40qP2w89ZdmNyZ0BWh1eK3hW+qHSXa0P5MM0cTxxS
EII5kLtFCWQjpqFY9Nq0e2JSyltcsDgWMbexfqfO4M/mxNnVQeN2qlNwlTuzCtKJ62UJOx4eQYZD
sApL6JdQN25/tkkw+hBqIphPXJTffLHHDnX8bBsaRRnbGp+1GeF3qB79Da7NbSlcS9vTXrSJ/nXM
x/IXLs4AdfY3xUR0mKe96iQw3NJgG3cx1YhGbohp9HEY7T6EpzOSRPtgQRkLEf4lYEvYv5Y3Qyfa
bcxDZMd7h3mEVNUgzdtxE+48CBVbdvNNCza+4IqL2kM9F+8mDEA8qTj+Xe6poqVbSpMAoY5jvldY
Q8lk3FKh0kKdXIlt0UZ3Fj9inPJMsnK4Ice8+FcPOe0DuBQrxdR1UNF6TDMLxB0oicIrvl1R/79C
vRFem+GgJiXP+xdvXrkhsUuvFvj7Lr2tHeu8SG+HazL/BnQrfWbPxLeXbMlB73Nm+HTCpMe7vIiR
r+vdDDyXpNbXC2z8ivvvqclZG2oz+kHmbYtOLDoPr3cFeIpwcbie2/Gyl9SSr/DZRTaWEb+VUtp5
zhV+E/v2MKWImvGKF78K6kGRoXnUs8Cxdu/YST40aaA5iOwQ7lLZSvZpZaWtNTPgr7AhCa7Voi6D
qLB7udw1WVyf4CCFZa6UuKzbY4j+J9UKfsN9D8zTH3aqj7TILZMMjGe+fPP9nLHgbIrg/KYK+XLy
DQYKZ8T5W74OHile1Jr5QvS7z1HzySw8403gl8X+u6HljcTciYyMoOv9apHJei+tKK7m1LIz+qf3
REoSDr3yilWQbanJGGCrBuS1q2hdETBJZGFAVWDrc3089CNdOdbGu3Cuqs/nCIY2I4pn+lQlLbAt
Bc9Tql7uAy3WzDEdJCBrRdkRCWCy+zm/cDV1I5xEjR/iTK2hVIlmLXXVtrg1lfcVMN/ROq6x3ThH
fajIGDV6paQ5iTKj+zF5Rx0nHSwv2TvJt9rSH3AoIABgWZ/nwUXmB78yyIY07OvDWm3G1+kKdZ+s
T/bMaAZHAKELzyn/6m76oAC8HOhxL0SsiYbKr7uGCVVlXO+oBRtKZ7aipVVU/YltQssA6t20mFWv
xcAseuf+Zmq5jKneuj336hwylSB8T0ZBZ3XlNZv3X9dEeS1y6/dgkwoGxoSMcHSReew97Ks6dSAo
5gt/VAE7e7pp915NHYAeNyeYA7CovxO3kEJaifTHHSyMVaYe/MlQHOQW2tSgL6b+q7xCB9M+VV1F
Yb/HMmzyHZjDNJP/RDdA2Av8DEACJ77eW89taH6qywULkHgU5XyGd2QyMV8FdXJSdap5V3Jl5MU/
Ru+0joETgKjPgZGlf6EjpTtApxV9KhxAXtMcaz1SsKmZe7WFsHUL4vhbYhZARfeGNSpDCr1hi9IA
UMbwRzR2E41BQrI1L5HRpN0POOtCrdCSPG2kbD2X9ptAT2cA7lfLGyl5OmXgauntzHAwYO1nM+dg
0VuwV/8sfrUKAqsjym4eMwT7O+QypT/gQaYA0BRi1p9V5dJxAilorbgnqOJX3LfuhDdeXi+IltE8
nOLnxqNwB4Xn/vLJcOalHf7m89Tt540ugy960VV6r6I9RpWCWeIx91tq5lcdMD2Tg2lwVQwhpqk2
Vv/Km2JRsn3OovmV44GjiptEppH4oA9LaqI4yB3DCEmXTm5870FAMPRM4s4vHmQ3M4FwUC5snvsw
13wOFSQa9rjC+dzDNSgxvbV/CUJd24/DbQeHwnJeMFHiv0xQd4wJRFX/xpypb57Scx2tdOUx+NuI
oimU6MUv2xHGG3hIbEMsz1Xi5MdJORUswTBwvW4fTPCUhA0joUoQk4gDRkAKphIsoNhmSRj6tKvu
8FyWSoNOmr5+dVN15PDDnEKRxeoi98kAYRoORl+dD3at3EOOZ0WQl5JWoMBrkPEq6kP/q5qEx7Yc
4W9t0b9wCK5eaAlIiQMGcaZNuZ160Dw1unEUO4gTI4fka0kug9ymBqEeSpG1RRJtMDVZsh2NKVlE
oc7Q4sTzns8kRLvAqsXslWtus2f7LCz3mdOtngSQC3GdZ1W6qGY+/WxVSueqKfhOGh3zNXi15KIU
iN1VDmC67pIIolZSgoVYL6TzRVw/urehdsL1grfexkxuY5bX0WZcBCfhamma8/Bv9EZy5IXMywKy
fhQzLSi6oN9R64Hzsb7OJBNESOYFEgqdBZsEUrD+befJX1AA1oUXfMuNtTa9GfYK3AX5w7us/um4
r/Nm7G71e0RDkjXnw3xJmZ4uAVoVDf0QQ2yvyjsuBeL6Mi+7ET8tCrKc7okYUVIthxThT4aOueo/
MIEaeob8SxFG15HYzC5WpKmCeOVjnLOW+Evox2FdBC9ogc3JubEHu4L4vVW25yxMjqd6/DQlgoYK
82XveuOQjIhxDPN+jqEzapa5x/+rpCw4aEc0G2jEtJmP2KQun8gWIZgTHskTiCYql5wf7F9CEATw
AtdnvqpA2tNaO9HyUXZchF9FF6a/sCMUciqJom8OvX+G+k23+QqHfOOSurIloUWQY0cH4a1R+9to
kwFJpJW2t8zYCdZQ57UGBDGUtzD7H5MeH5/LixKOWltc9KLLTI70TOnNP7X/xK2L7iMyPrDZwTOb
VcW2JvMdtDgaAZoX5hdSJEMV6Y/yVLZJXW7qOoLGOhe7MpowNVtHNCj57tv5fm2HD9ZhtX4salw0
wb1jt3VLRMrmU1sBO8aHtRKjT/xailjDHy+sGpPr822OB1JTm6KixpP9J1uYuSS5oAR8E/WBUCGk
ytT1DoLhrxDfW15yWZ6oYY5em95ykuYJPCyouvCCTaksjBKbw3lAan4aFUUbL/6OsTswfGULo02A
RR9GqmqMXUluQcy6D86LAcpgyjm1CYAZ9GKmAmTLlad0DZwk2geHD84qX+myc9Z7bNBkASN292Ji
mk9iq4xyirJlvoThuHdFCi5ZCaCHpgNh6HzV2KapA8atfatUXmohJGuLoZEt/4M2iG/UO3XE4jBC
BVSMdxFg68ghHZQ981r4N2MADLDRs+7HOSbPkm+yLXAh9FdTTaSBVAFtKBaNZAWocPzd2TPU7f5Q
jeZjhS4EilDzHYvJmfo+oF148xAE9EyTd+JFJwMMvSpD8/X3aFmBl50Y0LtnwseCn1MyPDLO9LeK
VuhlAVL3e3oSggb85UdsXmEA5kRnXzKlLl1jvA2M58UuoHvg0eWbFzWq7V9QK4shJ1Vy/yFy5jUi
ApyUwTdL73jXR9HNNgqEm3XHIX3KbPieEJBbzD2SKrpsBlshed+rivOVZnqUncvy+RuIoNntuh7p
i3U3gBJ4q0OfAQdmYeMGAGi/bdxpLV0x/jDJVOH0xafWk0BjSSP80bPHsPP0ZKHLnlU/qzMX1Oql
n7t/Dy3hWn4Lcu4oL+GUtC/OrjjHzfNwOPWnE0MpGR+Vum1k3T3eIAwTI2CztAmzmTWJ5+p4580/
Q+o+6H5noFhoSc6RHE52D3lEcRiFTP3qqeHty6D8RKIgaOKTb1OL7fDWn6xFH4RiBioCZBCE14dj
5nPzEehCDfISQBf2jKXZ4zoKtc5zSwDRTyfWwwYhxaP+s909SPx9JLi93ofukX0IKRVRn7SUu1oc
gZ28LXG9rQ191OQQTBVrtKzWjBg7VJxgBCgL3KE//ycLAw3Eub8NS50L51ahNOqDUstGlwqgRogN
HiKY34Zz7gkKpnj1Iwy+5sDKVknkCSBN7pAM0RDpF4q8knJ2EtSm0to29ELNoCLL/bxjfOc6VLfY
U7CMniIsuQilIdKccvITB2+5E8ebhfKu3f2MPqYfsUpSPv7Sh863Cxt8dm4AOg7EbL86xRWEVJ0D
RTpa7s55h6wZrFjCePSor516EuiqSd9+AIRVxhEUwQu2ojlIMRDRMvVFu2OS9knL7HOEQqiEDVU/
QG6QT+X27jWzTblWYcaqBqm++mSjaNh90pFzARyWoh/4O5j0Pg34S5eF+qgyE75IznDw8uZNXxlG
74DjYwvQss7IdlL0iz+aJMBvzxfNJgS4Eu3FZVUN1H7UqAi++jrcxoKszus6lJjTg9rbRJ8zUnbl
M9d/X2q9MEnn3xL4LdKy80KvqeK6o89YS8o1Gnlu50B5jaKp3m4rK7TgVTg4ODV/Vugv8KscAEXC
PJXYiV+lRsu5sfxC/KsNmydH+nIBt7UqlncGr0H87shy9T9IHs7kgZx0HH7azJizVndxKuL7VBJe
2evuMIAFbbUy8IwjqCllqHIKu5BNqdSkuSyPTqR7ZfzrSRJSygRDwUKxh05tixSh5/OEezaiVpbn
zUsg9dhxIvM3GkvzDYEfpOon74C3qpIkQHeEaBqrjaplsfqtsKXPuKZKXKglIBHDSikCJXz7R9kf
3xykZijQqChxuvrnG1eePX9EatzACuuwKY4f6VQQDV2ZhFpwchALDe/ZkD0UGMODX810CbX+HiIP
Z/xoUx99zsZROYeSvzkya06Or6hkNrTHnZ5HV6l61Cx85cZe5dfIpqnOxWgXfnvnp1M3p+l5Si0Q
IRees2pgI1KrLe/e4EMgXvYu3NgytHBA9yr5ymgiPa8QjLQ9p1Icip2p7vokSQ0bis1lgRmwNeOX
XCt+TJepCiaNxa+By5+w1SbMyzL4+b908suRBnGuke7doz9C831E/XuzFaDAI629vmVxTHdmgpBF
Nbz53TdkW9teQm854eh5t5go0R0Clbgkp7p5eRuXI96Tb8jNOqiEkKBuwOUWhmNy3miNi6FZ+2hX
YQ0WPfQPr12vbTXmH+gXdHY+02d0pgBATH3f3VTHGWwALTmVT5Qarb+Y0VF2qGrWIfi82lkylsk3
0htgZW9M4GtwXQ88uLho/bHxYNnrZ/07rcuiPBY25rZ4UULP6q2VoXx5VlzcJ8b7fuSEOoxlIy6K
uWTqLrXby1/hRgineMQrpIZvVFnM9QrbxogpLjYU4fXaoU8sbHkfGgFvhTcfNZNBAIyZ+wLIQLoC
APyOkUA1ko2hqcu11wZR6iuevwLVQWUPgXhX0rqHo+434DKYBTzbCN/vvfOdpbHYyKTOO0BPIcwk
Ooj/O+wOIi4Nh1FYZTovyMLxF1Kd+9dk8qrxyDyaHD9wG1nImZQpPNyCpFc1EgpdbmKEIKMb7EFp
++kv0puDPLFUwlH9fC8huBblqIm54aRzTRhclIEhQRQDrqDzIrJBNFLeDUznOH0cmDgEJomV/UQA
66jD2q2hljFzWI5fsDAViUS5h2UfJorHztWFfjSfmXzohMWXmmrjYSm+kBX5wBU2FfGFL2aMC8gm
cT++DgrshvEW2ULn4fnD3vz2fa4Fur/lq+ngOi2wuNp1qFri/uL27ExB8sdLdJBFingI0VHD9SvA
FZqJuhEwGulz+Jk/MdY6SZDgTKq4vJzyLWL1lMOK6jsxt2EPhmfCA4MPoNQz31Udf1vJWz0oTw1w
57grtkUVgQl1UqMH1gsR6voJqCrNXK28FWSI542IBl0ccNUrifXyGzRHYDcBX8QV2wZu6NhKlIRt
VkJ7ZAQbqYqkFYerY/gl6G1S4PHBiSktJ//HXfe6IMeOOLmfrBMo6Ga2889RobOE/mwA3+brHP92
nudDvxM9TnySa6Z64Ardx/5m3dNfeImDoVecyrN3X3lAzAvdwuoLq9xJUA3Fu47TiTW7XeA+1kHf
CvaQZo9wQeB9PyAyv/ek9fGlptH/luTUtVZZtMdjAnFWp/hO9ziq5UyYQwh7E8HRPebHG66+SP3P
EVNmwrZmjnGRWuhGJdZP1MoDNQRsuIvDWVnXfLmtlAoOfcIdD+DhhnoRUURifN/1mTUyz6yUOpuv
PaF6oR6WrTHCQQvhfRLfgVBT1OWX2oeQavGccaEEpeVGYebu3klJ+9YhtOUvgazRIcpHlpvvOyjo
w/qN0B6AHmTMN3fCWDvFcGqq2UDeFJF792I5YRQhMgaBtRxu0dnkex1R2Y2XPPWr4x8afkNknLPM
c7rWHIZCbtU53kTzfPmSDbBqR1jiAX8Vs+OXeIbiwiGTHGXzJvwHm0115ZaQKZ5cOpl/pHvMaZxQ
T+1WeyHN9hGHzZnG0hMQAXeSNF0joqP9MIUjptmqpaorT58JDpwsO/zS0VPWmcjofR37tBsWFi8s
4M16+eArXx7vrtOU6/z56KcDd4T+LWlPoiuuZvC/bdpcHnuYaTii/dx2GnFKq22dEbqa4YWCK2vy
GPMIOh9YwiEwrjjdbL5SjqYEwUB8pM9mvS/DyqNJL4InIfWPzfNd0/v4/lYZyIojr74hi2ExUf9O
NpF62YLw0Dj2d336rXrbKN40J/fIxExoA0QqifxKqmpg0+bXnojv1pfkzx5Jm7+llpmdLsdZLBUO
OEsqtDOPzhXSrokv/dBAQ0Pz1hGGKLyirfsCHNB+9QDjWPdR2LcmVL9PNZwVA5nbQv+IRGkzvCRF
gaSZ2zmXx0S0onYjerQq6qnw+pp4hOYf7kARCBaZC+s4qs7w+P4UhBEgOpfVomdTpH+3lM8q643U
2lraxhY4oqNLJXHc8fzm4hpTmwawNwAfw3uKDpTRLuQLko6O9al4kUZCEnqyygwaG+cq+x2+znc8
eiPrLKSFTVpn3Z86YGsMrzg2Nzfq2070M1Mt+GRvIBWQQHYmsV4LFUsZs1bRFTlkGFTWqrVlcHW5
vWSEMyRv0hXReJrVfXrvLjbOwqSo5FODvi+e4En2bwv4INBU172edAUY9rpuB7E+KXwLm3j/8ft9
9Q0NkFsL8vg+pyVNPytZgamJN5HXADe0gGkUA8A7p+2fuG/yDEWlt04cQ7AaP9MuuWvbtntOTQsL
0OjoOCFi3jOIvUavHGe4ol4tUEnD5kmc1AYGR1W4JUCrtZZAYbXpxtiENIvkFBDWXmSa5rCmt8zW
FcCTsQX0+uHi8eA8KEeexGJTkmUtRTRocsuDcvtVihmDGpI5fS9vGXea2CPZwjEjvIw4EfRWLgT7
/UyWHHaGHEB/tZ8lAH1pR3Y8IQqol0GCaEkrVfPe9jadS/XQc+WlAGuIaGh8/GoHKvb90voJOu83
NwieutxxG378UH0iTrNGmOYeLI+NHFXtTNoNFsXqCbj8/j91/ySE3TXgvFDfxvruCOjKPTBjgCmD
SKJwlAOSxTEZfiBQSpMNm02MxxgrNnLYwWpW+QTkAwkq9xWz0hXsc2J9g9ZlcgEAuVmTahM9zjMk
uFrLM9gc6L5Yk3KTl3/h1/z0ZyJFBX2Gq13kmHtVY4aX3gIWXPRq3GQmQBbsFy1y/W4CzHyrrx6m
s+XeyUOHfATZ0j+LHdT+Z8QQbSEsQGMggr7BruhcQPEEYZcqeQkz+414wS5SVrhf/tcl6j7xm6hr
GRBatFieZshV2R3BlAAWaEESsWmiCehGp20E3b7ssZUcEJiI0Zjajo6O8BCMjymzBk1tCZUgxjIR
nK9TKVEFTuuGE5B86Mtou0efpfrlAaa+2CeiWHfbzp9twfIVjQTfj+J5BiJJfw6PK3mXAQcv8BfA
yY4S7KJgIJ32orMLg6r9UQFEr9xeW+12zLfhBh7Z7gfaLqVEmYld5xAFtI4W+P33OU1toM9h7PgV
wvNAW3R+vMXwl8t8JwQ/4K0c6+uWW1M9vFdM0aE3NDTYYWNaH2dpU1judmXglR4m/iGBpO7E+UF0
xQGQOJYTAAIqt0G0sCwYliUFRptObhzwuooBas7hlAXsS75VKfc9rAH8SWYzOnZZevCkAe3pL5QL
IcTAVCbT9v3iNrAAfR+w2EaSbPh8yLtPEi0fthUDj9IHMcdiGxr7niFQydoeQ+beUEPCrgvE+3CS
02e0oY9l5il/Xt6QrZdpYlVisFqVeodg16RKYsEQpPjZLgZFHr5PcbA6hwm08A41VKvklrg5VzBq
pqIZ0IZ2HmjEEjsJEPc8cP3KxMVNXrgbx+3H/IrJFKexvzx+W/Fgv3GzJhnI7l/sIhH4R+hMPrI5
p/L+LPUPE9DPSuPYKVKrTJ8P8+5dSQukw/TAfxh8U6anNfeHnRVbav2WbdQsOpUzPTPTJ7bXAeqm
2nAjLn4Wz5aTMFhRJdj3i/W804G6dIbOZygREy3pSf9fJxryMy6k7BPrJQyeJOanyNdEPQf/z71g
OqFjdjcKjeTpc5bFmzYSnCp7kh0ISfsG5NQoI14tv+4F5IwhObFTbgs6tdVD2LTW0OS7lBAguQvK
EkU1sklKKAHk6QvkuG8F2g+YWvjyGFtngguwd0NcHNUmPvVcFaRFaAu0XHDD8JK4yy/SJHyuJtem
X6jlQrsbphuINCVcyX+WSlLN2l8xG+qxoP0iK3QO5KmacpDD0u+BazaHNv86j7fFh3xGfPnK+der
1+Y/MrmtOrLDdLYKT/qU2XMMDuaOcsJl3xk0yTtnxMISNoHXoptxXv6IvB/X8DG5jMWIEoU5heG4
cjnJ6el6grGTieTPIcH5PKhjcatBDSo3PjrQgmlqMIU+QxvvZTT0ifLbrynZTPV9fUpjKU6dDMWj
GK8SUAVe724XV1p2t31CzPPhrZxZ4DlXqvNLVabdJTzPYe6VY83gmcIWEKN6NFUUJYhFzUdqcARi
1BHXB83BDMKGIgSVBfF1cAzSU5oT6P5pN2W9M9cUNBh17sMa9qDSoN4YvxZDaiogJ3zqjAUuSBif
LTjT3pVByzRTjr3qyIyBy1fj6aja7YdGH3lKmoDRkihT+zZ49+4qF2nUdWNAWdrFNraf9x+f5oKn
2uwij/wWWbmzMzzPJJl9pLuUPYkLgMvMgqSuSMtndFNN1Q3pdz7RJTmFc2OX5Wx4jyypzG02mjB1
YApiMcC3ytGNKoxMYRc49TPSNyTs05GtDAw8o4iJSEtA5Rt2Ih0JB+qSuB4sDA9zD/7tTP9kkrzz
8FORkVih+gHlcAwNcXmE1ZKO5drYXeG1no8lHuBpa2/p/pct952Dey1xpKsVCA0nBaNsteKvw6Mh
xqGMcXMJAyZmMS7NU548UqvdQns8yTKVRQtT+oJiLzgFpGe9S5RtxrpkjtnTwFXIVhamYuxrgN5W
YB8HBVRpS04blnA+tq/6FUhRUPRv672ZO4TxUIj/2l5b4KZHk9AIHi3uqMB72Ftl53KhudIXLNDx
MOU5O/bSxrVfeEVJHcMB21YWvUnNB5bHw0VctPB/a+zmRR5dydQyh5y00zA/Or1kVWgPQd1Oa9UW
5NNVoZM1OoqXncmjsT7EIFqGqrnQpQvCaQuR3Mu0IWvN04jV3K5HJad7VrlNE7TFQbt+3b+VTuRF
q9fDdmutUZxBoka7g9rHH+C7G3TpQ/+bnMYBco1DQCrka5KUHEOcMTHB5MPnj4hL6CSCiDRzlifO
uf6ci5KDAdLyGOT9WkWZ1n8Ru/e/eotC2Uf2OvuTmsLAQLDeSgLArgf5L/OGpzSvF8T5Tjw8Ro7I
UhYj3bhKB7P16PT/WweSfsB0dzSSVvcafzQzr4FlNHZ/Z4uSJZUjBzy8Nc27F7tPk08oOPgpNVck
f7U/4PMPapg2A498F4EkDkTil8DVRErJbLnBVCvWcJnsRMBlK+NFgItbQNZPUvz9tpy+zzR38Nan
1+ahYjxnHqJaWu8Ze8Io5UgcsZjaRgTi2v/566Z+VhoEvDYcmWwWwR6oqy7Xjis0yKhAXW4XNDYv
wSdvznN5Ek3HTZUEq/vfN+4GfhTZHcLAUIcrB8Diaf292Efd8RRaue0uM75O4J1Uxba6y86mkDuI
8qB3zDSbjpQOeyxPXhHl8Ag1CNSGPsdhs9j1kchOdku17y7SGSNpZWdawUdO7c7GQhgApDpb41h4
4kMXXfZXNv/9WKT8OqoO/WPDoCpe6vzBBxRGyXRswX8qa0vbIu1NyM52iPJQQfZ9cCpPwBVIuM4P
YeJUbFLsek7eg8h+JZaruICpiidPUBk4sf7UPZDL3m/52C6UUQzsahyWqBzcOzaDY5on8WcmOqTw
ZY+k9kUBnGWv+VtoiTn0LVkQfey55tYL7IV8ptw1xHG9zjcfvUafiDiiuqZTPjEVD2ovoAl+6y4U
jVadbIT5e/mpPBuY9q1cm1NRZcCtEoeTgiOIvy8EO89kUjVwmlLpvChXjjV3wn6x86kQ60isQEAX
QPGzvXyJwHuw5w183qi9PBr6f4U3Qimyg2qKj4+2ybgOg1Hu+m8VAsncvi4AgnJBk6bQswmgv1OL
ZrDdp0VHhYExvrKG94rcpZqFc3Avuo+K9Zhe3fNwkX1ZAJZdH4i3hCW54HYs3LlGjJXqENJHxbGO
eEEDBzf5EaG6MLI+gOl2mA69ToynI+Ra0gsPpW8x3/41DYKhK3tO1lSjWuO+Di4qmr1HdncRH/w+
qcqijuZ8pYEjcr4+bVpcM/OKEKaTGeIQtjebApdHBkU+ACk1l+ptHQSAiYHxoNZ4BPRr5BqN3goO
/rtHrctJhTMkLShyfPEVN/NWdRl9EWqSDtuhHmgPp8pWy27WUshlhpRlpYEJgd1OlZZ4ERCAF/05
Z82zCvPwPt4Zcde7JgjXGQ2nM9jQNvoQjwHkL2GN5Yyn2COD7h3IqY1SNgtOgHQV8rkFMvsXrrXF
qgDY+CtuPPZusr1CIaoSZc7sWufK8u6hlZtSOTI8TXvK1uFMrSBTSF9W5PqGWTQZVLWodLLbTJeK
kkKTdNBZUzbaKFW5Wj6x/TR4KANAVV6VEVRrWx7ca+fSvItPr9T9kgQtDQ+F7vPNvMUSQXQI+649
jNPZlDUXakilrNjh6NDZExAcrdBcNTpuPXIqbdcVkqxYVlcXUNg2uPzJdwv+FNj4G9xMPFycHFZ9
qTg1lXAThBqs4VUSr/HEguI/TmiV+Vt3T6AiQFhpOFUqqfFW+fH4KVP5OeVfd58gYIyre8+9lqBF
2rKvbghM/lkp5noOKgHKrmuoWvCNN8iJ+Bv1+C/IQFRfq8zN4VE+xZKPhiPTHv8Y+9Yb5V0/mHID
ftuhrxnJcPWBwstRt7s+SwYzBBPt7SCg2X+4VCvKM69xlEhghoBgLEkd3Krt/gB+svG+XPFklTxu
ZCnfKvLm73musUSWnCSiXPdelfl1nt2oWpVVyr7qkj724C0Qrr5CaImmYYmTsQwJkmEmm0biL6Qy
4Ms9gqpHFVBLP1D5IWcEo3PWF6GEvlHiNNppTFuLTRkVwOfldAtyp2v9M0HhvNz//8dhS6XLQ9Ex
xxTPOlo1wOm61j8CXIyu131G5VyK5zY0q345pNUipgpRE6AcTxJ3cXq75x8Alkzlfjl9ab89yPwK
UDxHJNgTmBocYjvYaL8bw4zqu30YtvmHCJk35UsqBws1I7BOWr0qNcePmq/cxeUIEDvJTb1JxGKP
A6inobV7PD8LN3TBr2MqwgmkdoS4pPGlBmAP7171aXWcOSSLJjpf4o3abLk0YX70y7Wv5eE2mii2
b2VZ+/bZEmqXQebsoo3YNX3v4DszUz5ymsY+69/MabBM2Rx6tVwlk4ljHhrE5N0jo2muHxfZnntV
U7pWIAwmYSwj2s/sz721t5OBxo6mjGndG1eTYlhdj6MzGun3S2Fw9Z4ioe5PQHp6aJv+pbaDOw56
7siarmuxQr1ZsLPj+AOWG8xE2Oxa2i11CRdeZU4Tus0BAUULQAnlS4QDjnlJlciHlcH5fXZD4wem
qonZr/9nGyQuhk5Xd4V4zatKFm9OUVDMRUNylWjqvAzvQygmPVWvCndF942nm+sW+hAhn/vCtxCE
ZgP9PNr+JMTizMKEDe0uDWiEdczJpJOgIcQuuV3s0wvaEqnga5oIoBhQStXlZGnKTgIzmZpIJRj5
UPw/NiMj8ZfYV4kvlGou2krEY0bJumKl0CobienlssEekyREAZCi+h7MVHz7S+qkf6L2Err5CzHy
vfst2rYQv+ZPLIjU3ok7eB+Cz/99xJC77eAXNM17rtV/9mfsvaUF1rXQaj8h85svC6CzOi1fN1/n
Cf52UzZCuxC1/vl0NddHOKIMIhttudHffnjs9JFLr2bIiFMeoXyseKwXtvEh5Hqeu8AgBpikZ8gS
0m4a4+p2c4Mgvg7UYa6DIjX2TprHPgKhoAW7B04eC78TaI9riu6IukeUAnvQ1MSWehYgzaVhtnNK
mLqMqAhPn3CCBusHfQ87bFaK6hYkg9r1VM4y67KVEhn8NZWipvo/jN6FhRfTEZyqWfG/NJZnfZpH
hTYWat6k1SlNkoLWxKPmXAhu4T81YxgXjPpFzTG9Ua+3NiMilyJjjCiaDU/kOr1R2Z/UfqhGTqnX
9MC7oPXfz+ccGOFSH6/D4OWcrNPnK8WBsYxO9rClwd6jN2OTOwR06lKJoJRQpwhnFtwAS6FVejXM
OXWIUc1nVW5d5mp6R0vMamYNsboj/6cQGxbCjtXjPcFNZU2lA8X9UAXK8BU5gZfzQtHtB6UYYG5n
+2ft5vU0eTUbQxm1HTuGP7MdJfCITh548FmxOF5diQ4kC3t6IvJDhapXUzrCtDeCGO1gSsMoQrw3
zvZIlQ7d+8nsFi/P3ZdwVgs55iR6IflIiLjEh0moFIVM806e+kZuDesrRWIS941/8om/YUwzEpYZ
9lYjTY4nGicHQGJc28z1Iukne+1BTh4lO3ldPxZX5YHzWDgEXZdYD1lfIBja/qT5LEy/HBRd801E
LHpGRLNuLi+qx1WODKFQxTII7nwhEKoXKg2ud8HzmE/9UL4kGcP1g8Cr+p/juGKWEUwJl8nLDGI9
uHrJdA1+QBJyJAOeUtZyb9Rl3NwRrnLl9HcYsey4WK6kZaRxYmp3x8eM1yGwRKWP1001JD7fNila
MaInMu/KOmlkIFTzl7scI+I1MKIuYfn7C0pnESDzRry8BcHWo9hwvgxQT5gYTa1GYneLVtqBNasE
fWJQ6AhTR7eabxL7MBGvAA2zx5O/dDQ/lXA72jUXeKRBdKwUfF0aaT+gwNHZqASYq8xo8bbPTfF8
HTZagHJs0SG9ssjQ/ZMjYgTdwk/rzjihnLbPIE4NNGmRl1L8tgEetJuHGJHSTcPf87PpVffWrvm9
uC0GEJUr00leGYKJMk5cQwPuA/Fup70uoM9zs00zA0uZ2IWumgoHEEWtsDZ4kodlO4FWvFijWYaJ
FSlBUzPU9xLzItDMg0Jm1IgA5JlZcsGCHextE5j88mI9Q8A2tnUVFkNnZK/kCyIYta93PWUL+bdD
nSOa0n4y7C4slTxSKbp4nRWLwSlgcMZ9wXPf4DU4m2Hyo4AaaRCEYLyMy/aAMpN1oTpGr4Gjn28A
bVHxC6ywRn/pa2PRA7qlHI6RoANbVPwCUIptbCoY+FAKKcZJEik1trxT7iGAd+gM8OuMY403wgjp
qpvUwWkCejrFBZuVPtxHj7K7rZKO9Y3LoHHg/cmBVqEKGUB9D1IrFfwUHW5+bPbD26hCst1ExDF0
NWG7OBJX2xdaf+G+M7HXvVUwItbsfRy9wmt09u54AWJRScLeFpux7zSiGAFxFWyFoHDvWIaHZqB+
F0NkM9wdF2Qzuhb8pzhR5Np3pMQ2nLe8tC72imMf5NI9iABw4gyAME3uqnnFdrmkQvqZJAzdPssn
O6Kr+W7xjs7ULGuGDh6ocTfLb6nFHO82gsAlWmniVtq7I1NYO3GLGm1L8r/0ZJmXFiQqgnJ3xujw
DIG86FdyGp3kN+ZhmeC72euinT+S1YAbdVIWjGT3Kd/Z3x86MAbMtPzGN1QMTYJlZ2pm88z+c/fB
bvmL5rLLjjg17099SwPG5RTqoCe+MFhHNvz7WbRGSxF9N9Pm5CqoIN1RsjmGCwmfhLj8lcxkl/qs
DT4vTjfeHnlH4YV1uVVzKEE1jZpv3lmHorFZW5Dj6W8AF4BwEUbmqbvYrd2m+DZpKhr7QWc1uSvS
jZHv2dLHaUBzVep/LPOrLmvFLx/77LthqXZVuT/+zvMytpiYGxRq+dX1F1vJa8vD+MFEGuALC7HK
TbxEwLXr5siYKh4se6bqHSEz9Z/drfcdw1dAVJrr8B1gW22BluC8acpqx3f/xzt21UOfYSfpPeCL
nsVNKs41ly48yqLjgbgLBPw/MFbjrGI3XfXRqtLKORRsqZ9JJURASW3Tc5q2y3joBFKa+RdUWAbw
dLql4NH0YCsWCLdM7FnqSACTvp0RFDqBuRtcq5LxD6V2+a7wabgoYGPGMNz4rYSsIEdVfj1QvJ3t
ht30lbjfFMH/0Y0z+u8ZKPBweyc5K4zAHKXqjsaaiyxRL2SLrpa7Z6tTW/t9cfzNdJ/P+RRnjcFr
DnCxP2bepI/EjWzNSXwwwrNrHh0KZuOONNYDOloIQ9MvaRqayQv2JmCz9XxvKZrn9dhfqnL/nkhk
ckUMpK73vkmaDvAZvxaEG0uCJRCheQZK6IPFAYzedUukhFBBP6W2o6ChIBPkyga9T2/NGskLFrxu
rEQmG9d2r9SMeuk4VEvGMVLjfwMzsSjJcehCMAXH0EaCR57MM+uEC3Dpbz/Qk1gKEzXl4tWa3enZ
e05WK+vOh7jd3+tTPZE2fmSjPDgt5NQAGGhJCC+oOsEjB4Fh4F1G5kiErfo1BAi+g4Dn8BxsN/o/
xAsHXgf048GQ1c/A2RbTxtU2osXs0/k+kSkwQZKtXdCssxAEE/BSbbjHgbcYx+mEIItFIlzFyqY/
wWvd3nDDRoSf7zutT3sXVBQlUbp3T0+PN33f1I/j6W9K/EM8dtcEJ5XCsqTTqrLQXY4e5O58vKgP
udcwYSOov6xiI7eckZLCSH99BZZ5ETveQ3AvD4GBFvam4yA28ASzTsXtjS8whA5HUsc4smXp6jjM
p2B5vU3iMftXrHjI87Te/m6yWlMeF8YmE6xht0GSxdcOUhOpXp38LFccNAzTsu8nIzFC3IuLNgNQ
LK4oljxZLOdtXTsmscuQ8KSenFSQuhaaJfItwChyIQrAWvYAaq580cKu70nz7dG3mLFq/B13HUR8
sHHM1lfMV1EiEoraNgkPxpTG0HrrQruNNQATGxxg2UMiurdZjKy0o+C8/Y1OsZpT9Y9xPHle6QGw
sFwYFwH3Wy1RB9br9kgdQMJClA8cZaATyg0hyAUkgaO1UHt3ur5azJrtZqrkzYQFbkRoCTqLY1+z
6awjzXISgc5I0RhKZcwQJnj9ycKz3qKcGJOCJN1WAy6POIWQq70C7Kt+kN0Gg9ejyrE6IUP/6oZS
cz1OBD1fYVaR7R1YC7DyitWQuZ0Zh3bMmF2FTWB33kY/KeBJgFHfwrZDbQNQ+7QxQczLoXUrx/bS
UvsC69xTGyJWJs+pjGtsOwVSL6htnS2cBpeCkfrLT9xHyDLMFYDVkIGtuBMjmS7JwKwIFMBwboDg
zXXZNeXWDADWI2AmpRTAxg8SvJc7zsQmdRL4sTtNiagebkoXKRXIOk6AxxlSfCaw4x0vEpyifmlt
wXlSD3lOcj9LZcRWts41cItWLpcnRs53es47NuYe35clh5pnv/HaLerk+o/2CidBAR/NrXlpOGqz
xWuu1/SAr4t56IA8xEkVfSLBYR3y9FeCvLZoDumszyv4w2jDYI3VlapUzLjARF8Jltm8JLBeLNg2
9pfS5zuah7e66lyxl5ftbIrWccl9hT/KFWQS2+eTl/tPS96EtAzTCuFEmVwMTDA7L6BAnvdzNL3k
gfMyyCPYzPgQmXcbU1UMv3LO2v1hwyLBLEZhxaMRkGdIUjS8Gaz6fGSv3zgZw8j6sJp20IE6L2+1
POIPtZyEbWrAyBmZ0aOqCHCoGAkLk+z8WkR4WM4H8tRYYRWLPgwSw7rU2LB16wERqTuHYRHtC1qB
vEMW4pP8rwFU08c6/yk3WbLOOuJjgYxesbJ4JZ68P4Sk4a1cDCVSHeMYqOL8VnSc82OsIniTBrxO
+3DQIMAqjVlM02ZNbjah4zMud2jouA6385aMwHjbIM2Q96qYrmWnFWr3Prp6u3aH98y0R6QpK9hf
QEzaP6pQB7ghVN8CxHHXnciMPb/WVRseiK3Oxu5+Q97ZfPeVP7CMU+2kjEPM6TE6hvmAU0np9J79
JQRRNyY61zIREfDZH+M6Nnyn0bsPpZHpkI1jFgUjaf17TQoBq1Z0p6fy3e2auDYPnQmlFjbr6InO
ST2Vk0ug8FhpA9bl6FQWILdCGRRhZ9r6PY1Rb9RaUsInJeauDddi/6jfVh8D9hRHFJiNnP+vX7o1
1AjjnaDtq0PRy8wopEU3j3nImRinVn0sLhUQsktvuWYvEYCwTHtreBRfN1o+l6oub6BQXQa0jCQu
NA280GtSQSZpf8iemOOOjwzZ7SXVIk9kV5asT1is6ZW5oOL2tsUwfgcHyAJ/HYCYKNxFP4q38O78
ynfEacpEfzE8Zp3CjSx+ntJjsdplbjJPR07AxBF0j87AjI6A8GdANx0+TPLOtawG8vj0AO/rMIPz
4RCWww51hRj/b3KWrcTlIwNGyJFZtmCl31YVUAQi5MIHsL2l0/G+hC/ak1VzJpsBQLWe7AC1nvhr
J9ahzEA1m9Fv5R8yvF/Bm4l38wYo0dBzInERV3079XA5/feGi8bfdxnqkzlkP4/ZnrcWNWdxFl2P
9wAvMRWw9myhBFFInyawZHYSjHnp3jQDTOM1TNENfh57dUSAU938QvylHGF93yfUXDxvcrDKNDKM
7OWrvb7qiknYlzlX70F3lllqSJeETOYFJHrYlVJh0lC+pwiwzERRJ5OltWku3WhScb36Mo7OfTYr
7hMYQvCRp2N77s7Bbu4rRA3NTEJvMjnP3zTFp1Gg/BtAdTqZGbwoCJw6EMNGwSlrJV9XZTHWZp0r
jo8DhMUrH7iGAGz/LgwP4CPsntpj87jU4DQeeSwGgq3fXZipyRKQspAn+FFNTmqIaHrG/uaOJZvh
IJFfBQOD4rCn9BTATX1AjK8Jm81HYRe7wERh4bsMq3AfvWm2ATIHe7LJ5PiWRCPT6tsCezafSaTT
bor3Jbm2E5ha5DRBfyWia0GXiAicrHlBMNtykJcNvFt8asfriufHG3+QCH2iIcKP0tO9faLIUL2y
zlEmZJqhC3tCqI9uy1cCctejC5sSdlrnrVtcGcjy/1FKnBOgm2E/N8bl6MudIpDFLkWpuC19GnoP
zUB8tnB0tk445Zqkc3iFg9v/2J2p7KUlKIHxh7Cpw+FqIjr9W7Spiz3m9DVhJGfxzrwmoZ4yzViZ
7C7Av0S/W927iuTGzLBm5B+K39CLGrs+FZ0Q6NoyUCGorE2juMCRrtAJGtxyy//zkvpYYUP+nldU
orAdx/EbSZWkEO+l97oGlpTZewN7teloxXVm4O2vvC2CThEHp5F3jLFcB5fb1IPGmSZKQ+HixJUL
s1ZezH20yVYnxxITVikiMXrn5A8BdmDnVPjuyZVMCvwPL2GhZulcAeP+J2lbno6BO+eSXfX+L0Q1
IxDseE6QrfA/MP8XfBjNeLsZWAlf2UgZoUA975MLYo2qYyJICXOW16C28i9o4z12sO2JSf7GQxgV
lJXygQnHWtUs5InIOzY0vgWDloWmZqttiTmg00ArzfVfJLUj2RG9SxrakrbeiW9Ge2fscJZRmw3B
gfUTijDBtSABJX+BZ+bhHOys+p0GqkhOD064mOkBM/X527Dow3teXFxcxc+KH1aGTJwe/eenJFl/
Tv2uWMiq4iBDmrp/bEFthlwV8Dh4utFXWltmSVOL4fvQ+pL6Y4nQUC1J3JPeoYc6uOCJEM28Haaa
jGfHbmbDCIw/lJV+0olkds9uMX5jjXbzqSVqbgicG9JTdAe2bTtC5EA1gmT7dHawHTc93H+WeDU7
SfpWs8ate4yXSbnhC+ePPU1VRjHIQ9pfmLxHsUZjeNbCDqy59z0dm5jHIjWucZV2eQo9LDGhoGiy
hHkDgnIp2/YaNeH6DUzWLhBjty7juC4pARqFhKlPwrGuR/WWtpBvezeCtl5x6UhDqEq0bUy9MUTb
478DaSHv7gM2pTa8Je0obHSnJcNiTIxKw16StGWbT6wok+c2r/CQse4Lmr02RBrZXgfBbobhihko
kyWufx7FZ1OD6pjMP6ILe8vx/DzdNIsoaWiRsyLFadIn07CSli+jnNkYH9jorXrnwObuvsrl3L0j
1EVGkUh7eE++rIbOSLfihJ8xoMIfyvcS40tTZ+3aV5aGTDKtCL5VDFKjzOPWawcFxe9dCmEK1qx6
S6wgHoovSi7aSZ5KhzO98fqzl261j5yc3IX7+zyQCt+ukw+PaXAxcvUmssvJW8rrREEA+9//1dBg
HTYLdrDXnfdWnKntNY0DHnMfKZtbl86il0OZ3cAi/J4B4GCRy6N9o31UwuKLIL2YYQ54q1irlIIH
rVv5WprJtOCH9UevQUsQje0ARg3iuhmm2nOp22xfZQ2e/9HWGci0AfC30+wNbzsLbzzyNZatLmNJ
sQndIQG+Qv1f0SkynmhCXhzEngTZBrfnDwEBHGV862+bh6YrYJHqyECa5tJn/LuDtBEmX1eQ/X97
W7Ck13YPzhpLgNSDEJeb7+xKCHJbkNZSzEwxOSy9BjxJDCo4gWgn9FJFD8LUdCtxnzOSTtA1JnAo
cO1g6dx7zGUfoiZefkkxCbl9se4lfBaFNbsES6JLr0Lr6xHdfmtImGVktcL0FwxoQRrFpuq1VLUO
JqKDz+JKvymbGAKhKPU1MsYbq1zJ4CKTUbF0mXys5G4seo1iUKR6P6+N4TddR3ItoGwZgO2ym2Ly
nvFGhi/99jK+PKJkIy/mAoXRbgJqcJc5KLeCvETK/g0xmsRRU9n9eYV9W3oWfCt1qSqC5qtYHf0e
NT6HxODgCKd3DID9mj7Dq7fqccdVcTgNcQLOUe7pS88BdxBv4/zhi78CbcgzVs4QdbkLDmUY75KD
zf58niC3VxnbIQLjxffRIkIiOqXkc/3xUyIik0mPPrcDbX3iyW2jviQBiFBz/wq42sSyZeBiF3S5
r9LrpdyY39t5kpceuDuIrv/MPxYIyBgn6TR3fSb5b3tKgfJmcHam+bbrbXEJv4hZBD/2QhvBFLax
ZOCNXmRMedXR9fDc51g9kIckCtfizfRKYVRNSg6L/RYlPTpumJPYyQhWUxEqjfJD5rNxc+bm1Vq7
flz/O39NetL35zI2KeuTUtJQXM6YchyzJThbcd0RoiIeD81n+Y/nr1NGitVWZ4RRqCaI/IC9Y1ar
kl6Ke7ag8VcxXPsWfQuAk9AgXq1lsZfm1crJs5IpP947f3VktaEio58cA1RDIfZ/uQqrDpCUz+pC
kWXlRnR3YVJcH0WnsLmomfusmeO61Ru/1ah8KobllVKLKHdwdvI/LlhqnU3+0M2Ha7VH5JqEwua1
/aohx/ouwmJk+rxSdN1UVBp6VKLXXBWDJi1rnvV26Wp4Ibc6EclH3pNM7BuTu3rCcq/meJbILhvG
tWZi8HspAfQ8lWSCb+QOLwqaG1qz5L2sbJvAgM846WYaSCwsUl5zsL/n5ZwHqfrAbL56RxVVvmFj
lD57pKkWWGChp8zW5kapbWeAnI5+nhfy+bA8z2EsiJx5/KQHs2rHtdfaD99MrmTIMfSNJIfkA6UK
iYqfZp1Xri8JBMLlUl0xkGtqNlYMF4JpnIc9KtNHpJBjoxZPdEjbTe8d09YYEg9IITVoBLcenzW8
HmlMGLD9L+svo3Ta8usY1qp1F16l+93ZLW4H3keQjm/vezNH8JhjsUAYIf8e9SG8EPeHtLjLs9hz
MqXve7aFUc+v0edBoVIOlMzeTs10kZF/WwqhKDRwGV07XmPo9RzHnzKFTMTf4rb1l1lz4MSBYT74
1UucStjV0Flzlkic3HXm7NDLzKRBuZcrNtXGtM1JLGT05SYzLmwn45ZkVQyoasDrSZbJB0VQwcxq
5vxXQ+F+skR+3fEq31kJY+74DbTXzvF0pATci3FMb7ln4pENZGYmHuh15uVno6lJ+IzIEjgsamHA
MWQoMLjj7Va+yMoaICr90rYequo/8q/vSOMsZNNnwNBJjwyAkg0RW+wHkJ8WREjkLZOo4G7tT9x+
8qwqhB2AhgDOiNOSYCIvjnzcqVTQuB3lCVxA7Zci44L6k8Cw7KbFauiacjLfE2O45tY2ALA7i4NQ
Q/j0H5iibcHQa7QwVD/99xokOdOTtvcVFUTrJY5BnxMAetkOrOfWUIDaVK2BDAemeakDhVaICSlt
yEKNl/BoRY+mxUVzKbsJoSXDQiGKNfvL6TmUXOJKU1oSc4LqDkF5mNSizuXs3KElgGTB6+u6nBUs
9win0yvrg9h7mY4GfnhJc0VUqGnDEkagi2o/cD/PbmxCprJPSjMJczmm+Lf0CGVzMt9UjnLfXFws
EzTRRh8YLFoq6/afCcKr62CafzwQrNJtpYt4VGYAunECU5eii/voLCjrPMbWIDNn0xLiH26/qaZF
015tAyuFTgZ1de4lQ7qx9j7budNZijAZOJkuSdqATj6IR6c/GXwUAc+0CaBKSsgLWqbhPeSCDide
9hcNjznqSjPifxA4mBpjLpiHlnbUazrkH4Lox2XOrHIfc7nXViU7bMxd70rOdKjC7NoY2tZD1gJT
/rmsr29G2frxDZoFO7zscj0vgof3tjjMCtOQ8m+H4FX5q5M2dMGEnMW6bgh5dUFvrKupS0JCx/tv
ACmL7ItFbM+gSOVse0shPeSm69OsbekOY7lj0mjGKOOzasli3KEw5sdv5/7bTgIdwZWesWLRvd6d
l5N3SRsBvtLGy7bHAhGXOnkQoH1JK1VE5WlrekmOzsAeHB7ZC2MsSjA34+fop71oXy0y6x5Yh6Sl
ROXYy9MIfA/ReLakBdo7EcugFsl11nVIW2Yn2RHVVRtBNnoiF94YkkVQKU/mB5CfjYWNl+AvsWk7
NuexlEmmUERTLm3i4d6HPMlSkcVW649srOeT9BiAEbvJtOuw9q5MlqfMxiwGI8BzQHh8GAtTepmv
2w2cD7uzWfEM8+zqbjgUEBuPOSPBKPt3WDcH8+PtXsv2fWrUs8/P7GBtSp32GE8woNFBNjdGEY/P
Qt8gKdFrvW6cfnptR8U9HwW7lZdfIO/S/GXcKLN37kmz6H8Er6uxdmxs6+ih2L3BNzpcF/t9rILM
/m3+ZWDfYpEtRtFFD9XWHR9ageqJR+19LjL+n+uku17mxFXq5SpXoWHrrEeLZ70aseduJwhFBZlC
V1HbiUpeVsCxDA0TCuO7bkYN0GHYFWi5Zg0KG2U1sVDPuEHG5zjOSya8+6NJKsPGXGHi+fgzlCxR
NwDvShrVduFAa62nJPnljIuedgwSDn41DVJ3iVGzstaQ1jDr1xZ0qt2zpIpAmIbtFGKnCvrTu6QB
x/HhTdUJVmHFST9uVe46agHYKfPiCg72m7hIvG3IDrlNwCesCeMNjdE/JQtqyGevd6Ys57TkgTgl
cM824o7lkzs5lmTfeLetmQ7jyS0Zy89tsaUVuU0nWxqO9RJO2f3gjwodUauj1KNIG0+oRlCa+MGJ
u5259cHY6EWEUAYH4b5Ha5eeN9Qk7qnOx2z006+rxUQpSV43zP97JXr2owgM9rkHxFMLovJkw6wt
8uHuYpbXilxv5LA1fsiWjBr+edcS9GnB0ePbqNZ1psrnP0ac+jsokDH//s3zu2+Jmo4ZWUQW3r1u
66EVofLoVh2ZG+3FD2ReGwSwLGDb+9oKBoAfgngG+yz+6x7awhTFjDQ4QvZNuSHfGs4Z0QCgV2aB
vM4uNoDq0dq6YasFgTAbG4SFFS0jiGKNd2NIy2SDtNLtzxgStig05NyNfcdQfin3cYPpEplOsl0C
s0HcHNusGUdeYMhGkOJeMRfeOzf5lOoGsx48FxklOhTSwYxOyPWYv+A56wDVA/9qWU6bTxG7a/AY
mno8zKdjtk/0FZkdyUBDF9slG/HT8bIvq3cQKuwAZwMBFsLFbw0YnHPjD/wTpuBwYj4MgGAK38aO
CsY+xSujFtmo6lYjgcv9ZQ0XrI4LWEspI5ApkxsTq9mCBUZCWERI+9eCUrWN/7ZsULakw7WrD26S
PW/6v90mn2sYZBlR8P0azKtSGFVr7sOM+FkRgYmCCAB2Gq3eedVdfoV8xyOf4k5v+h01MosnYcCL
t7OjmCDMkCQYD1ddGenBQtL/ZPDHln/4u0cEHLbdFJpzfIRN16vXIkzKq8XsrKrPGKfHVuAcn1zv
1OP7PMSrF5paS2mlOMafgmbRk/ki091MHpFtq799QDb1cXE8Ask8N2WQVq9lGYkJXMg3gJ/Yq6kR
J+ys9aoHitFnTfN6m0LDnv97yyYsTKq/dD90wtKJWR2/fweioKA8JgzeaqyTmpcseO3LW02c5Ldh
vkvtpzWi/Po34jKZzo0cxpLNKdnyQWrKMqayq1k4p36twZm84LHMaR6FIS6Jonw/M3JrN3/+Eg0h
MXfZoY4bFNbrif5fXKNihHg+JRXgg3sao2C5I+5waM/C3GFFWZwAoG63u1VonVJk4yZubcmwEbRm
6GpIHSmUnt91FO+/0LP/ov30rcTdHnyXEMYPA2tv2t4B4ZS2I+MxoQKrEBaiCiWNnbqicja4xhoM
kexUIgiMxA2R8HnObMhgH1MXQMin0m/WLClv1D2ymrr+e5Z/RHeZfpXDru5R5wZrm2sL8FUJyjfZ
hsuLm0sCOGwkHszcS3K0vumIFca6ouMh7ivfYZH/zZT3A8fkrWEteruaK0+7LnELJEOyN18lW+Tp
sZRe64jx5EBA1GW5Qrenkx/Z7QkHSxoQtHLJJ/dk2O3aHc60lxHOyQdLzGCEJyACtKXCePYbn8Jj
eGdt+P21CcHJyQFptcRVBV5PUsq24IbznZ729RXYaSOHt+dd4R/Nwox5xDejk+buBqFDCf0MczUz
JR/9M03JXG66cfDY1Xo44ngrOp0eTKMG5Nbn0FEUg1SQuAI7DEasgzYR3pHb7XC7C7JP9A33omMG
Lmvygw/2CqGVWe+UyZCrDI4HwGIxGNXehJOnr/r7/NKtXz0to6jbkJ2FVzNdwYjiH+wQwrOv1Xkh
/tu+gW6mMNO38V4wAF18KU6atYX6HnbysmWmJYVIKgF7WEsP/82P+WPj0J6X5zN4hm6WGvtlEu4r
kcV8mVsJrPw8Oul2yWOIIB8J3PjRHcfLERPFY32JIsSP6gj03f9pInDCy4tKqDNs02QPVdvGG+WW
l+mJls5+kzojmwhVKqDmGc4h8G+l/+1YtNR5u0TKwIHudg7b0tTpIVMSiWsnl0NH4zI595V0nBSb
RxYUOd7Jl+jwV1UCwsAsYdj+ngFyMwcbPle92dH+mmLTq5ohDI0iBculuhKpNSMqsQoE4BB2Jtuc
raGmM0YmVnsqN18iv3IsrTu8NeRR1jyHupQQknTf4ASVcmSppTd1v6zqNWsuOIls3haUJzRJUYGl
pxk7oiRdkpbVa5OyAje6lZ3+2tYXZOi/cw8pZYHf0hpAnKo+9tLlH1iNy0/q9ojP4PtGAf3DJDQ5
23PqeLAIo02r8OA0x9nZIIn8xu2EjfQqIQDiq1TKzHBVJiA8QMqsOV6FPxagw8lBLd0hi7XyPbYt
NR/UKuHkcrYN96fCRCGkBgbZyDMGvcHOwb23x5Uxl2IVUEK02zaAC9j6TXZrI11Wxyll9y6KrF01
s8rrT6RzaXanmx8Io1qcq0tznalbjbCnmd0soBgQn3bv4YLJs63fP7Nl2ecKAnsPbNpHTwF42JLK
g9wtb87fcfEtE9cLRoxr35UgDmjnINfj2qEbSn8zjkPQ6NqXdXHF8GTnbXWjtkZ08iVv1ggg/mG+
8VWD8HpuDE9ElWZiueXytIA9EEmbl2eM31qhDHiCIGojy9+cv3uIEKI5OInsoONRee0m+cw0KcM7
ovPQshoRsddGauYwieaiB6Z10l7K1yTKh+1b2+ocY8U7P6275leGMUtEA8qr+JzzyX2vINcARnAI
Iq4w2GAbf4MDSMBc/dI6ehBfnjafgdrGxH+t61BuVZAxZfP2QkyvwlKZeWQXZGS7oNwpR8aBFQ61
hKhLFSgztK0cicKK4SEALxQ4YDL3yu9vQj0A0kufzcOttAhC4T7xJ0RgBdJ+3E5HCxYr8rmXV5nO
uQp1O90AO1pjSSpEmEmPNJ4t7Q1nh39j1I87gPCSY6Yf8LkA37pl4CgJ8NImG98mZZSGns46Q7Fg
Tb743Nl3OEYEo1QMvqjzBtBDCIhtk1KobEeiVEJG71RAr+r1x072YGjK3CnLJD1063AjUUSpWDsF
Gdy5K9lXH8+GD90FZ5+EsyhV4EADzovTwyk+5eB974FbCuoFcZ/NH9z7Qr64sW2yQ5vQpqi88rti
fMQAnzsTfnWITagKVMPT5gDu5mzbmi2ortFkIuhIz+q+MJBzZ2wtuQjvzfdgT/sZulC2oi3DmDoc
k7VKKOdsGatdtvBLAT1dMSR0y3yLHP1BnoAvrgdDN2pNXmPA1eu9ZX221F/e/VcS6dUtlX8mJjWV
7IqnKqTMnv11H/dweNkxdcjrcCPDFohZMEG4ia9Skf6mPxgJwi32LAZ2j6K9aMI9Yokuidn75UEZ
l53JqZBP8NR7fnftnhSY86+kWNTud8N0HF/Ezuj+Pi2cc3mQhU6BlMSy1WUJhtBzSKoY146Yuz/w
pXyDnV/T5B/q8VGLpdBk5rQ9CFqCtjF5oPKNyKog85/Oln1nzBo7YDjTH3c/9ZkMRs9IFTakdNhp
0EJBl2Ta9PcKCqD+gX2GufbPjnj6tBg2A9iLxEOy0v38ktLJ7HD3HwRsch7iV+ucEbjoqhxfEhNG
iUf8S5duQQyOQ+zQDp6/xUzoYk7wUP6u3CHPp9DrrZJvbQQih5b+0qIS7HCHVF9c71pzc45TAcLL
DW2uCbbP2NJy5uP8RpzW4CjkV0pIBgI55wIRyjHXOxlStEgeJwBI0gmanrITA5BuQgUMu6C//TEw
U+GPQx28UoCwaG21+m7lOw2TcnUOm0HoWlcO6luYP+tfHxHxv9NaxaK+k0Vre3iFMgM5FzL7gasz
nEtMptHJODXjAjHxT/o/G+DZyknELXw+L7cQcLnDMkCdILBIGV9qBOxR/Q7RP0EPg/a+5fSX0pgX
Y/X8sgQxCa19vfJpxRqHzzuPP8v+Oq0nSrQYd1ME5gldqr5E3oxUsZA9sV5iNREVpIvIfjPjSl+i
Jz1z1ER5F1WKzLmEOa3LQJvOWuWvZ2cMw1SsGeUsK3SOdKba6rBW8Po2oI5qIC8H/4G1tLGcf4Y0
dJ6b6K6ErxXW63OAWBXn5pN7IaIfHBTUWl8fvZwfkMHOwVS4Bi80KBkqo7co5ALmyRC8Ge4qAhZJ
f1vRjU2GX2LyoXb5/rHOvnzhjAp2oDG0qtOk4YYWhDUmvjOvtqaD56aUX60WhMAtJESEvIXcB7I4
vzN/ALWXr30bL+u0hygfb9TMrM2ECIkHrjgxYUXlVUCMrm60UMjXsXwljxdXKWe3I3t5B/7Ifet4
zlnzECban11kwAAR7TGu8cb4uq1XLcxhSQn2410GvfxzYfgVo7co7ceD69PoBpcjVbQ+0A44qVLT
FxECA6gZQlYyc5PHgMoxa+449VywLserfdqlgmPNOk50YKxQL1eYdZqOQ0/AV2VMeB8aEIYZH85C
8bVXeQyP2cJpf4tUAchj7sgO6FW0RyMHWInNpfFEbSiUavcYxoUaHA4v4dDSCGwPPO/pBY5hOHlc
+flHms49ox5Od3FwmlA2ruD9aV1UJPeEYAPtNkp5NgqmNzx8CQmekF4EaXojtAwDWGgkH5oP0ZT7
Yu6yYvmiN8DYqBv2ERLXLgVUILQwJ+utkf0qpCHL/9srO5QzH4finAET8SFEXcMfotdloCwoqxjb
r10qB4hbUUsHp2pp+sg2CRrN3CkVDJnokVtbPlC6auS/7ZaZI/4Mvk0MUs3PYAqT8hujXtBErscc
m/94qOdU1Xh1oTMB/fZjfEnnmpZm39BW6nqiOJiOaoNqbcQ4hhazp7qogSGm6b4K3F7lEXDBNVN0
Yx3acVf0FJiOACUhDj1gTt2NXlAY+hNASgSvncuQNDvMKs8QH4cNzkGw+0vMeMjebtTG6kSyAxGT
xKSxdJrV5zHZjiPoCz1R9Sp4SLIVtEigttmY6WlJz+T783yeJgRFRvIJGUrQpTNuEK4zQaoQy7tT
+ikPZihp0Hlxtv2dfzr1yK1xRt76NaTrV4yQTCS6NbeYhZ2VCn/y1s+y5WMDinhmwrApzEcyAIRT
i1HyZ5UX6ElA5UGSDPAGK871dz/MGEBCYwHZi0Bq/oPDN9GT5aJ8ZaD+oSgOaiblWspwO5bASw2k
wvFc//ajoo5arXOCiBmykFihV3JJnVchLo+cUy77JY/NLqMiUyf1F/hIiCgOLUpsDejmfAVa0dxX
oZGw0kzfSCyoUcHkVsMSg1NCbyt7Vti7I0EEJT1PzvnF8n9T0StD3oGXXDvFKW2PDst09cgSYFjJ
wd2CgVZY8Heuynvjnt/s9IgQ9EQXWh3SDWCKTCyEHGh7t9WRpohiJ8A6xaATU+7BTf40OYjoox7q
u+brWmA3bDk8oy0KierQ9+iWcG63izL+hbw26btwOc2Bxm14NJYdGk1m4vDPCE/GE9kAYdsSEtc7
8TpXCnZ0FTeCJ6bxDvpnrmHdPNf1SEXs+t23mQW985xTVfUiiguz5GI2qAprTpdWlcRqc4fjcghm
pp+lzWiYpWWT6PNuaNjnYxbURzXJy2nawUPAFLx2qepb7pC2mn4MkjvNY2SKpoNrF018TyFr4NXT
H9ZKPVqfWA9m6oc3/VeZbORzM/ur6OOTqBUZwyPoh20Fmn6/MjLpwuqDVwfBvdoUeB+nqloPAdVS
83+XVz2u2KehVhCLFj2V2g/ns98YUDeyDxFmvptdlKqMtcAnLKWYi+kJGTtQgUVlkO9Ph1ABrspl
FuRVvUccGpTUC2OVEJ+I++Jy11cJSA/GnB3NEmvYWbz+LYcfEgIQB8ZmzAQwgcErFXwO1dZ8mUq1
gR91JDEbZdH2NyO03CCmOnMPdlLvXC8hZptcbMIeCKkY1KsmlWwxx7tTS1qcuoxIgF3Kq/JQDVMm
fGf5F9gWzVqZLNxWiLBnVBmUfZ1q2cgE3nJ19qfCh2V0JrDb5A4gOMpJw7qPnu4AbexZM6alG16v
Y+tvZplYuEuoTA0cxRzxU6mP6FVODqwZVpuKDegEDjZior/z47UBviwz+gZyFbAhOaO8xiqELWkO
4hGd5G/t1fziQk3AFp0cgQqpTKhV3AfAxB45VYi2e3p4apN31eY6OwmfgvsZ7jhQgi4V1zM7T30S
SDFHXA1pTidAzu/GLy4AcLDIxJV/UJrzFf+pSSfmOzBmK+1TJok7GYS2SOl9Qx5dUqZTXGjV5SrE
8FlSeVoSXdG3J5slhiLOP7D461sMuh4sZGBs1HAQFO3fTtwsJuzGgJO1nTrIuPbV1+evoj4uDJ3T
MCEDiH8I0fTu47iGJjf9ALFsoQ8qQHfD7JT0aXaBKMkgqygxT1AuoYDusa+2+MaXsSgyNV39joBa
MwiMD5fdydITcX30Q5R+7IGnNc0j8QRpeUNzVv5o+0/s++ZiOlL7dUkJvDtdM8d+fBJ8LN+m9ZOX
Uqg2j4kyx6JVPtAr+1FxZcHpA2bUZTI5hpDh9rEkhK54m6p6MOvPoXDWnaZYyEoDL9EkaAUe/i2J
jhSsGMPcAq1Yzikz0ZlQgfUqp8q+PBu4A50Bf364kR9de8QXX0DuLdNDCRG333OMIi6UrjTBFVWc
OpWa4ZnudBAeq3bm0l4QVG/6Xx1KvFR9vkq9eWOawx9KVli1JYOE9JiZ8WhlGz737qaFNZWHeEVb
HPkvHQ0d/VErUfDkCJeDBNgOZPMjtcaN6GQB051avF+86WggsclGWIGJleDe/OPJwuav+iAP7mLj
VBttDBC0uq9teNqwYlsRrOf8cvereg+u0PJe6Orrnm0GjfpWfJN51j3Ttr2rWu4XbyPFipxsaNDa
B5uy8t9xM8jybA4x+5gXRUwW1PzSnT8E8SY0RkUUAxrwVCrvBtORbaNnKrutgIs4bttxbqUR1W+M
uXzo7j9oIS633f3WRCVW1l/GpojGBGW8alHykVGoqyYi2YkSzNc0YOY685/Z2wB8+L6A3tscUWbq
KE2Hdd3QXJZ1r2AA3hX150l2hpiQBNFkocflyU2f6bBog+/7UY23SZpRgcO3HsEYJsr6CCDgRjXu
ZvvVmOaZyXYuXmPy0jx7IPgatRMPHr/EzF+kq3xMgc9FBq/40TLr2M2RnsRbOimQ9bDxh7hZclwF
aCM0A7OyKc2NXViXATInnMfyKxl7y+0IUWO1CuTWm/lJg2MCXo+AjKnx7ROKsFrGXGDQ9DE+JEaF
rEuCdfi86dT+XHpWeuD0cSOsZA96c/rPw0OHwELAJePgyCECuAc4NfDCM0JoPgOC6e7skNw3nm5R
v0f/hDQiBxkc76MsttHWemJsVr9RfoGcWrOjpXaXzxpCtLU5RjS6UMgZuNhEemTpDXHwXeIjQ0Qr
APZPfh4zbUYv6JFEH7XH7Gk3QT7UmV+bFDqoN+nkGA3ttYvlHR+Y7cPYTIGYC4khSFOoL0NUxdTx
4ClO50AielUFD0iabo1KilA3jMjYXhNob9IgWXx2b5UWelz82RKGK2IAZuudXwpwf9dHUbaAaNGe
VpsupVduMerGoQmI50p5eDV5cjlg69leAba5TTJ7yhSRZWB6wVMs9JGwEAS8JXuB1kUm6YupkrUo
Yf5blcAVnXne8wXBpB4FrizfaGK1K8o75X7TrO0VvfQYF5/dnqhtZQ1v9k0eaBtwZsf/53Yih/h6
uZFanMAGzf5zrtllCJ6bCq1v2YzS48HTC49v25xWOPl5/j4C+Q0P7MDchUk88MGL5kGffpUXMDy+
a7i0zAQrqiEYUJ5X4p5khpE8nPA0OEGq/lW/GK7I3TbNOJ8PM5dtG7mcCrzv4tVxsAvUE3yMSPtY
GrmwNsVqK9o2cucJhO4QFzjENGTG+xwXdN9Pz6Hn3GWhUaOAuRRsCljlv9LxZEOCPNDIZDkZfd/Z
e8PwJVVHLNWpGpjKT+gaNeqAi6KqhzGwrWwRL0u6pCCMiwhCIyRFwcd1JvwYWqrTz6beGwhcIjvP
vtklkbI9AiwYR5g6trHqIV6SRzGwgIYb2P+Hx+eKxBsResW+bcxswtO6WdBTdu5WwFMRjmH3v2GR
QTvs7K/XRo76HXJyebNKzOaEkwMBJvN/e4zMHSF9lz/e7F/99wXyRgaDcJejjjWsQKrMeqfdmvyN
kOc4oh8yvwrSitNTAXpzFeA2VQPZlGWt1BwPf4pgNh3XQ6CMrBbTC0HU5irqrg2keVc0JEVwHLZr
pZRsXX6eJ/l80yJJTbxWlitGT0kF0uEiY0hcWBcmVnAVgfbpcui5Yuk/4N+qN6T7a8vMZMqLvl6c
BpN/tMn3M1PEOZv1Jt3nkPWD9AtWeUURaN+LwZp2J2426jpqC40xWGXy7KGqNUCK0tgdYebe+wTl
LETnEbKsiPqVpM/K7GHTTqr0qyf9f2sRA3uH2SBSItpoIZai7ccd29YDGHTk3aqzFbsKCpMg4c7G
T0/dAH7qbDZimalsNysWVAzopl3sieNULNcalT2pNmt0nfGfIO0wZEu7DKUzeP7JzSFPGH5QgQAm
WBIlwO/o1U9b+riDcVs3RpwXP3rust+IpJ1dPpt2omibSEZIs3HYLO42fkxTG/cxe0SraUi198/z
EbOcx/+8C8n8bNCPL7G4bX8n1cP60IdHWVzpX/BDu8vBE+OZPdqxrnZvDFj/Bp7FPNaXhecZiqDv
tn8mc9G6XK2eP5Bu4NILUF1P2fnKkmcerkafOBcfN/l9SOfCjsX/F9L5B+dvwxCX1Isb8/4kkvb6
9V5+2H97D8Zvwj0Gn/u+hAZ2APDN2gF35dUyCowlP9Y5rKsikXpJX0SH+IjdSP+iddzFldYV/Ooa
nZtzMvfNmeN6dTMdB36OdId3CqRwkstcu4PJXizJZPyMwO86XiLU3NklFfUd1WcAjs4HSWx7VlxO
ZXsh0uJuZxeAkrgQz2V7hoo7eeg3jAAIt7pvLrlb3k/ky5Ww9+H5LmDchoAwAclw00YFZwb+HdxI
+75eSIsmGfFwtj4rwjfmnR3bbgCpYKwB9L+f4AEGZ2P+SCr3ogF5nEBiABwbWklk7kwHid4C0FSX
fZvxl1d8haMfLKrd7cPM0aT+levQfJyPE4T1oTSA9/Pgk1zBQIngXdH0nnvovE9bPYv4yGSVWT4b
u+jIzVLcK07eDXvFYsitHvkNmdqSyHWnjdimR64Eor2qAWDKzTAYluvDeIZGdbZ2BhQx7f7NdNjY
vu4bi9hD4YEfAII01L6NALG26kuX8InyDwYBl4qI+PQQI2plSjosQ8gYt7yUxDloAq6zpfV3LgCt
wpfBKmqs8ecb22KmH9DyGpE7Mj00VK/SXQlUA6JKe+YXyUjnuGTTei/ltvIM5P3eChweE/LGJEnJ
AHSUK1EZAY/9wxVij0a9VRqP3+BHHYvTrkVyPa9V85vaIVWzp8vd5m0JvzPp8Y7SdcLbgzWUS+Ng
JGam38+C06vezmmfl5RyZ2XPiX6iW8mIoqxyhKkrMvnpVboisBgM3OJvulHZHN+TmLKLr/CbpfIr
DbqQ2NjbElXkuU9V1s4B6WD36l6W+TdH3IJvy81hQWw8zfjQRGbiUGPji7Ofa3wUGPxuszs1ZqDA
t38u4Tko35jtquf1vQPSgTL4mSTq9ZOR/zhyFfSI3DRjkp0cJqrXqu+tsji3HkwDz/pjKG50KrWF
2z2aOFWymv5Y27CviDjYj5EdkM2IJirwr08bMxZ2R+/KnbDPZNBpCJ0bN/UM3E1GSyMwVp9mTn65
eNf4DDdEkTeU9iSSRPjyhvJ5nwCJEB/UIxI0TcNmEzqc4MpI9o/3mHVKuCOHcukN3QLtO4dn4T5Z
9/J4khX9hLMQRIxiWlaRK36LxnB1gvxuYz8XLf0igI72189qoQr5Ca4k6nm6UdRXFkZutiiEatTl
4L7CqGiK5RNMNBXmv3uiVS26RXahLckc08CpcbshiazlN133HNIOD4a5CVOMVJG7hXw2V4aFBkPa
079/wBZV17FLnTJCcZy2gQVV1Onk0sbN61xDI5gWyBMrTecwLMxmsL9irKKjEtY+rQv6xVAX5l9W
hA4c/PbDpNwwDQV1N65bMvDyJKnKCQUAhIcCn7cNLwqG8rxUQnYLgKpfKqrzgZxE45cb9jptpfcQ
X1Odka2FkuN/SrZ0+FgCcnH2SfJYPyZ5/PqyAc0YETdGs+anQgwWTFJyiUc4jqvznMITpFhvQeuV
l9MOcSSTXaFttcdTa279BS4DnTLGHQKYRwIW/FuyfiIN2SSa2of11YyAy/I+kwkxZaDaO5Meq6Nz
dOBJXRTuSakC+IQtlo1WUdkSMNTEBnlZuOBR8dQ95Im1xZb5xz9aOScwl88rblhQOW5b7/v5ghNC
xHlezUfPo/mA5SVGm/GMUFI97Bs4jKTtao4MvUnuhkMKm16aYdLC84/gbZ/tc0iEk05+wzaQTTpW
VgiRzmVa8QJZW1XmtasmNw65Fv+gScoKeZTIpAiHq9forxX2nV85I9PthxrRSas2EXXNsVDkcjp4
6/aBiTLUP6caPIAl3x9g9JYz98+NJdhYGqdUduI9A7W0hFTc3x623G2lR4XX2BzbErWX9+JwLPno
Rmj5kpTjceNkIXQ6cKtJtMy/nJB1uio/C4SowbYTQtKb4N4DoXrmTN5xRNchOTDeUVgjdWceGZpN
kcEnktWlZuOkGwf2mPuycIo01BVIDBHtwzu0LcE931u8RKqQAExkULvJ2GBKHI9cBSbjx7UsNsL4
ylMwUFyfPRod5kJT5f8a+T3NeTrf69yQJ1M8A3vC1RFfEzewg5aN0dTX+32LXf/dPVzO90KTdHAI
y+cSOwrtKeyji34fzGEVWEc3PDXqChLPAZorNSYyhwHhKaOENZ7a3ZUT9uHon07WDNbW5ocqNwTk
TYgKA9F1TE0iFpfbHTCCsYMWK7uDBjhHMwzDI84cVBuh/g1QswNwbq8juXE2bQJTlBGtzWYNJGKo
HZWe3S3aFaKvo5huk3+5d71kPFg+wmpNfseqq4D0RKKzq2NlE2388GAOg3EMomnKz88fVWbv6TSJ
Y0E+MnUbqdKdD2jeiJ8C6Y5vUHP20Hj4tGqRVO6ZwtqZxge7f/JVql8HZcuIsqisbJHPduT1ApDN
HElrMrqYAJBHCe5iElwQ+06Y4XvYtdPcUTW903ilXASSXlyQ8T8uMKSGKSrg13YgvEh6pMzYa8YA
7xAjTGoM6r+pxofGGv+F2pMbHOnpyhH2tswZLDMCGAAWabG4Cem5VRUM1b0f2yCpE036EhAk3J+P
vmPKVlASFoJbKOfyzd4FCaVOm8/LKFZqAzQMnTk3Hd9Bfiqu2AqiWcnUg9w36BxYY523xknV0TLp
OrmSBaKVmWC0tho3xZl7LUMfM87EuWZsaGkC+LQ3gIC5Ge/OV74SzIw2NGPxi4sCSpO3GKIRTPSf
5AktzX4Q7REajqUb9seOONqp6i48rr2O9LriXTGr/UMJHEuOsW137+FtiPFyk5Awjh3k0DSoUmM0
bIXlhpBpaPujqKkXP1cPV7dSLQUbRjg8qZebpNx0vkb2ZqceesuMBBUS9H9jz04EsnygC38LesI6
IfPl0z3p4CzBSlQ+lSZBnHXlYyWDbYcHbW6x3SZn3MxEzipGulR5irPvU7il0r8nPU6UFpvwExJF
BRdvbKBM8zOglK54GsF+tA6hL+WYz/iq8RN57JDuGMJy+z6FMpIjQ1U+TpSSKYSWTPsMv4G5ZaZc
sE9E9oYP0iH9aIJByUSMci2Kr3NRUj7HrdPZ+TsW48f4yPeUFlR/IhbgzPCE3IICiFX9VfbN/S+4
Y3Igoeu3/OgyCGUcju9/oSkamPHTpGn3MgnkLSGasBWU8qLQpNeU38EwjABNXMELk3xAAX+ge6QX
KV7X1RoIcTnvvxlkDv3M/N4pCEi+aaMLowkHpGRviRf9WziY2Rs/hqv60dJgvZ2JQk2Al+8pKWiL
aLy1XqAP0b5boLtNtnHi/LwZexLnpozcw8dOVkM8R67HiuYv+chJlzMxNSkR4pcrHW84IZtD8hDA
BYPDU6QZeKTk3UyRy/V307m1rtHZTexxalmvulg7mssX1gJtG+il2ZmnL1YyMLVN+7cQsJPCURBr
G7GhgaTRy3OerrdvwyMn0ibAob5v7GqFI1UJXOHmzPbleiEv/D70oxeSsDAjoMqmWw04ctpKNkjy
ZycsVna3FTMrlTYKDk+a37CP8/Z3jSOJNdfp+nMSwjgZ+T8Scstl8vrkDMfjeMhXcLjANWofCN1H
+nlo4AhnLhk6RTWM56rOgFdidJpC64/ON6E5XqjZyxTrW9k5pl2BPATcE2W7VGtvvcASoQ0pxydb
NKGAXhvD9exoMfUj32estRMO+U1Q8PHxJfP0D8BxZ+kZg2VvOwc2GlD53eVnZ16TH2p0NWeHLRru
abMzmuh6XwawQ0Hazmm4nezSor+RKGMZJa9mDMJOvNEX3AlTpxKbqzG+9jy9o0aWlZ/fCn6upWn3
6h2ofR54L+sUfWUf0W2PNDevSsjum4GlBcXbNjiS0/Rw7D7L7yHdaoyhkBWPmvpPHWRRF++BTpBC
33t0P8sHIU+mGvPLhMiPVuozCdYePmRVtEHHYCLG1g5fDliTsFwfgpjjbVS+c37Mj1h8xZwhSv8t
HXtRgIUJa9hj2aPbjgbuDcJt3W2pSjN/VtNHzyozsuDXGqe2dEqld4r3URGITbhYG38V5fvoFSxd
KEKloWzM318oMctDW3Dr/rPqb5UqWLhznu86Kx3coNu3fqXbXrhmEqnI12U/kNUdnIgzkc6x2V9B
32KCR5X+F9bu2VYem/tX4RRWcQfrOvqwW73PT6Dyfnnm0jsKQFx7QM5m9f/Y3zCWGU4LdzfKAMSn
H3ZItGS4n4CtvTwrSWyFpzUZTVgqPlotJNhb6RZSiLQeIc80Ut1nmGvrIgQpfA4epMj4mNTKoJDX
2eOQWitSIvlGRsDs0QxndwcKu85o946Gc45Ba1NKLwonY9NPBX7azvfFW/TZy8xkuZ7MEOv2iPzb
v/rb888nLCkPrffVn083O90t6LbcNXj/hdoB/ZTr0O6mR3s16I59oW+asdbe3BSIjsjpQ3g925dl
c5np/UXkTiLLzf5aDbqkOpUDcQIcOodDNhF/jSAf8aDlj2fhuMFn/MyB5yYVMsa85etGX+7tfoPC
j5l0jMBdBtHv2jRKe36JJBC1zDsMa+CsS5kTH5OZJ8quA7KFjU+ORb6MyywcVBl/sI43x8cqr/vJ
PtWpoWMleAu6pQIf7vJ/GGQZqJQuv4xw7+MmC+ECwxGCUZUDiZSafPtw3jqWciaMd0ZCVpYGVq5a
C1zPRsAemNYsVMTTEFe6Hu/y/Eu4UxlyG/O5LVjvyGJuyIK7RDrcWwREU7NnCiHWgKVGiqRi+uUK
/OW7GZawOP573YKUab6cj6kJc5Xp8ANyJ+YpxMJNJkvkGFOZhLIxnJ2+SSDwBmeTP52EnSDqvFZD
EccdM3UNavJLjK/ALHZgyu6zYE/uFODPuZnPkJ3aPMLob3U67qpSTMCJa53uaMr5Nd5J/Czz3mui
6981yjkma6WRu5mSyb7sPF4zjZ2kLOJN/luV9d0jt44QOqCYpGUjMzbPTFBM5b+DBmQPjw85br4A
K2ZVGbubs8oHDN/piE1DswL1CQ4gCnbkrNSCPNVSfLGG3M/P7/6B6i1VhzerL6DqcNdWbAAbSAnb
+jz6YLJ0LIgC2veZS7YV4JQDHbG0r1EldlzjFqedjlTi62REuoUjEoZIMd5woYK/8l+u8ThojNzY
TUE5TwPIBx/rMyHNDO7ikcP36fb19/R3/URgjrbrL1rXPzuIk2+IzC3cw4iACnhreVXwTVBZmrto
Aug01iAjAOBqvi7nzN2+qgKz5EoFmPgN+n9fH5cb72VT4/rtOuxVOnOSA1vs8VMFtjQoM55KirVu
zqIo6dttfNF+cv6SPWpRvxj6M1nB3LJmU9OsqaBlnvmHCtYj54VopiF/ZcKIsibtBKt+KbVA9f3m
qh4rldtmaD6HvLLCp2yN5CzhuZs/b/EDlsr9CEaXbw9bxK2Rekbm01Hs+KwABaq6Kzbdt/EJJGyO
q2MzzeiIBa6n3ROTKYex3PdweghisF1DsikdJXqmFCwOcSwLNvRwGNVMdNyYpDuXW5hiAkYKS+WY
ExApx5ooRbhDjlvZzKW58SYnGQdvVip3Vxe6ShoKG7KNicAXiQcS4CKEWEA21owh4YG2V9fSjxsO
Vdz158h7prujFh1ZkbILJgWZGMVEMRnP0MEloDv4plGSDZ98i0FdlFsVf1G9IH+03AKBzX+nkeK7
8RCZlsaq247OTK1HrYXdv9suRN24+03H77rqtzr6bflJwX5NG8IHxmg1ApO1mPvHQG4ebZO6RqK6
mhEqxpynvHjBe3oic8e4Jv0VnP/zhOl88+Yg4zpG+5m+EJ8+CouOKW217LUqfuCgkbHnsKj5ZDFC
BVHGorQy1g9OgP9rqx7LsNRSC5kpPUnyd/svIXcWumoo06In71b7tbciXihl6wuy/Io7lVflh8IW
cAaVhrQKrzuYY6lmLyn5lTT/QHsnTRLW1NZ636tOc4V+UrianeJG+71AkpPZop1CE03T0UajrrJz
0yHnXIQm4VxZMQ2DN7yK4AG9ux83AWkLC4CcHfXJ0v0J6PQ0bQwNYHLG5OdcjJ5gDqs24gd8EZeT
sQCjlLZV2KE/Kl+urLrUF2wDfs4iVufe6wN0iUBPDrajilIATc7kvomgiftj+e21Bthgn7dNhywC
FeIe4GvtTChcfnFebx+s1nHJjs9LcpkitWU8anJRdpG2L5U1KS6FkTrZ9S0ylbr1o1vddsdFMUoJ
4cHu6oRTlDk/0n02atXh/Q7HrNhmJn5wBVvmUDugTuomLECxHyullgxJWPG0XO926EYmeuU8p5mN
k1GEuI82wQR8wLMgyBZVCUM49RSIIBcVR6AJBMmhfbNU0JHUHDqpbsl7ZpHeHAIQOUv5x7nqucRX
aNcHARrJ5JI5qa4lruqN4BxKs3C6kiv5mJSX87LCJS202bWVQxl9x+Uwl5ALlvIHy0iFSFi8OlMi
o23Mj5Yu+bvLPyQP3AewYzIHFKXhCQ9JCBoG+UZkS7mDVMVFqF3E/Bn7wxsPryWWr1/LoQM4TiOV
hSqnwmq9cTeQ/8Uy5cuP4u7o+WJHRD0WzcHpqMtFC23+TanpQ0eaXy5/VhsngkxTfRs2psrUEQ79
0jqZiyxSpWknDTs6xO27zfI/VX2FMxFhV61rDHx6dMp6eooiF3fAJnFOKjeNAqSWXc3vxt5j1895
jkfKoGtFx5rYyTXN9l2FfQBg63j8FIWDRP14diV0VbRdqwiNvzoW26P2pcOsDWDl8HBQKzlp43iC
gm01pUZQxnz5UgySgRenLcVAx8+uVHOgEqThSQ1m21qQhUjv+MkN2tp4xJ8Qlgmf5+Z0opOmvuYS
ptuGVF/qFfdfhSYkivuoJYB7/LOjw/82fK67I7ZCdDysZdLFSOlICbbgAS5wsxX1wo9Okv7APTv0
IvX2hiD0vuRFSD/4i9WFALrxvi9F8eY1iIwfVw9bDMGBxxQllg83IoYvkKbYu9p3EpGJ5dAlEaic
x1X7lWpxsRSAsSajVSJnIaQRxE4ib4vZrl5EtCJCWLqisupxWwWPF/Q+M4JkzN+Umq8iXFKHr7vu
vN9E5Ls5fAzLfvbgQUpE2PoZ5HNAJslbsNtgSiHKyugrDkTUFiPvIRVh8z8MZr7CHjmfaWDcQi+H
4yQ1MmMTAVVMF2JPfpZG6rZLT/V6wBSjEnLwiiVn/54SkXODCK/Vs5DMfEf7bgz5/vJZA+lQGMNx
8MbU687uD9/WedSg6GTs0UjFDt9oHw4BA0/OdpcwL/3onBAGmTy5xm924OIQx//2eo55xiXSRfKx
1OokCxsZcfbeuRVwTIxpTgEsB+/ikcSCeoV5DPBwgtW2KprAzOb9eQFhR4Adpvria5T90GZi8m7/
mN9pn798M9wjHbWTwj+MEn2mr+grs2wutE87jqjCQTcLMdrumUsJMJIaZVXBV3p/+VBorBSBynQb
W7G0QYJ1TKysKUIOx6Ae79rboBXW0r61JOaY61dRHzxRrKDv1absHxjbkNcCRwP0HQRozao8tog6
sIkWvDF1q2J1IVfUcFm6ulx26J7v3Pb7n+iK9brp4Lnxl/8f0CnbhqWPrHNRs019Oupv1s9sFWPh
24AyRpA+V20lSvxRWWzJi6owH8e9xVBWeuTmpOjZS5tXvZ4z4X5JVR+cI3aBPAUq0FTxx43HX37I
+Ap4n30OgUuZAXX1pQlh88cHgdggX60/0f6e5ZoMhEbtk29Z/s8JbWc/IhpplcLGGPngilmi7BJb
PEJwXrQ4xhm84CyNwBOEe24BLmcZsDplT6lXsLNJQKrss1wT8dgYMQ9SfNVT2ZhErUpUGVzd7zb7
eVqssNslHO5lbxrzdqsrGA5aFV85hJlKP9rbMp2IprBooF1ICtpQmJ3bkjKR6hFi6vOE3wryiuxU
y+RzULuWTAzmRpJ8TDVSHXPW/0D+4tjApUD42rnTNi1nj8Jpo6m7xBsoCOuZczZ3Ce5NFKqsX/EB
6KHKNIlqWjN9vKcnOXzaBv2owHyEEwOBbYTf+SzaQdMzZycIFNwWnUr+AxV6Ifps2CCGtesAA46T
dXc3JARF6ISSG31rWaEBvcQlkavczXUTfQ4O6FP3tlRVAhXP3e+qxB+2C0Lt0gPzt2sLmhq6L5m3
XW/SmRL2ujNQqSeDkFMeZnwAi02M692YspXW8l+xyYzVFs/K795IWgHnd3jh3rlQCUMZxOFCrrcw
2+E10i32kWuiPzTK/9cd70ibCfm6RDwhLaFzHTwd0wAwyRTpX+ht0t0d1VK+rb4zMwKN0DoeB7/D
cltNm72vWfCPMSLExdJVTBkq0SxSlRtPIy3hLEeVvC1X/8ogYzek7wA8BO5EMs/yckuhxw1VBJO1
oCzKkEm0yGyyG8abkPW06ULbCK7qmc5tk3uA7kd5gikoq0dpgJ8i/cP+YAvQi29ae1TI+EO2iOhe
k+x2XA9DHmrXDCiltR8RnZJYUGaS3K5soa/IZr8d48fxNfKY9nvjkMyGY5EH4oZyol5aSWtnIZtq
ukxdVntVnvf/6FTW1UdNsl+K0lILHHbI0CvwUE9yD75IsKgAM7VunKQmVr99QG5LhkgcMUUkSl3S
vnAJ2F+6vRN0JncU09htAJbKuKpCA2PGIxKhKDAPBnSk18u4IB2fRj0rowy85+G1IhBKeZUuJ2QY
wAYeJ3JhzafmVBa199OCcwWOrTA7otMonIgKAgRuNfur9uu7Au3IOHeyZQPYQy4rGYO8V6UP66Fs
9X7h8nYC+azfA93DMUp31RyofGkMqoSYqLDhYtxJqcRmhE6JQpwXx/YWdeq405TE6EBjIj+IS52u
UxYNEPZjwiFoQz5JuBT0hnlewERmTrk8wRGeH6Lzl3zV0I38LgGl3bJildDW1kVhXNX7aEGsCELi
Ff6QyfOb/6ArQ7Do/nEWJYGwuuFB5gj88vymTLH2ATnpATea085L9kXGlHSu19kWaG+C7n77JWCf
XZv/5e0uSHU8ulsTagDqWfTR8cOuWVrrO4On2EUN2RW6OG7Nb44BgGxOk7dN/uPvbxfnvlhTdrA2
38ATW7z6f1oW0mFZmpVOB3z863CAw5YQlbSMShNviqkIMCo4wZQPVCaqdEPg7ayv43QOtNrVJV85
S/nZ0XTKF/Z8XZcBd7A9Cq0oSMRS2vFUVPsmnbET/KUSFuTrhYiGtPMr20PYO0XYy1kapSXXhEIJ
N6tqb2OFwIXo7Rt1laNrKsudqG5qpyIghmbpZbDwDcypGw8rDEjF/VHVf2dlR5g53vGsQe4UwHkJ
76Qq0w2XJ8doqJjyfuSFFwa7s3+un46A7rJKM21EQZg4q3iXMKmXyPp3XE+2MZlOF9f2sRLSH615
Z7Ufv7BvPiRQWeQ9jDBKec0mQMNydlakB7lF2ZJSqe1xEgZ2WUHcWnPaKUxa
`protect end_protected
