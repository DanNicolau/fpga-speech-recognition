`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jw7IfBfWXP9eJDuWU0e38PqfKe0/Jc1vUm6Z2b7ajxwBXhYgiI+Sz2foSjstQTL6xNNGBaM9nbim
6poWjyrHtw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
s+ibrI1raLRoUd2rXujunmHZHYRqHyC6q6xfhfuYkCLERtM0bmMep7gZs/8XI5Je4ANgDCpydZsl
U28Jfc0S8MV4djEWWBFSAlmKeVRGHBWP0LpLNnTTuYUvZkaVNH66fUun+nY+m3upFmoNMSAbShNc
YQqOatcoaTDzwQfL/7c=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QiAvcnf7YYAw7dHZozDUG6Ouaoy5K/7e2VMEuxSyozq3yCbqzgEJkfTYif1wYAerTxFjLelgOz/P
fIUF6c8qwZ6cG1hho4cCbznyjNbbhgFBcr7pVdhm8u5bsPHRhGGZt1OTdziWmQ03rVaNWt/E+xAK
2tpmylpBpvIlXpBV04KIuEyJFGltH4fDaDNLvXjl4dNOCIDp3AOl6AfseOtvrB8PvAnkxNd7GIFT
zW1SCUM4CqhOnDhmNOg4zg6KLwam4O7m2ijAsioJCKD+ccys56O1pvSwdkohzNTXBwY7OK+LoUIc
bmvY6hJ7xCXDzqzYm1sgri8TY/KD+geiq9hfcQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aOi2FDycSQnhCy3ODFks+ZP4sdvIEAHLmaXZ7GX6mvs6Q6ZTP4ZEJR3WCJAJdhwPXcG7q0+QWmE7
OGotW/RcGV2M5tC1E65qLW2Mi6S5XvsJmvZPwyGzIrA66vbbJMkruy+HNo1TM6vtP3glUekw1WQ6
SVwilyGWWOTRb4Ai91GN5zQJ9kFJLYAfkaqm2iAfFiS784EXZNqzOO0iJUcN+0xpVigWMd/5rB07
Ey+kA+Y9ZBT/y86WyZz2U+z2/IbpZp3gery97Did3kknQ4ixUCkIBDQfa4f4Wx79ACBwKSz/p17u
hSXxgT/kqjqTlc2LLJ9Nvk6PjMEoX8rzknDG6w==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DENbXRqduWuu3V2gTVP0xpp6dnSko/i3HgA+Nyzh27hQybmHkq1WuSXw8LBXvWbOSmxHnowUJ+hG
9kbuLMpQiIkX5fHrTF++zOQKitTetTsvtvcn0ZWTvMpPiPiDdwGEoFAFw2K2n9CiC9in0iUS2ZD5
8Q66v03bZixgVh5tCfPzAzbSUgjAqmKoFyIcvttZaO0aGfQE1GwV6nM20DbNTK4GSo+9onQTHxqa
aQQPTSUQhG7DUSHKGE+pTKlG+lvItMYU2Y07wDjl+kZ8YqLXNhKqD/Kb53swOrFYAQjTiPo592+b
WfgVmkXQoTRIXGgdSA+zqD8acik/NsnRte5eWQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kHR+7qlDSuLko/NNQy41ELFqgqVFFphzjLA6veGbrz6ycAST3f1QKZfFayNpXMzI7kUNiL/8+3mk
/pXMZj88f1JdFIx8bja8PWtg/JTTbhFr8Jq/SqnMJBF83+t4nXFchuBK9L6cQj14+bG/SOd1Mynr
W2VnhoAFoGpk11Mr2Vs=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hfo/epns40sgO7Cvs0UsIdTROh12zhQ5gNuynvZLBmdb3Fj2rN+hjVOeLIQMZ6xqAiRwNwirFQo7
QDMDslVp7PTlXsYuM2jmZGPNzRCZfVWDr5l4NURNe7vv+zaditiUsyzN941Bed/CT5r5m1E8wowt
0WkPeUqYkDYBIX163OvLeS8HEksQbEm+pb/XdOOdEcvNuEwkbV9S1cIQ93MQ5Czq7dJaIcuVbRg5
ZREQKnqDtzNvPj4QqQhMBZtme9o1Voyl3vz3END29y/Kq1YUmKItCbeoRwdKRlscV1hSdx6D47dd
9bg7O181GuhZAuWNF3OTsxjC92lWHGw3WXKRsw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 681248)
`protect data_block
bqvrpHTMpS0eIKgBBO3joXpcXHb/zihEdb1XbtdaXqmMfsgRH0Tk3P0iaie3i8det2caS94J7fXv
/0voqKoLD+rekmzzuKTbtJ4Moq46N7TTbWGGs8zAaWFstZJ4WYMPAZbY3XD62SQcnub3hee4adv+
qSpBlA7v8RVxudGCYwlmvxw5bkv56HUVS/Zsi0bTW3PZy2aESrxIWGfWyxzSnalxaR9nn76Mwh29
vFKdXkAhgZMv8et2Ga1U9yKV2bpNbQaU73eOWllDVMXyVHrdiwZWag1RNtOTzIdPBms+eDijvU9y
wvQ69fPMCaQjQ/alisXIzfClWO2Y1sEyiat7cX90hcFMPEBjRnsftIimpJQk3ZNXQgYJ9GYDpd5N
2eOtvlv0tNaayoIJWKFbkF5Gy8M9/UkQY7geApnE1JZtcSQEjO+Qh8aOPigP4eVH+mQHgCZseIj+
6Euh0JjrOb6fptCOS7dtApfAun8f0QmisRzL8EU/Hd+4cZ/p++7NzOh+T5lT/WHbuMIDq69bs+HB
qAjGg4Ce9BsIfdll5SeiwVXqBdFJisooTsgLhcIkrki1WfkDUdf7Clh+FnQbSYXKZal6pZwV2lzF
5VMEgGCc7hgLaH9KyOF6P8gw/9HVIVo4a7HH26FJgep0UfKtZdFN5AaUO7fnDN5U04tdL2FLYKZc
DPqVx/q4ymVPcGAU7FxQmN61cMTIQ+Inn7rUtrMDybUn0QxNsoemSqEgvSmR0Qjt2etRDgD40Qy2
xP0KdfNMyk/pc90s14OeYP0lqn0WhE8V7i2NEKwVPizLH2l6FG9nf9Zh+Zm7joZth6HqP4UKO5Tc
2UtUtS1JgJmLzpaEwDCsGqYshYfCTPWOOHvEwymqGHrydvFTZAYfRRiwJPkYl6j1ufo+KWHIFofe
l8kQtAkaUIkVltKLYoe4RRnlSDX+4roZCCNFSUF0AUDRL3iJ/Ps3M2WDeYiFr2AvoKInYiCssgog
CMVdFZuClPb0Lw9gyH59kHvzHzvt4jHjP9hJ4ZIa9ZGW0QoBw+0ur7YPzz9cYFQ1+EM8xoOrun6Z
06SmVUBu2aYV9QE30PMfgBc+mPeFY3L3j3dj9noY6XaGeL6+vqItAxUxib7dRsz6mKCnI0f356sK
gWGUv21q5NCQ3GQXXv5vlpNVDTVOmEcadY+GXeXhltMnLI/gkQtpwSf1MlRdbvg2XA8xVvAdCV9o
A4yO9eifsH7DUOMnyZIdZax/EHJKzlOQuKC8za7h0ti7Spr00AtrDyRnWYa0Unp0Pkkpwc+DNN/d
gPuBPn1BYSsURPm5YIicozdZRSGGU3aNFkvgnGPexUNp82OFzwP0h+DZ1zcFky+mAnk9YekEV1Fs
x8JyRp2lI9SDVYp182FKT2gaA9kuWsnJ8Rme1WryRfeKkQiIvIeCwmaPVJdQI1+tSMvOIjgmRrbK
ucFttM8VLBw1py7dxQ5nLUiQMkya8EFAKFMDEjAc8EFPdGP5JtBLE9RTBnPXrudiFC3KRqxBZi1K
z1tbTe4DNCOzIvfEvv44tZcYm1s5L3DT19bDpHMmP5cYey7YtiQ1Fy5AYvzgmUVIp525tKckjXpF
oEXDvSlwzRNPr8s6/tV7eW8dJad6BkEpSHvHbfKxSHFk4F/1jv3RiYTbd3VLtpijWrnB47KCtm1x
wCVUJIUfel4NpZnGRiaRYozxcItlPbCfkd7VqUsWPj9S1rPVQOdYoc0bs39MB1SIVRdcG4KZmrxR
OvDm2j+0x03R0l3cFQNL2UhJoEjRl4EuGVVK370IpVIweU4NHB6A5VzXW2mT2Nb7kLCdWrv4bEnO
hD40icf0ck6SRyFlQ6EXT2628zL5WdzflS/4c/O0aRhG23P8C88KoDkUz2J1PCjpl1+PFYRnNQPe
fADIYAGtrTkyPgmhfJa9k67bO4KWc25Dk50HWTnAdKwbFKJPHLVezzqQGRgUSQTZTbsVLooCWO2l
vib9HU73a8VBhPmZ50Wk+Wcekz+SpZOxGtmcLakALf/Z9Oa2/+OR0jwCPW5aZvOXEKbUxE0w0yAr
uUJUNDoy6/ME3dygQ6rQ3yXvHsZWV1aTwzrU5r2h1AnctSxMz6A0aaAnO0TTpprSkRY41QjH+T9w
gImDenTuWrp5mtixV62zJcaK+EAF+MlMdIMgOBSap2UFXOdjWq7/5+b5rVQ/KfhKa7GAgy2Cv+Pd
a6fBIXd7Fd8xP16+uXRaU9WrlFj+W9s7EMhY5Dq/zF7ShN99qDaRuRV9l2MbBIKlQqm90rCLbD4B
PwGAHyPJGQBT3zzQbFSlMU66MhWyhZNCchu7ws9efb27ReLO2FxtTG7KrTCwiaymopslin2HMltF
w4CeLtn15/Y9jYzEwMrMnxo5gh9Xqq1opp7VWpisDg1HyV1Cbw03aFlqTT7z2UdjTL+pf8ijkCDq
Pppwjess1fou2VBNG5wUao+BXW+VFjt7mT1ZXMZmMHHWQBuBe832V5qQFs4CoMPMAaRkwaiZRlFp
J3wgWvbDowidtOkBcKtwqLiCy65IrBTnb0XL7t4t+l2OKwAJvUk5p1cYAgUQW6xXBrGgZGzWUt9W
j65uxpcjPQDyBpXb3Y8XMTW+SnpDzEvCfpjoHzsXmIfc0OVfoFKiYMYlwNY//XPMdXkxOSGYSpxm
c/Z4IcYez/I4gj17B0d+y4n9J0IPkx/1xQ2MOu2D94EHMCnhOGRix7fq7/LQmD479H0XLhwWjtG9
7Udp2N4NxGDKqIgf9kTHUA3pC+c3qGnw4VMzbxQ3KxqmwDYzqrOf517b34TfqbUy1f6w6rJgiRVY
Ku4RdN2Pd+v0r7Bsq7MnTt4kQhq9kh/m1Tjx64W70YbnrEuP6ShNXgBPBM8rX0F5LZMvtlc03rhr
lmIyrON9cM7SKHfeACaLnzKP+Ic6Rish7Ewqbxckw2twF0zczAa9z76sKBUc512JCojg2PljQYQ+
BoAKmZwsCb2S9RB7ceoFz3yyVoRhameN+fS/IsPrLefp9+Yc9/rfuE1JhSPd2bIJFuQcNdJZaskR
G1M6FxvIXxnjngFZbDQD75HLmo1p0Xkm2hs0uU3/gU7LWT6U8jIXklUlKwEjrvmcNbL8L7O8knek
LgUa5NlWcZlcOoSgi+OE+K4mWXFNr1vlW7HVGFML2zEwdbmDA0PFR7b0rmsex36tWAu1q/4yK4T6
wQR9/QfVht/sPmybNpeCPRj0mydtW3+QP2A5hKInW0qhHRxreDjsW1GNqrmHF9svHe9znebQtTUy
bTB3cU5khwziAr7FId+teknXmrhTxpMVh7rIuhxUCNc5qTigf9/wTBe+2p3hLmd8xcUCB1VG32lW
YyTjobsg8qmDXrpdoRlV/bUgQG0JuI0/9y9H8Y5iVtNYsjwPaJzn7r+89zYs2m1CgZjW+aAgK95y
DHA6+qSKIBtndkPUXFY/xpVyrwQkr+uhSmeLf1+aBhP2KdBsnRsRybTgQSJddn2OGEKqvyDd1p3N
7qRFU5hy+0nB8yGWSn5X7eTn0UAKeqHJDbZCFWdms7CynKAvrn/vVxRsD8EKbTYk4c4ArTh3DFiJ
Tn33Z302yqn+Jda0tsAql8evdOQ1lXM3KGA9bTyF19mwu884OpF1ttXQUV2rMkxMChWOa92vVIKN
DyBG7wWzmFkGohYuNVgRZ63jQNSUzb5TJ7P7fUMH8n3+sDlIB3r6Rb13qU86Xz3iVxGJYdK3R8/W
trVuv8ZdUwsxUBqWnwFhCpct7VHfp7Wz57LqXO+bJUqthPdjSJwlGZW+FwKTbKQoUO2hUpRaG8+i
nVtMBuxrzja24RXRoLo/CVxVpuJIOiIwyetuVdoB1dOl+hPUf+xC5oW0jWGIWtLIH/68iBF3AGsM
wcdNP+e9hCYiFqdH+/pfbYTSAexF8ztvcUS6MSn5sVWPWpnnGLE3HjE+6eYkcw5wGhqUwPw+Ucvq
KlgF4lA5esy3ulfDb9rB0ZGJHkGlbxr4VCAJLk1Xl1a0PBKpYKwCBLe5jA6cF9Qb3fyVRvqw57cQ
4HupQ+Y5R7zmnS6qOSGZKUfRBZj9y5SBmTMOqT107HYA3P5S9Ga44GrUMQnJOK9eAKsSczNl70Ub
hMnI+7gplwiMXhYg3+W2PGNq30Lx8oLc8Uw6hJcEuGgUHep4KcnkQ9g/Tp+ZMyY2nwS2POLA45Rj
e+ut6nMttuH27/+vqMz6s01YO1t0zkFeqBYjFzXX4Bv65TyATl0uiH6g5D4ZmV58gUBysuqRAEpq
rRM9hyTE0p5KzyJNc812F+0BAi1/wlIeww+ry0xj+OFqlN+1EMluDHoikAyZ5dOQTFk4w6U6BpxU
pu5o+eupn9hgJ/uXRpLXojqaB/e85nHZ9Hp/7IFCAv39ZHuqnQd0iLjwfIQc7PWV5ueGKxvxM1V3
EGggwSpiX8dQbAWa8IAAn4BBX+bBF8X4oqyvFgTPJ7HPqc9rDPGEdOi/L0L+VXppo1qcfcuoxhVE
o9T7+l8ajyjhyT/4R8bcGWqLQCoUTJ7gT055xIq0PWXeVudfAeQ6o/0E2FOHD1+Rud9W6Kj5vYut
piGN+yC4r4QsbWRWOhB+bS7dLtVNbOBlAgDDLoY8CRi05i0EkxgEstGyXXNqWgJnVjSUS15Bk1lE
eHw6C43tYtTMNJn6cboW9Y3j/W9yknuHRRvvspwcKVHUAA6vS3doMw6rdzD72FDQ06ZIvDK2VjZH
IHt6TLHJgZwzzhVczegmufx80Ff7mUQ4z0PH72kOj9U9gGfbAAP2dUnNzEeTBxXnBN4pV0L7PW6m
yOfPJ/6sxbLAk6GFpA3aiKcJt99uCucS8LpAu9NmYlLBY4UGiRmHjql6G/wR/pJlrpMQ5UO8xUxo
ZVbGa6ePig9MHJRTe+duNMCVkHrkm6qh+cyrB33MsuX1wAyMe9uJ6qp6XuW9XlyxPtu6SpRyMlsD
Puvd+DEG2xT6CVaFbfKt0j4/NHb/XE1EOg8r6vKo7/9II+ZspoY12RknvwMkI9MxXDFgUzseAgOo
NYN6JUkIrHDr5VW/60td5gP39DnKCIDhwwzVCQ28wSk5QxBkoRBHC0hDLA74yE2VqKLVuJ/MwuH8
6tMwuyOuJoVICCsKL2NvRR5Eg029Oh3fVjTJUdUXDkKd3/vTdwkNk5zHTX9+2r563wOCBpWCmAWE
4fZwa42piLzG39EJK/G0P0GKMUPqOFAP4fWC8I539SV1j0USmlU5PRL8hVjS/AdR2i2XmHcAGxkx
4u/3y+6FF9S4T+xsRzclXmGRAaW1TAP33ffS2++U+FcXwAnLiqs/SVGCg8DZG6nGASbH+2YqzAln
pG75QX1v87KQ5QIbxWVPNEHL8mJIQqiZVy2xXXaI7arAgB+P2HoHbh8evPx4yAe1TB0rP4hPW4dJ
Mmgt5QpOyns6DqkkjxorMCb0A3aVB3TocbX/S+kHAqQw2YcAYT83DuZMvgFD9LUiQCY8Xbyx/NiU
5ZG8Nm51fgSPz/XFXqdM0XUbHu5jLpr9ZBGC3oaG6mrobEyfrktTZqo1N9roA8wykPChJLDdvs6S
hpKheEmdgNDIFFb22z8vdTFu/ICJoNkXevBu4oxj0F+iRDKs/z3RymAW/NDqI1pcXIl4fh9VPYqs
QrUeJI1EjPV+ItTnioWy+D5ZDOQaK8EO92RZ/X8k3K9iA5oiYRlY1RS4C9Cb5HflfNv9EVPDne4+
5fEnYk+XLBGEyZgFCivaGS3oEbpJzw33qyQXqAyHREEALXchxxz+fgAFZaiCvU/taBfAKwqN3OJz
5DZNG5u8CAbEUqhZqHf3ZH0rQ2R5JswhlQbA5GeKDB30N9ZKijnK3RGuPqLfQbW8tnNCIXN7lsUp
pN8UAAJMFF1Ziww2kKKpRCJqqAlSL9i82CjK9Y44AS7MPmJjl8CGngWGqn9Jx9a4t0Vxl98z15Ug
AK0AZexmI/mC2tEidgWaGlgg36eF4Y/RAxnzLHZZbP5sE8oowj/VL6BFf763eval1RMxmWZjIXgV
ocIxR/cEZ597Bx8Pzxln7xdmiIqVQVs6KHTzz3bl/RwocC+IEWcd5/9oCQeHbcWlGLpibPXb36bo
iojwo2+tCoPdo6zVeNlHvOfwItM5l7sDUs84xT+yO8eCknDDha9RPGud8dmaCnTUKL7NAoVhywrS
zoxY1MEpn3VyBOIthAnUlM1MIo88CVHfdV+dI2uTbO8M/gY2uMrRaJ0gZDjENOn7xQjh3P13TY4k
F8VDBztAjT9nD8libqAb/u2GRxVFTISdVUqwK1qwonoMf5KKMYnHqKfcelVjqXrBo7UAAAUPFew4
TdeZQMllAkBZRovUJ4QW/z8S0XWbuv759J0Axcme10Y3JFWCE/gwLc+2Yf6xDtaUQO0dR84utar3
uZrRVr5zZYMXj6b/oZ0wyKXVAMBQ3z2upV5bZF9ubn5veutn19e7H8ik1mdbquUdygWw2EJSlCs0
/msTlVfMwJk1daskX22SkGGlKVshVHdUTHC+A3pdJD1P7JL45ZRNey6qq7sixzD5fOzCJ7v9VdvC
LKVP5FlYlzcMcbf2d4iBhAauyq5rXkx3LMMkr++orgh3jNao0MqIl5rTA0GnqDVY1DG6LpD2i6RB
xmbfAxbKhdRwOdC/JSPME0lMJvYJsQXoYHrIqWpecWIuZTLS6uSBfGRHZj5zjJo5jNaPTPqAdNcB
WutpTDjmOKeRtM05BDNGx81YutM+tRiDh9APd9vnKLUqUXXt9h6+2BxwXZutP6fhMAA0suDA+Rvv
qB1y2JpR3wI7x3Xr3K5XMJkn8At5tq9+y6v/ptSmfRYpBzGLtpTsqz+MZnkPPO3jxhA5HJeaWWkY
QHXM7BFRWaCWdQNVZgirSeMigCP1KcCI8SUrYNC5rsw3UZ7Z7H+SeU8VnffN9xy9YxU+OX/MkW5N
g9WA9WkAaKJ5v58dbSHlXX7s8v4hU3FWcx3Pz4BZVu1anjtsZUTkThIm0iR4DItJifKp80DP9jqb
xcrKT+kO+bfo6tBpW9+R794G8KEsrhVgsEplZ0pz9vRtXNh1WbEV31Qe9BcovS1giEQ1WScjyI8a
n1gyDowWLmNO9r36sb2EG/jIhxy+B4cmPUXp9nVKEJ8udufBcqm3O/EkwRtkUeXQ+BoqIhTtZg18
4ktBzMk+WUVdZ7r1CMIcHgwTfUx/0D5GMi7dL7n5CNP8a1TWfE7lNPkX1nWYRzqRAEOfZXAaXh1g
3whvf6msqCoxm/LCT9Kzk8NkX0ZUsM0LgNk+r0oWwNP+gQojrmOxD+8z8K1ItsLW9opTvvtAyHDV
IRoONpTzDVmxs4/POHEC9g75metRzpK8X8uI+veE7OAGJbES0GxSuo4DVBSNrduVlq3BHfUAkU/t
a8JnkJ1qHWAUfvsBQPjv9iyTUzXTBh5L8PtCKgqWSAIFvhy4zIbX06JTsBqLVj873BKgyJ7xUxwp
15C23Vu8u+WavO/nV8qna0SoaN/NFnQORRflED6ZmlFMh3wS/jGBB096YqQi9TZJOWGxy381Y1A2
qa/nvMuBM3Z77GrHgJkyXY3Ac62ZUD4j0OIwuvkC+qPyPXDjUjikDUZOPhZNpmmsqDDz87ixdw+l
bzJOHDf+fRy865u5hMWUY7DPgmjw6h1RzL5GDeIgzEpeZJv18Ggx5rHAXZxmMwKWyzowT6bNtOr7
RQ5Q0aTAFN1/lNfpstwKoc+JUfGQk1oznyBhYHE2ZERA+Ro/1bC4Nx45S4Uo5QW2cGG0u/zE8hYp
f3iK2SVukA77BEGm78xzUZQF7Whin126UWofpeUgZ8URinJSxiGLrCRJTD5yrNIBMqX+CY765BCf
KQqIEYycm4x3mcA0qjV+tKPhHI9AIMHGWrW5duLeeg+92DwT8msoLfcfAuu8mUcC3GCgU2qxEVh8
1mHPk5TnMpAF9em3Ut6r+g2CjBAcmGuq7S5mKMkeyjVp5zW8YJJbVcdubOb+MUSBguOB7TuaUHfL
/mWdrHVJecpi3z7edH4CmkO3r2nBtrE4P0JFjsPGJP6LoCWvI4VTPwMX2/N8LiV7qudmkrMACdx6
H8ZQhVXiAR9Bb/FYII/7TTgBWmlGQ3p7anJyjVO5r5b8BWihqYaniGMnw851F8fqwg2QKt5NGHQh
Pi/ImgHbpx2PJ+sH8+1FSgSEQl6zCjAM2hPXz4yoOgZDIJQznC6IFlB9Uo/2v1XxQWjZnXFkhkkd
nTf5lxW6HUEJH9nthjDQyr4NBZ37S9gAoVwqBWIimcygQosNCwjcmuMxUPM3R+AqWfb9sVza40LO
eVGICH7p9VQFPQ05a7QaMq0QuuQK4Y2UhVh5gOFsXmcQHOyNnFTlZnIhBuORFsDogjihwu4XQzFk
BSCDJTKSPiMApwestdBNhWdF5yVEXBeGQ8OSdjzOGosC4JGBRPa+kaXprtGcBBSf4smlGSy0gP2O
ruewwDfq7DnLPsGv7dV8L545JJZTKPUPgTfoU2HnhGea+a/gdoXiQzBwN1Kvb/sGQPNczVIJ44Nf
KyWEoBwabCudJVyssYQLYp/i59f5FFt+8q2uuONgQeKfXV0RsK+790jfs6GKGyt+McogLVgujJBk
baV0SJIkpoASBaLcMEnxJvqb5KF5GhupJOkFWFlZ2XzuTGtx3E50BmxjNikuBY88tRAX5agGbHx8
5iDm0T72wgz4BQscuvrqJDFHG+w/UJK3YPZWGndSlvVlYKQJNTpqLV88fDxJZmFEIxbKaMmV6t9k
sgR0EBCFIxB/EfS8jXuNChS3ICeJbro4KtmHmJtzqN3nAab32tyY4vS41WFVpj7NU2eRciUj9Ord
CRjERLF91jmo5IWnzCfj7k7f3HYYiB2NAGG7WOT63bPjLWWGyVyosnhuoOsRvtShb3AzvomWCWAn
oPgTzDc3xkhbMYLW7IW1ubCoUiDMViNv7KbAtRUIiU78IX0yc2+sZm2Sy2M+M9DX93yp7CSFQ3q9
JecoKkmgH1H9N830hgkRHijfFUTDR/4fieihHwtzQ3YfB2iVOFUs+Zw1LNgouj9gvp4CcQUSuzf3
wlHGWVf4NMclOKXmrCagVRwN9MMvjxwJqq2nlMYQZBVsTJbw7PPYAV63STmUv8WAX6u+tsXW2t62
G/FvSJ2sb9BEqP7djnpeXHaaLGLpPB6a1ZnS8TgOGNl7d3ATGBXQY77obxesnG/REo0OKrP6wcaD
qtnC24+shbF5+aEwQbNlmX6QMs1Zsnn1A64Co3jtiuCx5oEhd1Vzk5XVKaojh8KmXdNJgbwUhain
ujxyiD9PpaxCO9wpMVYKb/9zvUEdrmXtu2IwdMW4cMLlkGFPFgdGm4pBl8N8cQYylkHWZeGT8ihf
ciquT//Eu9Ije87Boczrl0BKmKpEnZXhBXrfTLopvYPk9dvownMrcH/F4hTDo8h1RKAcAzwMO4D2
V6z5i+7MPS7UkAm5XqxEpr67IqB/8Tmyzm5WxJbCqWULbKJq2gWDUcnk1f6KvHBg66KumtYD/D/v
gTzFQzYaflbk5uS3L8DiJy0IzjroAlwt1TZNFEXWB6bXQunoLnZTJaqMGeJTGqMTIak3N1iNj3et
COyZgp5jlLnTiI6J877l/zUgM5P82ThV1peg+xDNPxdBUM96/F2jaNiB/G6drUxcJ8iVAPFGCZ03
GbX5lu/fquOCQFroHLY6OZxWlzco6IByDZ364EEpkw1G/0lUc7seD00oL6ExjUzWiceDwDfLHZYp
wdKO15x6Hk13kzF9khdqR/Xj5RcufmiBHqNjhICDyVujPxjM8qw2FXQERCBg1tnoSiO+tpB3N/Oy
qUOOLHaksL2qr/6Xm2dmiRO1tcSQd3lL9vhrQgTxx0qeQP3+DpqLLG5fVXccnaOWDiqXvz3JaUke
U4fUblznlU0yA5cMKTm7dEorGuVDa+yOmcdy8e/ZVip1T6ydIX8IGNeJRrU3I2EIuwXFNe5CoBEy
1Zy8q1+ayqIEnLqOz0XWZsrck3Gr/uyq7HcZhQ+xjb7igQGxdD0iE74GkE3LzkVLcgR1F8yqCC2/
CFFOQSApbOgsDNOmgzCD4+4BCUBpb712QfzsZPNbAljmduMZQy3FyMm1LS/SPcgthWQdLp6CWMt2
wPDnFNQkTOzd5ufL/4yBEk1o5buPxxHj2WwEPcx0//OlnoFh2bxcp143e1xedjgNDhXuw4mfo+QS
J61u1RSLHXHi0e2wCD3AzrChipnKu1AG55bVxGxEJGUJF+DjDKGD5odOYh7EeJ/wLkjg0S7df6rS
WlGDK4frDsDFkXUMlfEYEvvLqHXFWbuIWxs+7N+g3ajPrtuLcc3hF4Dp+bq1EAkxSRmd8m0MZCtu
uLR91w+JykxMLh3ctjBTwT4u9XXyfU5i6m2pPq+jbC1Vp6o9uTT2A44cyerfzuQ8XdYQbLvijvRT
yRwRQmQdphJYiboW3CJJ4UcNS1EPh6v9wsdFtyLx4tR6tvoMYed9DSEKKji35S4WXWumqGhuh5zS
22BYvV8rYgRrlT4aUU5MeV3Pg8BzkG0+AKV7wIej2zvRlxJsVmBiswXX7Qzg6e/+1b9wRH5NqW0Z
5fwYygT5UwGF/G7uvSbtXUGHCdDLnyk4O4zzOvkNrt3Vds1yzPUlXDwvJqFbCDcPEqPLeO1ze/7z
iDvEY7nQ6Rn6bPpDamyftV3R3x3aap8+kTHGc4BqrD4OBBnj3Tgk8XDB03T098xA0VFAwqBLguvp
I3HbXBuYCiWx2pmq1JMzzj5RDgzgNjDrQwfWt2Vws+nAJNGDe6FTXIb3fxJq5/d7Hj8rK/Y/y4bh
EZcPB+MKMye75v9s35hNNZzEYwr510n4oaevh18iu7lxe7wxfZyQcbofV7wM5L+xHA7vBjBuxU/N
85rYs3rod848pOMY9Cuq9RafoMBA8FDixJY2J5jT2LerpOWvAH79w6fJkcU+zFia/kG0jWgeEctq
oMWsyXCHy/Lt+JFIq1IE8XDNgAZ/hSYX/4ecH98y3i8RhmOqbmPCzSvKkQ+mi8l09e5HQTodEKPp
gCPfkIUJa3tBBIVHdI15LCTBkkSpfleQsuaYAPkMkFJ0Qto35Ushwo+kDqCe8gtsrNKWr3vlG2Pk
YIS3Z1N7Uiuxj6qwRq5uenKSo6/GDDf22xqJLLuHt2IA8BkBOjBi0mkZKlH0/Yc5qQjc+wbuVCNU
+rBNsDRf4ho/61xQ9ACeHHR2Uq1FWlLCKFdM4qs6W0e9f2jo69Ld8gsTkhzqv+0hP4Q+lWgUMueg
dI0AMwwpayyKzqEJ/EqJh7h3eOkseOOELNm6d9IeIEgV+aN5o99U7iEkss6z7dojYg4o+QS117aI
lpSs7weZ5xQc8Ncudol0xJ7s5zvVo9bg0NCw+yDQb4bd1yz5gdB26K6nTH4w3ezpOokOy/P2GIoC
2eqXkKNzwYMI/JG8F+F9kPD5AjvVDDCEEwml+U3EvvllHNOdC521qxqKIPXkS2cRZ9++1oGlRxrJ
pNhp80TRo9iILkxSkgF8F2U+FXbvl5i/h0vUjA5/eC2PGUCqRT/8NjHpluVtVdI1lKzFxpAsvd2j
Mh+4UFQCwkp/8wor0RuJqD479T35MdThOsQKUDudvs48iOb8EFKB6xEwZ7Anz47O54SoZ+VmlS2g
m4qQh9Zb9UKhtVVG4Ta1KJSf4MLwc/Lw0cuNul3UMv7v1r8CAsfQ8QVo6cDWzh9p9gtvy7Vb2JpD
MEleBG0AaGJgjQ1j3D0FXaMirSSBSCVaRJFe6lQkSNZxd0kdnlZyR0sktcdf1Sf40rxHqclvxxYv
FB7bGX5j2Fz69tX5kIVJ0XlY9nz3gVZaBtL03KGlttpX5dWIphe8paZLKSYR+O2B0AGMVgj1oAzA
S3bNbscV0GqNtMa10hlPo9VqE6Jffh/iYpP9elxTWwN5SOxDO76/p/3rumDKSWPm53AFzcAyfMYF
z+qln4eZMl/b7oiQSuxiqBUNRVzuVlWfnsDvg+CzatOhihQOwmDCRdZztsftJwpEsux7nGT8PNaF
mDxdBxLQJNDQtkTW6Y52PxS3PIfD7tKmqF3u31lzEvBE0pdd0dCcLV6UeoHg3BPTPWngxPv4vwc4
f1U7lgSZbTVAgjNweQC6jrn8p9t6miFFCQItn2IvzQTN+xxOPrq5h2VWSqqr0G33Y5AqWHntLeJn
Vx/ols53fVZTCwWghDDPy/QZXjA5K/0q1tTNByd1VFI6BsLKyclRkKV4SRz2B7MTePF8H6cmlm6q
25ka9eMOzZDValkCUPWpOQqOQN/FMZXILABPmj+rfY/XHmtzll3IcYRcqRK3Pedj5LsvoPeBbxVI
IrgD2/jwvEliW3wS+6MMBQVxD4jSFhtivUWCYOv0OBy7e1vnYgmYi7jnGnLGeL07MGAmwM6oZWRe
Pyztph2HXSXS/Vped8pw7XjBC+NJcEDvXIhMtLJ0ZESKZzr2HKbjWO49cWuNGnV7wWY75ThMemfE
pLVSEI2e3zaa/xfBN7CautBNyauPRMsFPJDt4ZgU+OXwutjWSf4SdkDpDAEsFhyUD946YGDSgkpD
XBfggbTe3QbW84l9FkNcYm2/vz9VklRT+w7FvRn9JP/YUPOcXuJiAG6hbX/KaPfbj+EOvp4dttrt
RX/Q0O2ul8vvPMt4sBn2diPV/xd/kHBg1+m7clepQSIpFnO7TtTQABJZ2mMMKZtGj/922t1lQjPk
tB33cg+8NjdMmFVwopipTzX/F2Hy2NDaqVXjaAXqN+d5IaW+q6oA3g6qJLLHh4msTsY5Rz0zbTgD
1knjJtkbcwxKuUd0Rr69b1b1nVFhUiaCDHIF4ENx8zB7asnO2uBZdQYzEdNolgPDWQU0eZvbVkXN
mTbJHKsqy7X579WMaWDeazey4jTkwwHLDHRpr30pg0FB+Ka7+Zx1UPlauamMo5SVHRYheBid4prP
2Cch+t8rInttq9Imu5t3YEMy7YArrnzpuPwioK8BwAZQPfVgA9HcvpiyohyyOFWXBjGRvQFEAUP6
cPk7OVwhOSK5kGI+zzee0/K0wGwrzT4ARy5ohfE9lTu+TQPArH2sC4aihAtrGS+x5EcolHLe3g04
VHO5PAwEo52gOBXEgo2FKu99yk8Pco4JqPtj0k4EnJcSWh9ZY/6g6mIb5Ry5JnHFX+icsIhsMvlz
/sOdNVNE+l2yMs2Fa7E3QVsDMpKuC6r1C7jVuJxZLEXfynUu0NQYGr/eIQV0Noqq2slcrZZ43Dz/
c07NncUt25Ow/GQ1tq3a2h1qkn0AAT1Fq+1ohlVKfSnGl8/HeRrSeqPrAjk356mJb6wT2DoHkeF4
1uDQ12OWSjBsGRv/mW+p5LVudTvDka9cDKWSGHjFSL+VBEh5lqZ/vf9h/Ea57E5HT+Tx0v+ekUw6
QZG5CcUQUcBJsue2/TTypNLt4ik+GeYL8iqQukHBYExKhTyNddyhru7R8tUVGbpM/phgYAnYePuV
RZ1wPwRCgFqaq6a2nOrEi6y2vnmLGLnX1eMZXwT1xaTHwgE7v50dynggAWSGw1UIRtlWJqnQn/io
bE/GTyH76GWcYF9CiWWnpa7jMZYWEn88YkBRxNLLFiom7WmGbgzfVXT1ZmSV6RPfW661+8DlXJLx
LHBANG4T1s3XtzTGjwZyZhs4IU5nN1tdpARCZ8l9SqfwU8BrszYVpCswmRD5HDSk3jSSyIk647Xj
iLEdOFn9LxlirWyw/vdkUTm+fCmaPSiUXrx92kh6QiZiXQRk72GhXrARVafBUNw5kHk/How0MQeG
XxohWGM1VKEO6lojYfdlnjmvgZcrwUAvqq25/9a35hcjwZ8ueMmVpQgWY+BV/Ul1C0v9cwPJsq4e
ShA/SrON4HiUVEY2ysx4bKCsZETFTnJftdy+9z3/tVw9OFD+UUAY+X9wUdoPRwemFiiLhUjfS1uM
DvJIxC6BM9TVV4NtYJeaPUBuwpx+twA3qpYpAeNZNU9OR/1+R8g4uFg0OTiX11t6d9CfwJc7jRMD
7Ig9Xq2Cq7sha4V0w+RaNz7PDxXGMzoD0Urp8cWN0iOAbtD54CK5agmpYS9IlOQy5N9DT7pw1GYj
lGtRv0FPbcOZl45z5SIk4MtYTCkVm/9CxK1zvVQWPc/IXR8UN/sWSsY7FRibwobGr7hVx46qFY5R
Cz2jy054HHY4p8OX4K8bft67qjrtxy1VENniDAHA5ewVDuiziZ+i04UUllV806lkn1u5fGc1hRAP
zC0S0+t4Yap6wMHUq762w3G5slCflzTwFvLOOXiS/n2N7drX1FTrMcP0fm25iM2f2yVEMjHUxrRj
uMNy7DKKHP6Bk4tZvifyyN75dzfT5nxUt43vG8QuBZYTCVtc/M7461nmstYuNGMu/jcCb3imEdQo
em4oIpMBEAn7HPITEsa+JqNrjqao3Bc0/uf4In67sc9d9KbKtBl4q+8LgvcBEXySQTfDdunyegsv
+ljBNohWScEesoW3lksX8fN0hTtFZT7K19XnbcR0th3Rmfbn7rlws4ogSw2YBvJjlQZRD3a7GQqU
GuGPp2OsTOt2v62U/PjTsAogVshTiydRZH3CGIBEEs2QHblzEjPyf9qVF0N4YtW28UrKP3Pr+0zu
Lm5VQ5BMOMmODCTD5hXiGSOfOJJgrtaLhM2ehjnY4YNZctZG9yDZ7Iu+i/wuWl8NFhI44eMWK4kO
o+UNHfhMppzhlVTdEwo904IP+CmPbvrHSQRIvxQta46pH1npwjmIZDc9zwYqphAxaQ0R1MoK6Uw5
vTC/BxbL0Mxitu2uAk1H53Y6Rx73WS2ifrR3Ys17XN4eJKpEFlsbbu/95VvT/0i+6R9vP1lfLR1f
VsTyBow9gHC6kEABu0plOBHtOBloNvSCm7z1ThBGacks/o/7/5rhXmDm+bGeZDaJbu2465qb5qiZ
lKIA9loQBonKXq8phjlGDieOc33Yhbg7IOmGJZYxdQX7BpKakTse6AB60g+jSvGGgEKLHJ0LxEAi
v3VBMyrWu3HzvnBj4IaAl1CCoRm5GoLtALgRsgRXW1NL92nxhkwRfxhHP/kudk+NmoB49asNhTVT
1QEiDcu4PLJG9GwUafB4cpBoraNAO1l/nQI3ESWlyKbeS+FLnbxf5QBg/QAsC1rQ3ER/QjePjrh9
Ci5q7K4L4ZKGvBDJ7XMfwPdpZw96DeTmVKq8BExFSM47cXLU2DfHsOvRGR3htSkdXoX3AxaRoDwA
H4mMTRquziM+tD/R5IlOr9eKBob0Q007cEBI5nXEh7Agc2m/MtgQg67lhmLTumIQG0cRMTXOjyRB
rfrnsOaT103XmWMVu/1R70+Xg9UATjEwPReQOb5HpcW8XjvasA0EIIUYxmiqt282h7g3YNELLsBU
R/kiBQJm+lA4LzBA+EAKGDB1xNUbcCFny7auo8MTDjAw5KChcpxT5nIv6QMIY4vFhz7YKEX5OWBr
tEo6Y0IOyzBs2CFL81QQedBvDDhsixzW5Z7T+j9lLiZK9HG/MRdDiiPzm1pAuK9SbC1U5Qjnl3w5
KULE/covZ2xOUYg4DMCHqoD/0ECnMJKvfq3lJn1ulsMC644d/thiIPzuNhYdQXfl0KZ41WXqYaoC
CdGYPHcIj4prau8gGeGJL5192QrZSqsFa/PfD0jw+xf9n/Cf8v+TWb/RR/zPTFMHoGl78HO5cwQR
189F+T/FkpzOV2KimOuDlbsoRNX/lVj2z9cTOG2StlvPiHCsqDTs5EEe+ynEUD5t5g+k98afuV5/
GGxNgy9L7vWHyfJVwpC8nZ9myNRKu41SGmsO37GTb60u+lQiFcY4xj+YDYf/Pd1f8BGIKhOh4vfx
mpRGglOPAFsqFQ6zt31O4ukqL6oq5ZUZc+zy6CYpre9oQeCHrN5Qc5ZZRG1OuCIfxHz4LPpAS7S9
EqM/dIkv0Pe+WaCEiVmUs1wBFVn5Gfu0Lg2u+1y3AsLxvJzCgneBFZ4BE0gdOKW37cl/1NmDU33I
J7PDZzWezUEXX67SljeAl/QhuIYpNpppgLpVGWg9GJpzP10YY0uf1wDGh9ZPzyDnchq0lr0Ehzns
Zx7HYaFqa/scgscBmRu/tuUGowFshV+rZV/78GN1Dkgn03S0yri83vEaHFBJ3OBk2Pf5MeiJQbyM
YUs43vy5yIhg5To6LemoO1pn/hJPCt+h/eLH+1/irINII2AK/Kq3C8XtLiYQNCkBcXKYSqvKbkfP
saGrc8hr0dp13rnWW/E4YPNA9iNuOiFeV3Wa3NgZ+qz4Al02GxVeuCkeG66g7KmKneV199ArdApy
M2aIJs3s6uPq0wLgL+TNQxumeWZZOUDP0e1UOriK5zoFdm4+osS0IZrgyphg3Hh25IzwpICwyNPr
svx+zuPLBVTCq2tBT77tGGnyX4FbEsvr79g7caI2CaFg3OBBxi+I/vl9Wj9cbInee02GUpqn7NbD
lwfuHAwSnXrh+guE26c129efVANwBpv5BV7uM424yKDBbkd6KH5fvz3V11EqtY7gwevy4gFSbrre
nSMyy28kr79uVbFlMMg3TSiw3IDHlGOgRbHiMO3Hi1Tgpb1V+XGN4hIGGHLa34bS/IGIU7rtsysp
cIzEHBT0d/gOdRPymia2XAF50/fNltPB6SKBFAo0wN5WIJ25HwrAeOflmDErBAVpdkBSkBwmOKj0
BiP8tgVYSiq0+/HAhF3An8nwlEn5zmc+QHqsRsllZUoJKibBVOuy7eNeLPmHUb3Pq/TugZk392po
xdFvKYo7ATYnrTAvCEuZvtORQFfcL+wHrXQ8GpwzwMqdea97P9UFPeDhI8lm6wBA0jFMWwFUvb/0
5n51IYVsL4IRm+fbx5I749I7VNKJag7ZiAMAoDIKpC5sOHkcihUEA3J1Ehn49WF2PicNDPKA14Dz
SAcQQywWG297eIDuwSulNVWHF7Njpr/nsgqtNsFQf9JiT1pqMBaD82lY5ljRCi1aBYiWuJJAwUFl
354xwDkikMOtGJqMyTQewIuruPg5RC+P75JbmBvHmNA9ClvPFYh8+GlCLDOUXFf3ICvb1SDVE9Bb
MLonNEYZu86IFCCb1EgwnHOdV8aMzvfngKsSImv40Aq1tDz7HV7xY7XmJnE8kM+MvUdbvSc5Zpw9
khVJegPQV1e3JcEq+fODDchXZrQ0ykYyemsZtxCv9Y/+SG3tMermWZJ9bDa0KHebPyqmbPOFZb5h
SqMQy82UxCLsXHpcXlLxSAtAhzBsa6b2RE4tLxKvEqHmVFnZiENmbD3UgCELZKxB1hCeB9Muc3N8
BEG0H6q7W/EFG7cRfFvBswg8whEBjh8IlE8/Gs5dYavFDNboUjU9zfSrKccDwt4MFO1BNak3Z2ar
Ozu0aqxNtSgsZV4hXY0GaLFel2S60LwG0Ej9USDGgsENQDGNHt/FBma11IL6kY1riCyQJq3thDto
CTiNXaxEqE+PbCiwixMTdk0J/+odn+4Cwd7JSIaNa3QgLB31B5c0qfeJspTDlrdXCtt5H4sd48wL
r9cHbEfZhp8BedjzxDTibxZSV6H6n6fqvmm0s2GGdu3shPtwmVeY7X/r7YCe85qIgsYCkumOC4zE
2HrnsGkLZdQ6rdcmqE5Ln9kNqUoHmegl2fjO8p3jyergulKYFxNz65UJPCB3KbXlFowTiv5AwfzO
+mCJMG6H7yLeeOy7PYwOvtp7ova8uVz/251eZOGpE6hdZZ3mnzSAxmASHyLtCabcruF14uk9eCc4
NFsd+RzBlY02RzeTGsIYww85DCwYOfOesKISCEZgD+HAO/+7GJzghLiqpJtPfyM2ovJ1WtTzJThK
fggrAzdW3LQcwlRZmP2duJoby8Zm+ZKvlveWPhgwof1+tFfO80sUtf613eLnFOYptJHYxTDA4VZR
KZKyqjE/goNnNDXGobdWY5Znzbh/j0eIQF9oSLUW4ZWNUPMXD+jhQ6lCSs3HnhB4r66kcfzgqYS+
i5ryoEaZZoaEpMX9NmDcuQLQJWePpSNfunvUmOexrwcvI3ke900QoawYSluW0tc/f6yVIA/WAGvV
bDx8MJNVIiM3vaNGOXIAQiME6whiTbVAFBjCj3aIzI5et22wMOVxjNMdCsh4pr+jcFEvYSqURPBB
tlKYPXCscYrs2VUXB5nJjuXWQSZN3AbIGfvn0vrrMprQmy5a4xIUjDU2m/onk5RDPRfH2oumuhk2
gwN0WdYBAd3OfUUUjIZkMSx3D796kyiCH94mhBNCQY6dfdoLdSkUG5NegJEq+IxnWamE5c1ts96W
yzJxD4puCLP4h65FhohGCZdMf2bv406VaoJDCKe5UanZVxMA+AGlz0e64Fw9JXVDGianqUOdjvk9
45i/gpE84eW7zTSH064WlxvUJWBJm6ALTMF42qyVdT+L4nFyA044ofrxdLaxkyIe0orvdcJ0Kkl0
jkSR+Ush2llk7yyCf/meilS6PWgCfsuUZSjO8OcL3c/TBxi6GeNmGjRyPFLUL7a7/862XJZB7XSz
IYvByBlo/0gu3msL9gmfFDyiyRC4jLy1wEc5u1h+nZWlyO3z86FwY10Iu5U8bwkT07f+pWjHlSLz
xubGg4lHCDr6jfNZewOy9EM+L7Q5DR5ub5IHpbMSem/9FeYCDMJhM0CnHXzG6SnfUtW7ye5L0Wm+
u4xDlRO04+Sw1RoQWjjNAI1bOlXQk9oByERZd8Aeg1aJJPdr6cYc1BvVwYyJerDyaurVAyiuLopl
+HIhMGkpTVHgGAUYOpe2lsiUffZjZCpXOWoTXSeL+td7wUWCpr2vJrwxN8CSI2FTZeD481mOWBLg
VKcrwCXbWUYuMQEBY5LsTDDZaAx3muMv9yvDkjc2FJCDNHC++LcQy4hqmUhJ02DnZy4WARU2rvcw
AW/EwhPKy0pq/z9hpsURJCSr5tste1mFE/ek0zj1OZws7w2cKS4HhG4iHg+EwnNfYC4gUqeeF//G
mDx3APOpOg+1V0PHLt/LbhBVN4e5jMRTJ6pfIblDDbXmCPV08PpScDHSFF3D/picHABVJQYiwmIO
9/ndBqXvhtzJC15vEsDKljgfetWlON4+EEzA1Kn1yNl3WwMMbfXGIMiWOVvB1HY9hjH4Dc46rnv2
S/Etn+nlDdlyPl+HICdXY/zWU1BtWjZQP2L2q7sNwj89IyfQ0kpoph7oZIZgmSPjTCz969Q2m2sn
e7WNrwUQU6K+S7dldqoZ3XJhFV9p9dDig+ZsuW+21fTipgoSJHZnmOn3Xhd5yXRTl7HGAwCWxr/9
eTdhglDqT0O48aIzOM0L6NHK7eGEO/sKNOfERZDbgKrCsvj6yA+4odXkH/bKF6J8BfczEsoCsyYy
Kjm0XGDdefgmfXGQvdNgrLTYBtlJJdMfvILRz67PQ6r1xwD2yvRdk69qvd89Hbwy3lP6pND2dCmg
mx2g8ueYFAyVapnrBvfqP3pWbVvkL31w3NX4e3xVhNPLCe2F8ZDY62QhsehmOBEsNqPIuh4F+hZP
ECNxL/kIEK/Jf1AMWZ/1+rQRL7+MSkhC4rPibgzwsp9Ox1EJOGOeQpW62isZecpXi99bcMnstzso
K8vXCAuEhCwi2PdHtq47VJqiDRmf9UE5fVqzu70b+L88K4DrRxuVUOFoeDKFRzs9oTgZDPPvGsVT
RoilDZtvmxxqC6wMO/VrDqbgY3wj5gW91bHphmCYE43TDkvZMJO4MyCsB6oX53DNVEc+8V4Z3KIj
Uk0ewaiiChqTRbdVrOejFHQl3DFxQxyfu7wPQNRcpYoh1SVn1cedL1SAfZV1j0BqspX5wtyOvCjW
B2g8P6Txh6SIWAOE+wntTZrm9dRXiUOjOo7ivewrUxv1e/oh69XYLe8X51aKjLKtjF0W+5xvZxMI
kTKEbILSY76WgqZUGPK7xGbmmuRnfXx/zfCMFEqeqeRqW/uHh+/tAGLNvO5hVbJ6H8C5kEXqk4VS
B18Ar//TMvpLDiDmr++E1yBmfx9FB1q+VNGXpSDj9hvhiMWJuI72LJsyXxwQvt4S2RJXsct/fQXx
1opr+ToxHkoUQP2pSDBzfiRAVeyOiwvmtsJ+8Qlvsq5mmmR/cp/hJ6UOJ82uxwZlrAOyyxzQG+uU
LNenF43SjH2XWYZreAToAg3BOw5VS2arOuqpohNq5nXpgxM5pFhvjngE2RGf0MwX0b3EVfGHwik6
coxZVfRnnCx5VnIvzhb+KcdLkOsHbV2v48G/8LuJF3Rz27yqK6nBJmxjXDqCh2Xm6Jl/m9fXBe0l
cJfKsgUXP8Y8zQx3JaD0d7pvofDXYSVK5/5MrIrNxCZJNNThucjRrUtuimjPKZ3Wt6/kvx0kRjsa
yoM4dgPgHJJofiWy0+GBt+mphDAzyQR6Q4ZPfaBkgHWj26MGnvFzN1mvH8hgAGc4hgsT0UFs5qvW
lCm8ZAtTtP7peL9LZCFI51MmccNxxCuGAWqacaHErqFVv2VblBiq93Z9Q96v3Q0ir7qbTISkb+J/
zODOKMIZfCdAbU0oVWrB1vhZDJdww73X6tH0yx7BWJNubF+NF4S28X+/gwq9Sqi47fJdzOKHDyOs
59jijLTjcWz8OXP6ni7WXPRoNt6Zy0gxH1WgR6woGDNlohMKZf3CWFsuLuZVyxheJubvfbQiwORv
At0qCwyho12fDo3TLTSs+V6D5OOK4vPDSR/2vafrZTgsV7I9XX8F54dHXeSXBg0K3t0pjEaD02O2
ptZOYBPVkQyorRinXQKT4DAjZwng2xa4xDS2uZ2oDjo/rPmbwe+W82x7aa1k2Jh7J+m1qP1DZ8m9
l9idcYwq5Icye1cvNR7sT8J5FFg+EwuNcoDMnuOn7mMAlRUU6vNSC7+YZLNyrJj7IKAQCQdPhzSF
ygjLYPj/FXf3TEeF/qqJK8kfcwb+QsZwDzziD7LOBQBeCkeeMRxighQYv8nCuJ8w5M/4vG+lWBvo
aQGucWY++qPUkXkpttVkEKsHfAVjHecJEse66ZOjgJBrgH+WMHFgmN3VcggLTmNnikIKqGvNLVId
ULpr6rFzMhpt4TrhuYgrujBPO0xqPSBdZiEiDID2H6mVljiOEJpzP+pA0LWeytZEZmXQS9LQ4PEh
l+VcGZokOYLhjn1ggRmmnkvn8CPlXY3Vf0ylK0uD8fYjn6h3s1dNQFC9kjvuDq7m4RWwWVLEUinv
mELUNZA53XMIPx+qLCCZnmWr5PQkvIOobAhvMB6uqEdC5KfOYKCzs4OJrFjeuVIJ/tXRuuPz5G8h
OEgLktPb1a28jd1JQY9VBbRo71G9ic8iCUnTEvoVjSrky3fobm58XE7OFArQ7XZeNYaH3nTyq9el
Pwr6Eu+OeAkDRboBvVFgSGLvQFtqa/mpxjit8a+hR9bQsASgD16H7iQDye34eIbjUmSKOAkplf21
amh18CaRSVlQLsCDrJ4SIk9q1nKRnoz9l6bps5mJ8TgqAdF9A8O51a+QGa0tPs3EZpv2UQ7B3h45
HPIrcKA2Hb2HZfQnDuOfeYjKbX7LEdP9OSpGCHEYXKPqvSvTNsfmcgcYQFn5kuQ0f/3+zs69C6w2
l+eN0rLJnDeurBydKri65zoq/Iut14E/qy11QLXNUQtKWaP175gXJwH9iMND/Td9XAEtB8jQsB1o
cIsMVDXuoOcMg+6IGinzEPCgiXwFMdXgUQqS3Q2ZoZJ7Of8fZmelvkkxBEbYTVpcTm8CknijHcuP
530pgXKrI5peplZX4E7R5cIIBD5q65UNkfHN8Qp7onSBARxD3FJj+/R/M0O0XtjH0mEYhR0sS/G3
ZucxgS/qjLBJDzyI/zpZwPEHRVg2Uc+GVaDsApVWF1g3x1/hbv5fX/RzJf8i0Uq3m7HITuZxb4UC
V3Mejwu+UWOBTFGNG6H81QJhDWV1yieKgQLRGMwcjYxQUhtWQfgSMkKM/UQaxpXRtucvMRhD4qxy
52/v1j7Gj5J/FnpBGMzZuXGWTsa9lQ4JJU3g8IC1+g1aWu4PQKQMKgaw6YR93CVxHiLAOl+aB4o+
ZS1l9N0Drq6RhT61OeKZROsObq/EAGEZz+TvQdbjet7ZMVfjGO9qMMmxktuOlcnJ71LQPpCDvULJ
xrcU4hXHixqdx25KEcEVuAJOFE5f9mp+g3hQT79FEfTeXH6YvC0pFjMothPL4jBiRbbSLYQKMv1N
5SwtbRdDFR1eslhoa/2JSkrDf5tOReRJtUIXzR+9mympG7WWDA9Hf/j0/rnjQva8VyBq9zkUKZUY
MOLet2TunjiREZDIJwq0mubaNPMTniB8u7cg2FAi4yq79Op8YkuUDcLwr/2lTXjeEgkRGwegYmGm
G6e73Vvftq6Ah9skSckWLWZuvyB84remYMQqexLyCNjxc6YavNCKmSZkpfO429t7vPUcRwRzYKCg
u163/Mkr2gByaqfkyejIyVlHGBSk9vmf43lW59qMN1ex9MqCtbSRzuBVQ3m+ks7bIWig2Zjj0ylW
mzwUs6mOdAtK4ALc27PlGxU5vYYYqZngapip4MSoJT7e4nts3M6XaiaF+RNPOSdfSOPm/uAgkE1X
Zlk/eiVr00Nz0DANHVzeCyyW+s4szZpiRVegifq4Vd+ec4PUJJ8rCTPckO+H5ZxL4HtGtcUnPYBI
yOsYb9pGMWnv1L5qMO6nX5DXlz94pj+ilzgEebC2LPpXmP2Vl3LdjVMjd1soTmPD8btyU9+UXSz9
X6Z1KcGipocIydStaO+zxXlcluyoFDUdBD1o3J7cxXpkUlWF/z3JLH6zfk5j0/o/deVNch+jXASY
mGUMTS1Fc47eVY6zt2RFOSQ/MU9hP2zA3ZMewCPURfnFhbYgvRu8PuxTKLL3WT578DWUG+d4xUD2
fUe0SwURX70BCLWqcN5jM0xItRa5rLz3N0WKd8Z4KtrHF+q8kalMqG6NLEsRf2kmhNODtSLek3jY
k4t+jFBHa3dq61RupAO9qabqd7xEoUCKIQM9jpaFHcdEuaGneKOCnKfNaNOpssoRBEOH+UElQ288
Bd7dGR0vakahHK2shzNzasi9qNNfm8yorgLOlsS5b8oPMmst5AmVJBHXCGHJG4FhvbiZTi31IJCl
TX7CXKiCD8zENCPiZ4t9RSCnosmQXucRmBacOFhFsxaq4GxousfQCW3Cz/V6NXSQNeALOcsAZUwU
o9Sgu2tqtcjo24O6hfhyg1+Szk10VXKU8MD/hqdJ12vi7T6UwUumiwyfrvk4FSlAhoRwTLSO3lcB
oDoXLzfTQaySalkaFZDvvKm6k0GbbZViHvGVEX3KNw0KNSM992+177VLtqKCJ5R6Wmxj3EkCa8Fg
luj+QNxCyMVh2ZkPYj11hIYWHPZTeu8jasjXmoFLbiWA8rKbyjncL32yljEc5Ar4QIAVubP6LpQO
sgEbjfaAMzkuhB9yVzHopnvrd55s22alGT6n5sq50am2SSox6raZQDH1P3ocVCim3wCAyfP5/izi
weQT7NMhck+tCVIKY1ufKLcCvI3fKkimyqR/gS1ztzt5PnmZJ3396pAVVAHxl+xW2Gzb1kLMPeVi
IB4Q7xym8jum3+Y9WZ1nb1vqsZVCny0XGQybSp8swghtFVjkM3FcSXoxPSeReRwMIQBDyCGxKnMy
TGyRrvO977ZF3ThBITwH2DHhxOG0eONVwaBB/qPMaO9HhRo6oBu/PXaTBoIoeQs16SG8zdcvKYid
18Nu7WNQjHbthVAcELYazoupKt6sg+lS79b5TLRSn9x9j4WNeqxFzFf0PfeVa0tB6q3HpIXNjy8X
M6mPSrfLKE6rZDBgqUW3KqGu+8ufKJTmPzzm8BN68zElBXniU45QB3w63JEARICn2BoL4MM9iiyn
GWgjFHKuguy5WRoGWjwgp9aUW5Q33lnqvWXOtrfZKC9ERcefLsSj0GDem0VkRiUBEM6jP9IGtQvb
/j9HY2Ra/qT7WvQJkIvrZOwn3tc6m+mOZazuv8Dxkl0nYSUTsg7UkDWq5XtE43mZu8pJUDpncpWL
msyxC0+E1l51Cr9W2Abb8VCHVvcDKQdqfo33UbNOvKWmpTgF5cr1en4Qd6OguoG/z+guozQOR98o
MLjXz8q9tUdzhhlTiAMsdWxU6lOInRANsbiU/wyyKiqe0PGDbBxpajYLfPIY8cGVj00I6/Ot3ZU1
RcW6+YUodLQdy4aCebCl6bmdj6gBpxzZ0fqiCHGAvseUdwKeSBtVbpqYPGeA7vSn++Zj1PTuHd51
TN1o9yoZw/4FbH8kAu0aFsabwnBRlJ1zvJ1rBFhqLPi40bLBQ9aAiuVNJW0MctB34BF5/O55fzOR
iCU9qqfKiqbN+A8QozdQ7MlBNDqXHh1wUAkKngY1FgUOmvLXs0umn/7jjtXgJ01mq9Nkmy0k2i5i
MRj1kpEHNBEPw1MyKnmo0RiUGPNH4Y7Asjr6qAyvQ4Sc8ki/7ajbp2Nm64akmuBFr5khy3WrTzql
DdbsSIh9dqsqpDDV3MHsE/2rx59MOPLtrEckD5F+KSDxaZvxrRmtm6q2HgSzhNUA6KdnOOwkPnDx
A85yGDcBcgKHzd5p6LW5mbf473AdWWbw6ITpjnNbcEKpNZ0TeZLaq7q1Y8SPFfX0lcJxGKY0RAUR
OLX+KNIa/1TQDyfDaXPUlbK43VXr6e8j0/TsHnchc4qG5uZ0KQUyv3kt/bNE7XeW2876mDVQcV20
NWeKr7wmNM01YrJ2Rl/PG9wK2+iune33WIKACoEm2i9hpZixB6aNkuSxVRApwR9bxxMwrT1w2Bea
+P0tRZKWIibJZYDkQMdyIwtskdufUtNxUP410sy0+bVigriglgeaBQ2INqL5u6lXZIxDg0zYYgqG
Z6qdkMl4s9HRT7qA1Mi6wOxkcWE+Y5+R5zp2Q8PN8M1wWh0Mvi76br7FaBJlExiel7KDS83FdmzS
OiQEoX9SPKCw/8IlJEfjYfGVqtF3M0De2lmexmTTk161zNiECoVfBqWIezBo1y6n763ZyShgduTS
AuixN8zQoEvui69AQ85ujC5SkYZK7iWF767PhWlbbC+LIaMSyUWV3DDPlf4IcgZs84dKzqoS6jQh
zujFKHbchWlecGv96agozde7cQVytmDhtGkCyhWE0MBmqO56O/tuePr+cXqTBot2b7LKQqd2O8RK
DcXBndExrTexz8Ip0jN44oyubeU2Bi/otzdm1mL+YN19YmYeIWsgFQZTGXQAguRfjC7v1PW6mtBF
s77+L5vAs9JbEWHK9YZ27TJiM3vUgbFzF019xCQSGmXVDFzh3/JpZMlN9PGNpuBJ0Rj/3AqtJJcT
YqcJXzKDQOfn+Sua6vmRepKrIxscJtv4kIyrwn7h9S52DzEbFJVBq4ILN8HpZbioDGiGKBWkovC0
xvj0Dt0We3jv0oWY7B46Um4a112D+Ys+YebouoYbsTE5UzmVN2k5uEM3/o3zWat+eAQYnVsA42c3
5hZvV2+3tz/lPSHutklrAXsSEf3jk0HaymovcHS+7gZDBITmgoRj98Doyo9+zlElm/LtP8/z+xoC
lyflLr/l2UrHST9ecgPsCTWoR3A9Kwv6b1LMyT7Fz9bY8/zfaQO1ynXWw0OXGL/R8LM1DjXZNM3e
hGQJ4oMJkONHWfD7PQ2VD2WtEDyoly/g5KLtrYaVthz3XU5HDZFRERs1DB0rGjFfDMnRSXofYy7O
VC/Sl9BHRr8949nEkyNXy1SngIBxFTrOvhlKLTxMrhdkcCdyEN7c251hQ6Knyw1kTOeuo8FLnXZD
O7LpVy1FdvH3r3wHlxJ11xh9xxWIUXiKXhuTWWg3GISGdwHT9hoB/fPKwspgvmdR0LDFsxljKKSV
dtkN57HjMnc1DY5ctRfp93jOiQziLsoKke0xyCkk91MNxJWmBORo2OGc1WOiQHm2WtvNwsbY2mDF
3ne/UGbQohw7dlBtEa2MNUmBQlvG5WE/e56D1R13PKHbHdUpSdzSSINKjtqazXtIFezt8Uw8YYJr
uCrszTSobNw6HyWNXLZASfCoMzZixGemesK0tDRKpdDCyM+X7B2n0wh254I31r8+PGumZJJK+ZzW
JG7qmcLqtvbEsEK2bFCu5Kg5AXDL/71nT/mgKGOIS3olCRME0arpLBSvszYkjbaTDVtSeIPevmFU
Wte8nUA9QwuB/+YuTDf4uLVkUikTMIMx4iWPtrUMskYaoB4dGOoSLP0gr6LYqPUFy0I2faw/616E
crO4/jIQ6vQAWl8SPMqBPt3VrtVef6bNUOm9fKPfwZP8kN4MRc5b65xP3XA59qv99cajQmgI0Cw4
I+YuNBQ2a+mftvHlIHS9i4jpnUMU8nk9E2yGRGrQKFU+a2QuQFJAS7LWAxjTCbSNXQejX6T8yvUa
9/TickDPuqEg9jECmmhcYTUYZSO+OAcLbEYOLd3srSF9mpSHjqEdnGzqdoR+i+1YlJOWYNgEarsh
xQpuCTiN2FT/7ZUau9U7s/TNpDRyJC6ENdxc9uIecvpq5LeUCxDo5LnNalKB0Ki6X/Ydxrf9x0Jv
pULX3+1L230iXrsTLGVBnYBzQTZKT9QxXsoRn/ETf2PuNa2NlR4yWDCLiyMoba+DIeaEeJ/bNWyL
cK3e6ec0WtWs5Ul5Mog3OxMsl3JCdxN1LRuB/YrlMzlwuchG0Y5l/hK78AVnLEBNBDRc/5ZcE5A2
TAROD1olMB0t3Ssj0vUcHzoRA1ny4O2YrGctqnA58ZKGGXZEI+/1lfQcx0jVjC3r2O3060H3l83x
CV1hdzZFHuNmhfdoSirwP5HLyBkL2aqLmjjEDypoJKnCp0Gz14UtxbYPOsLnLXw85n6q9rKfU2Zc
SEwc5re2h7g9SmFHMKVh4NOnDQJuftiCG1cRAyCvRBwJei3uS5EOAtbIgNDLfy6TUmNnknG0Zddn
Hn1RmqkZ9jNBULzaaFeUs6d6XjUX0kb+KlAjNzOlq8k1uI03PJvYPtgXDlYJPbdkKd91DW/fhvHJ
79iLXqNuV0GhQeb1QJ0RnGojByJidkzD/v7mSZeit80KtTEd8z8lpHqxth1+9X1CwFvXjC2AGX6a
4aYshNGKjdhVIPsRi2NsjTnh+rDOAIykd0ZGYQ+85C5hAVtGz3nF2k4OlEomTiJh8fDifjg/fCHr
cltYMGxn/LJ+jn5O9q1mDiIje4PMm+pJks0WaL9diFfAF2GulOeUt7m5Sv55k3TrrRnkj5+Oj2I0
udxx1IxI/Qss9zrDf4kZYS0vr5Twt5SfjxGCyaAbSGBwpFHwsE8O5v8DGWxF0ipqtjZpbvQkb84p
JmHja92uE3edwIGjC8erYSjdk2WxPeW47vLe3IbOWsEAuTBmXg5mscN9PrlfjrGtZBDpt6G6CTCd
1gl3hXvXRk3FTh8l9eONqENLNhDyx3R77Z52tSTPTmQ8GSs644jVCXnPXbKlIHuPnRrGcx0GeqnG
K6SwK6S68EBicjteRm8zYLrZDPIbK7lXQGgW2LvGIptnG2vqQbePWLdIsZIcIOEUNd7+1cPgT8fN
Ehcllyon+zTQlWJoXcFg1zs/4axefSAJ8gwNSznhkhcd8xQfIp5JdGCZGQ2ykK7rAoRrSbXBkNE4
anaaHOP+wHN8JhWeqyTcZBvCJLDnXpR45DV6FqP49tb1CpuhN1PQoMV52qmagf+7cLnlX5fvMzzG
kSjO4y4MYQtVILHJEB7Z7akP8ya/+RX+KpM2spd2BLo2I7RXEdImUwxLPwl9mECb/JmBj5QEA+/s
2O1Fnjgf8niMw51FD6SyTe4duOGlFLd6NtBiUU6+cLYEmhM1fhmEU08aWmKzWfIueiXaDkdqWwz+
OSx05OFiYxKpNqODUSng3WMhIkDkq+/6IM6nkBNVkkBdH++NB4Cx0LQqTPnncILXDcaVFS0n6nZK
y8mR7Uo7YV4s9j0AB2KAYjlzQp6AWuQwAF1xON5ONKuV0A52LqyWfr7wnRa0S8yhS53reGW7kyTL
rvVHTRopSX0XJkhKuveKVAKG/bmkaVjC4vi52KS6cYBm+DC4pNp0DGSIeVJNDSWSOGt+U9nIayMY
cGWLfCGCwHvdIOzRjMK5DBXWUUVBmNzCdl6cd1p2ObhmzaOXX6UMI2p9/GaYjQloeMFXCkkWgJiL
ipybmIzwC5aObGpxlopU3FPSGup1IEV79sxN8MdK172U8ZFPS+67kd5OTlKipr6FrdE9cqAxz0i8
hVL/E3oUcxSQIEVCX69Ij9YmVkXjFw2sqAscW85ZkTst6RXKuv0nV/ofVawCWqkHx+kuJuPueAzC
QU4qjAkzD7CHXuRNIsfBCRDAYsqMqHefdsdZKIK5r/WYWXaUOU6E4WrQGI71MbUG8lnAISHLMqDs
aCIRUz1Ir6IDs7mSaJDmBIMLL5uPc/cVh1MPCMzhCjQK4u/hhs58y/Yn2d1H12QqvpNYnS31NIXh
h4osEyByC4C3dnZsat1W9qhRwdEJtqqqbeNirUQHf4jPfKGWzfkazb/bbXJSlyzSeAAuPD+KaxTu
OkAF6rE3w9ogh+ju4vMgWM2Zi9BivxEIeHu7SdvosDC4iI9GL/jO3+WzPpr7WTl2ZqUrNoZ5wUqm
DkyGm+Tn/8UzQLQS7e7oypjXrRu0m16oyC2LC0AC3EEujCxRqb2cOtokaLwBlP8OF87B4zIWYvif
Sa6eZMygsYo22bSsUPS3ZwqgYw11f5sJfnTJMkN3XkfbKbdpIYDoyhC0Jb0XMfnR1uucYMGyUNkY
8n1AcuRs3mcPM0vncAkRWIHCwHuEsToPlfXkyG8tUKSKOxiI3ymKG6wJQOjWIIXD4gEn4MEczxxp
2P3Bct5e2crZy6Wl2c7CSCZ5ItmoCZ0MBWkX0SW2ked3O94PyIcEtwKbceXPGsfKhmCI2/xXL+Vh
GbF54PvC9Jzb6H7MH5v9ChTcSuFI3ehO9qn/JsWzGAL7hoRT4EITt3Vbaw8B48Bycw7neThR3QBz
00jRjaJl82xzq7tV13sGwQHelxGdZ3eh5OfvnuVFFDUnwaqoPhUbnVz8SKTVbAfObQT0X6e0VZ01
dfbC8jG8pvarG4bzL2HrGBnsv4waR74yNkbyzSxvKnj9NrCTtmNSN2L5qBn5ffWbJO34EyHXKM8S
8pFdQT0v2OIAcqdhr+s+dpumlVVPH2AGKJcTu1Z6EzYKVpfrouxrQjajYDDoSyLQW4x0XDIqW0bv
Rfxc4zEKXUQlvtAcSJ+pFgi16v4ev7GRWdtPYTVl0mAnet34ip3gVLZhlnkE3WX0nAiYCTvrUb/C
TBFGTR5EFkzp//VgMxAw6Pkr7v5qwkomIAM39k/WWWrur/B+FU54B5tzcIaF40eKdel3bYCsUGRD
WzTkUxuWFztEHhmEPVU31HgqCBshlMbaCpiTKpp980iNzOlHgx5a/TyY5cIAcfw8w5RTNgmyrWXj
x/nX3vEpWn+mCg92V5W/tOgBiVelkzOeViz2uZQPCG0pSnD7NDwF3xOY0jrSSdnGm/qmDOXCojhV
Jz24xvV2kd9Bt6r3bw1sC1NR22q4reef5gH4qoFyk+K079LqyMGrsMqXEcIWGPG2yiCRLDpWvwIg
hpXK1cRBGujApotHHEf/FbpZB+Rs+YXDXO4u+LoTt4pVumDVQJqBIdsdKlE+UQBhZaWt/n0EpfZK
imlzeoZK5FIo6J7C6tdpPLAuGsSVsprcu+MGKHB2jgD3FtK+MFHpMiE8Fk9KE23Vqko5c/WpivA9
p2UB0j3ZDumcNhX6OXa+Y4278B4Fqz+6ydXOH5mIcN1INBA9dZOs4UaZary149hqQq9BX7SjyAM/
WrTQtfAY9pbLZxuWbDV6Jgb4tEbBTKwxT+0HVgbQf+vGPcSKRTE7xoM/sUKcuM1WS6v1ov6tzu55
pzBd8ruUAXFk7ehsd26Ozzfsy8KMyXkFJpbcaMOWQ/ubKUqal9tzfgIcigM46W32DmYgK0p8fRX2
NmgBPx3QVF9w7iR3jAIw3B4i1/SRaZXbAuYyQZkmXVqAh6pkQ9M67YKKuAAoxGmqS+5jF+oKbhaz
OA7OsFzVJCpNK9nAx2xuUwQXWK5MX26Ylk6wqPQW53++EUPN3OO3mWzLPsQbG3/cqK361fLds8PQ
PgRlgZqg1cKSOyR9poOe5CpAjAZynzzvjgfU5SZf7aBgX/9a3+gT0t+4gTMpQ4uWfwcxUAjkISRV
HBOtihwwYVDAjyBfg7UM+h9V+lPRXtimKqHyk0Ex+vJQMiBn7gQjFHw2gnvOLV0VQx7MtA5SXbt8
E4uX0JwkNdgTN5jd7CzGxtwZmcgv12XHRcnTVHXN4tN7qG7wBWaZM2bl+e1CXkmlX2xf3TjkrZ4b
H5WDqZw0ZzVNI99GWJBxDBMy9jrwsMTsWQYRAsrO3D569QCS4ubnRID84plaX08/j0MAQ9NMhK8L
rZwDElZBFQR5P/KTqzES2QUA6Z2lAjfhE7cuLG18DwFqHCzUIA9ym9lhW3jKtgQAsJ7YfgxG7rVK
/QytjXrrpuW5Cs1ZOfwNAJ3e6NUslzzVoYaqc5MS9Ac7unyJUqQ6EHwFJMfo/6ZTc+5Kep8jao6o
56XlNss91ptyAghERNYTwdJZY2p/sGuWGuYnUbHRbRObZvCI0zUo+t2HDXl4G6yY2diXPP0ZSzn0
wvo4vqE001d9uy0yWas11YCPjJY1/d27ZaL9RzbUIHQ3BWfh+LqzxBczBBFh6AmQLYtu91z21TJb
zWDvU5ZSAvpdCXFjh/8+airuYOlZxCuWnJL33PYf4XDwnPD7ovy0mLal9twnaELlTN/kQCkm4ZwM
Rlx7mgrzKU3oQT8zcNScwRuaeIY9ufIDoqVQCzLSI+8c1uCzExQ+OCGmfGiTBB054PANxsayzE8p
/re/oaZZcWeBGpBxSBgbO8B+leuz6MPYHDVY4Jza5D/xsSyiUPN1aT3r4mjhi1oEwRs/KnFVRdFD
pk++GztM+taH/Ca3nzn1eFzCzTTjUOJ+zN96JBMa5iXfMZdjT1iIbIg1O6/8dVAX/HiSs1LAP6YU
jjk6XAaNpWJDl2l4sjjbwzcREar65+iDdSx0Hu+bdCIZXdtZHAhJQCAY7I+BfkInHhh+FpOm4/kL
Dk1j863jlS4MRZV8vPYH3HWZW63yHg3v9PpbEVXs5H6lZcUYNYOt7KeP0/SlWDe+H4IinKbQJ+4y
te94kUGP6SKYf2dXHZ49FIUax+cirRHcIrO98E1XPzkCbwksFOOD11d6ljYooqFc2PBzxmsZiB9n
GhMeEFBKSq/lJvmjJrDxVDtA51CLNZFfvxtHYz33VvGsRz2AOPJxQApx8RVkLRnERwkSxbElrn/3
8WwKSUiVV0Nz/xBmOsI/JjQoQwH8nz6aG2lqAYDVntMv2/M4eLIuR2ubqMCuVCmFcY9rFyBXzPKM
vlMRBzX87/USnwcrrxphB+0YfcBTXGJ6G0vHsHYlRdPJeaRCSID+i9cNkzcFUhLXh591HtkgzJ8I
cF7xBBIZgUO/EbVGLvWQkKdiB01uUZnwR0QJN29bGhg78LxYWkW48pzLEI08ySSWUZYj5CiGOgWr
YTYVS8pd+4NqZtOgkmXmcspG9XeT5kmAShek+oQLPtxIKIWEu8PaI+JlcK60HgoSX/I4zOF2A86m
vJI9p49wyPDr1sP/g/QftrA2qY967fREjD5JHBXZpJzZ8xvOZWF9wlbnGnyy8+pZ/bNdHW9H/B0B
oIvGx14VB5l20gAroNLEU/KY7zgkpWRzq/mJa+xowzGGuJg4VpiUU3vgfWlIIOUD/RxbhXJT1Kqk
ZO74oO0uUmiLGSFP1ASTPEIu8/xE5kgsY/NSQQCtgU+YFZPEtmYfC+I1bQo4Jr2QOdidPyH6OiyS
dt0Bj3watMQBg58h8ubow33K4N3RZK/EKcgU1BWC+B6Lu7XmcUX1yKX8MsUeGOxkuSu5tcf8DaRr
Etwi9P7bY2X7zswNLH7Xd84EKEpHs7iZ+13HJWG4i4DF5Bxo06J+oVOLWXHyhA2cyGBNc3X+jOek
QXYi9ocWiJsEkc0Iz9ubb0bQFSQOZxQa5+v3RMJdwEgJJVQl55abLSVilY8iYBNW/0JEKqmKlYJb
Wdq13NUPcdf8V9QhE/RS9Wy1jNT+Fd357Zoq0Hn7EaaBbOfhfSOVU0s0FGSXCziv9ZnAN0Ei4SI4
W2c52wLjtIuOca8wpxN32aptRvDDZJtWCInfCu48xSvgrb5/fsdWN86WGDdyT4q7hJKFWpluf8Ap
pEYGsBRuU+vYlVUzemsYd1TfO5DjLk6frvArqxmb3J9G457Vvb4Zyb/UHZLhv/RQ4RkDj+I6LP3q
hnyrJdfOAcWd9p6NBM5J+2cP45SROjN31Dj0LFLa/dfHIqJclhKbKvwJ5xGqqB5CRuqbwVqnVnBL
T3vIktdN+fuQa5dqrW016Fe0vdfDtCk6PXdWBgSxOw9JeH2YlK1he8axru9wWlGkGZ/X/EK6dvOe
Wgc5WmyrR7l6u2QEICUzAZffoM62k45tWEuOiZpkg14yYzl2hdvzYoTA9kBOZyfGziBTukX0NHuH
cdpKxWsi9laRJOBQaX3VppHJba9DQBA6zZ1qgUJKxCYhGkih4CvLgi3cfLD4YxlGYbvlWFNAUF83
+8DVG1gj6/g1ldoc0w5oVw/rZXlMFUWTgLydzOBVWc03wq9QBUWHC3eLJuKnsab93BG/TO1uBPiq
752lJ85o3TFfdJVXRzwIaPBo5voeRGrIhEs2Oqx99C5HbtGUkcWD68WUCeeunj7yA62WJceKdldw
6xssZbREWuV9PbuCjo3DbQqqvX9kLmkDgCR+0rpVChhwgBcAT8Ya36si/oa/K//hjdfU8WF5kE3P
ZUWVEU3qV6jK61c78NzpUHHbpPKkm4NWWGPxrURJ3m+8V8oKaCwRidUYHr7bnMtoleqO4kDpgy8Y
WBaj6aA7a1BNK+xw8dJ6ah197KEo5hHvgth476hKccbweV+H+96+IH2UveRU9SZ+JY7wgisc0vGH
tUkFwJsWC1nnpUQfYwMvW3IprZOAs0BGIiYgrB0n20XlM4aMvvp53MmTKnXt2NtkJ1ZjnCwtv5b/
b7MQIH4hYgjJE/NxEbmYhq8u0Hsm8T/XZfXmIuHf+hRUf++LDgq9Oaux+RWTmN+7N5wOWJ+JL/BO
SyfxBGmdv49GUQE+wVbHUeMkPt3cWfPlXEjTN5t0NH+s3PFVSdKq0alxXzq2uV/uSANwZUaY3qZK
XHaefRYWGwejWJqEc5oeoTEY6JBi51RkwBlpekJORlqwi3VX5Tnl6yvJNapB8hIio6llkg5oujqv
oxTGMa0EAvCXJFSKuSAFVg5JjkGc5tOXdvy/yOjPZOKNdeKlQuamcw8B3P8BQlchRmpCwRl6J0q3
0pmG9G15YIMQH6h8UEasGbdVg3C6ZhL4kCStyqT2Zeq4CE43xlsguGQ0HocIMZchZ1kdZMefLUkW
2Pdo5jWq4KhDVgMQrx7PEn529ouHKHhf8ZLqq5fj2jgnvck3Uxru4kA+Fqr3xNxw9gTkRtT2ozlx
pY76Jc3H1aFhBOp89PNQ78452YLoZZ0GZC3K/sSKEEmfCZbcH0qX2hrpNfNnPfIaWby1wHUmC6dM
Ull9jA/FTYQLB71KDppf1DXupe3u7gYOQnngNk9oLV4U8RRY7lDVY4s63HW4zx6W/QAk7ULELMkd
A9ORfLSpDS/k9kyvXFwFTfca0mbC/0ANfiOAqrQKuzFny7zXmSvN8T4eJEvidCf3oruLTopnilsH
30L+OBzKbxwY90qyWQDyddnZqqfbdwa9FdC9EOminZKS2mFkdEx5uIoGTalduF74q1b9M1LGevpn
8HEByRcfrYThv7PkY0mz7F8jvoGNZfWJ2qrr0gXM2bcoixHAnZdmpQ9HxuB5m351GwoboubK+Bmg
w4/BnnJiuP/Ml1YTNOGm0g8tpGmz1hQUq2oYMfaSfvvZf+rQUphG/vhRRaVUMkDpB+P3Kafct4r8
u5get2ydUYkJ48hc8Y0UHtJTWl/4+2jgLSn5lE91m+7PVu4uS/6c8T18nALaaxNHFtzMw1GLU2oo
OJdq9muKvZeXX+wKOf4D+soSiPLuaLNOyBZjb4mg8qSXO1xClvBcrjlhfjhIZCJubf7MeBf7vc7r
HdRwPypfIVGd/C8cFiNdfHE2VEo9i20HC5vJpD6FbE56j6IMPUEKxCseO/qoNvC3v2fzGDs9f26D
QiFjoOsdMtll5zDty1BBDOy7rodFLxDU2aHSKEAvT0cxTC5kxX2mwnPYVQIzGCGS2KROzpVh8dG2
TrzUP1CD79FMCExmiHr7Z+SNFrgajRA/B0Ym64Tb6W8lqUOD/V6UeHiMbbhaxTRJXaW5h2eElrVv
79lU97SSjFMi1bPvYAxs5L340Tw3DgzKc688QFQ7bI7NwBeuTC6YX7Pz2xStuSoGDSYfwCsHh6PR
N868pCYOkxSTw4ZadnGfEy3JsG6256x+vCjBthFXpLh14WXmfoOuggj8gs+uLxWm2ryrl6vjmOeX
aHhBE+Sn2JQxtHgP14ZGcYytiXi7T6JtgqwuqM0aHhj1KAiDXH8gxPB4py2Ez4Vd38R1t6DM/z7u
g8c6sgrePyvco9apxjUAbrm8syv2BhYHQnbCzgIAgjwqfDELreYmMw6ah+sdoWN59Ju5IJmOZp/8
2zOfcIlH6ZJfJnmKM6Q5wWiSjfJu7An7T/V+Q9+Yw7bNbwia5EHkO3lxIrhd1jg53YZpBmRyi8M0
OnrPvuMAhXOp7clnusLlUl2mRcld+ktgqperyb1QBTVTlTq23XQ80bMnj6O8ZKKaIZ1dVDJWeloR
KV0bEhpahx3BSIB2Pt7AjHF4lPwr3xTVcucZHWSQtGE7piBD1ccgBczSeG8Zb1iKpF+Q4ACfbrqL
dmDsn/a5LoFATBUWKsFyS7+l2psSnIdIlUCogQMncR3ZMEMWjI/w/5MAnZg/GA50jLmh9f1JOYgB
st1+GxQ0rYAQa5y79yGmp5anM+RRiHodIsJ0Y16F9ogDy5O3y47x3ZytMMWwAAH/7ymjtRfcm4Be
lWvQjSb55BpAdgnje2fHmshlKQeQaVw/wB/5xchA64E5vbe413aXMgh2Yhdk2qEGtq50UkrqEgbQ
/wQ3JON9cTN9wsve8zkNPa86+Z2iPYo0z6b88cJRcvsBdHVciFjYOcvQtS74ME9j9y69mXLW3yjN
Xp5ZUs5rCFq8j0O5oe01td6vWjk/RmnWzjJvh7a/fgvuzRUOJUhmTSadsfd/ZiLpTtEQ3Gmkmfkc
DJWwMPK68Op2wmMvEk7+DZhMr851QJ12KJ3f7q8Y4YH72YycZpRNLRwFUach02zqAtEN5KA3KkR6
2/g61ErVr7vdQeLHPkXz4ntJePjmBVyYGHbDWyu6LOgCVkPhyP7VeuBD2W14aL6h8Mgtq8TdKCXq
zZY6TA01oBela04ty8MQD+VPfdQpYdyGYde41hjGYDnT+aqi3ZtskrF74lA7feRjptboRWF9Vlyr
wEv19+MuXTP2lJ2ctX+PtjoGvzGgdm/Hct/HEPVvmrB3s45Rpu1wcopuNTBj6zM/XdSPR2qB3Qkd
Jp9C/DzcQ1iNJCbmgq66GjaQc//YS+j6PwQXi4DXZahxjobEjy0qaavxY+8ssVLkDlW1SI+ddufN
AXk7xK33Uks+dpAJDR2+Rn/spPXcLjdN55Es2riL5Sk51Kht7JRqTQV6+J9Zh0mOK9DO/z+u+4BH
FS7O+mOziybDJKXvKZYnfkLagsY/kC8qRVy2vUyqc/uPzQ7kKSX9yGnzNa7/bUdbGls4nSkvFD5i
M4H1RzLuYoL6brG2n7QIihb0Y8ZAMtACQ+n/y419AzugG+Rq4/pLp3ls+WH5yrxEGLVZPaxCC0m4
dXsJ1bvV/i81pT4dVXqPldnN2zHQHcfqzb6xKvWFhVH+WPWKJRp0SgvXgeKSsgxVviDAtan3n6Sz
nXYWTHlafajxgkb7aV9+RFyh8I9BdFnsZ4YOlcQFWT6Nx1Z9H9t457z/pXVDd+spO/UoaE9mMVcS
z6FQr+BnikgeIdgm5+dAWK7tHGzVAUtfMTHBiASQn0UNHu+eGFYApZVlfUYY/H4V564i9twwB22Z
qVjBU2mrz11PGk0mD8YK8sGIwTwloSZF1GSLRUVGlwxdAYtV1hIK5g6T5DCJX0YgRxwf7CENlw+P
IqtV8fC8nmLz0aAFb5AMTS63zQGkSPGHOlPYIgn0R/Q7m2M+43euz+IovdL8KuxG3xDSnAnSrKjx
Ab5ZMe2fVxzpTTCbHXMhe+ORz9qa80NG0dMGTPMfLVnN9S7sBxqsbjRkpR22oODHrj2oPJrdPCe3
A7ElN97rrp1x8fIe497luDJrUpTbt2SL6fq/bvkznC1Znc+IaZ7ao57nFUEun2NS7SQpVqI0rxiv
6/us16q1xFHsFEUMrWO4aMJbS/fkOFKovF9UcZE9cCjluXqQJ6FsxLhznb8TmkHKbjY3hNJ93JC2
ZqY6eJgMcrUnDPtB36yyWquBWEijGu/2cDixGajQG7YWwCeHAcJ4lhJDRf/G0bDKWAs/rXnqWxrb
vgo7jkgeAXPu6NM2j8u4aU5r0ixusBq0elLkkK+BdWVT6aveKrIOPrjn9fdKFxxFEpdB36aD6OIM
JoTIN1cFLoNnt97+VjaNoRCzAnXacyXtXbBB2XxrzsxKIiXPs96RBi+e+yTdmH7KCPbfQAAcraS7
H6Ltajbrou2up+SffyjdbPqkgfgq+TKhv8/FJqjJJKdZY+RlC58q6gfVRydj+0SN1L+CxWOxKcaN
/bLGSxSZjqaYWDdr+FyJHeWPYu2pITFg19bfciVaA8Bg4uUW40ea9BkGFnPhcnZnjqer3TVQHmC3
hDuwlOCnzaqCHhkcRH6WyHNufsdLEPQNereUIGUkvEc5Y1mWqWzw06z6QI3a1S1jPTRrA875p4dH
WW9KzQVl/lMB2TmvR/w/8tiECKw5MisWrUPD/DQmvi0R+A3ZhpoBIGxMKXYwcgLaVW3yBA5MbADR
awJLnFdy9n8lMlhw3lhDgEGE5JFi5Tfo84i9Zw1hyMMuqwyX0N2So/XMDERYIlwJhlI2G2OiJuMc
nUMjRMk3b1pA89hSWSd38SlHVYw2kXYz+9fX1xXXH3TuOk6U5s4yM5YkYZ4JvHCo1T0smIPgQV8g
v6nNyARaDLxumJ4Azc9k/AoPvu01MK1BNchXKGrZRjXDNiA+NBF44ZeZBuj6DQTNOkILAlBA3oeh
TzeAmCjrDaHSLus6AF2gFbXJJH5qLAFVnO83Nnbe2lgrrznFdEL4jykmd3eanfaPMB6d4YPljrw0
zVN8y4WhJcYACHendZv5k/Ybg7ctX8HZJarhlBKEDJHJB4Age39UJ9w0MagamjK5lw9PFZFoHHEB
w5cpijIznpLzOmrER+rwrqqsMi8L/ngR40Z5m+otishGvelQAhXuRFXx29RBTdai5PAUdD5xeFuR
7PYq9Qtui2X/bs0YBs1VvIwnwsLDbmcfDMjN82ycXdxZG3TTgQC2iBqtNRosNk1MD6lIF6PhrR6I
nB3x4U/1D2DA6a0hHaCov1HLlx7vP8LRTSgynWjtxIc1dvucs2jfVeInpETkMVKuYDFaGuMce01H
/5TENvVHNdvYrhecE5aICd6ZwLoffBgMqvg5OXyVxhOORL1rmgL6RZQqryApSaaQsE/7I7YX0naM
4yGIuXbTzVRALx2p9Wulmva5W8UJCR5yUbE0pUC/LPXNzVMCYQGvtlRT0xJVfqh3snfACIKAQQHy
h98zTNwVeYiyywCtieRvsbYESsk6r2vri1Achi8tzoaAe0JALzp/nnr5TAS1YUGN8gYqFHSZ29ZD
b3GovuO1bgph3SFl/bJvtHdSWroACl64aA0zkdV3UfqmkbPgPaZby9CaxRKl+yKJRLOzpDaErDrX
5DV8cBv0pVdRcmPYH+yy2dUIWImMccIs5qn/GByBAXMlzO7gAAtZqoHNxY6VifuuRPh66u6WQf+p
adphOG6wXtyWz+RtE/ls1oEWfyIHBnvSL3yyo7i99Xo0xtKWB2wrs7piTnzYehkmjiKP+34Nk5QB
EzU0TSfSuSOymnMcBb40LPfRa/p4yF1lDgQgBbSDrD8SstEbv9IXeUwbqAfcjPygzr+D4XpjSFOT
MyB3yB1jN/VyosUgIXYn4vaCKjGMuikQJxC10tXp9PUMt+okomxhI3dRTyhO99cNRytmtZcLTiCw
nQw/W8Wv8WcQTVyESBv+Awu85YsEfusRt+3PXYJM7zqep0SwbpUJyMAqHbut5ekZNXTf7a1Cyc6i
hdD8ynlNLce63+uBYT1/46NBoGu2vxKYGTnCi1e6vSE845mvm2BabBNWRfIdghLaBuMz2l+4yhAl
lVSblwT4i80pS3W+0X7B5RWME7vk/fOnFu9MUnfdguFjBoKn83mvcx9UncetYup3fXm+85Xq/0JP
zEo0r7mwZL1WZ5lgSL88GUzPWi94TYl1SZOJBJa88j9UT3OLHaNv2G8QJrRA8u6K8QOsy7P5x/kr
8/QpJW384FUYvwYvIGpwppt3lYq6cmdmiTuHvmQsGbKUvmBVm1TUkRSz5WzFXcoxeByhSlmBTyO6
ntZLJ9RB4SA7dntMYrBePvGFQYFU/Q7U6OsIb7wEJEn9fA3/Ko5wgKUnQi/peIrSYgOcIm6QeLVv
R0wVsHL0gYiyi8aQnl5127ceYTQleuH0g7RYcr5jrbiOvi/m0B78OrW1Dzy/wDr4Tyupl/9vju2i
J1A7gFAa/seiUlS3jpffW4JBK4szCaOGFrzxlrNRjPwt5SBXZEVsuHv80ubN0wRaZbeL7waK8uDk
vM9m8gJEJhVdCYAGC6HDcLdBPXgCEnztAlpgd4NQb0j+XPZzHFfclC95hmJLSlVJityrAFVNmRtZ
WnBSv8aT+ogrrWJH6C0efJRIRFB+13uUibmBfALZepSAJHMxlEsC/xq68SyZOiQE/RABHZbeeExC
qbgTC/ESQZNlOfTxLQ9fxey3abK5JiwaYpYYi+ZYAuWaQX9Ern3Emc8xWTd3xx5krvxPdBZ5C4ni
KbOkEn5dWoJM3jIVVC78buCJDmpC4OyLEzTA4PEn/qwZAyOCXXj+wqUl9KBVz5YZcNI8dG+E8x7y
baJU6mxRfWBntDNRDs1xcXHNJaA7vu5O2ih+0nHOHdAk4J9VVXZ5Xpcd2L6ahmG/gMPjFe1y/lAo
t3JVoNHVSxpbNxchgwsq+8APjvGaECqPheuHVK1vlYJfzyUHdyQHb2o6CtpQ9C+25zU5z2p6LmNp
hMpDKkWcbDWfLTkm84XA1qzKqAFyhgBTkvfHkbTgQRuRziasAXrTJesa1/aVcF5Hf/614FJTCOKc
wR9SR/m+9IlJzDW6M77INXiwL4QzLODVl70ft5WiJFNgE9tgUKESP6ckso0o/iiJRCjqSsbCm9vC
HsEfExjv9lsHIVIygqW+nS6RePpYHET0ed8d3OBHowUPj1Oc2GiOLepqeNvK7fLx4dXPuIAp8Acd
f5FfisF79zrxRMBQfGgwfeOK1Gxt+LiL6z1ZC4u1pB70Gk+2brAtDhtZFMky2OJMKy5JKT1JNkqu
9OYMOrqnrT1MrerC9FcIO2/4jl+Uy8qB0UcDa58IrCEX8yCf4HpAakCe62/Pb64DCZXs4ps+EevA
znv5Vh3IkpSPFcp/xgdL6i6RQaaq/NVAwyLls2IrVyQamx3c7xZgMxWdUDbi4yvtBVevqo8fzNIf
qhDfTwkaGNh0RQ3XjTwBHN+lygRWSYDDMWCM2mPoQ+UOYeqcY2mHN6JkwRsvFPhgt+d8TNgoLk6T
PwvsDM8A1lIH0Gm3yvgRBkYrKNtsqjT6L29kIedS9UBPNAlR5TTbrFQ3b3FfumtkJ9Ep+ZZMkaOe
An2arLC/v14JCsJtDeTJV4Umzby/w0/sx/ao8XcfJK7ODUuYNXxNyIe4/rJyTrBAbnXVq76tMbae
f44TLsXJWZYsSX4w6aDYyPSAJI8/qoDADXb1po0r9u4iC2ZQi8q6LGGS5t+KkU3ToKsWunvjr6aj
WgFUPRFpS5VsQcmUo/UQ3fFvGIsRD4/EQfMCHdrX8j+vk5j++11Ws7X7iMLsXkjLbbofVIPJPkjE
s1ZWtUwWvdhfWombBL01+fsW4pZl1yFICuI7GDNDJGftPbM8BB9IDKd4W3zavMeXX5ldE5tUA/vy
9OSjh2uEbH7nZTDmy86rphYsqAadMRnAtcRRMF7OaQ5tHh/d1kkUWHEyHzSo5KA3Yl6zFn6WTY48
z4TiP7+3fLeHrep8M8ewuN4HfdqNpP5xtQfMnmPYrlGOsE/BJ6a+1Xyz2Qv42pjHICSHLk6WL+FY
U9pdc3iGdtd3Aec6mBPeJHrnWd9ZTt7qGlfzoJeJJdpRwEVhbi/8Ci5BYqNsJPb+RLZKhCTEf4dP
a1B8UT3p9npfkXnKykaQz30Zf+4xyWnH+w4GyCjdidjxREtz7AuEzib/eoEE6MrHWrRlXb+v9Auy
+vk4Q/Lyw6s4tmnJ10e9hrSCObneCak9xMMNuRnWwNbRou1l8ijarHFMAmHe4iNyCpYVwkzAUh4Z
inJt90r4jeb3U9/qnfGXkHZ4Q3m2vd7ekF6rn3tlrmX3pXuXi7oTfH8j4pv8PCBlBZeCsf6Vfl1v
n6lUFAwB4es0nmGmR9byzeoL2Chvi8Hj+WhlZXVBf+o2ncBTPODin7PIx3trHfQYKQV7v7EIM+Ym
oZu/RmlbMnreZKIjDCaC1UsKitQLAypJahu7h1dNx0De74Zj4zZRLbD2zTu2PU1/hFskdgLF/Ga0
hbaUnHTsKAXeRJkMu0VQjxhBxC7AWLBYfrXYvy9Zm3kLdhM8af1GNbbzU5KNJqHePpIe570VaouB
UMD/JW+RvL602e/Et2aZFBA3BSfCDkYrlxGuedXn/yalRNpC2fWrDljhy4fnFtRlIGf1EXPRCjdR
zKVGfFknue7M+vPo6p5xzDtjq50Ma1zWsN/jMMaW3xpL9fsWNa4YlIuUGcwE8YM5dXrQ+2jkeoyt
WK+i85v8kYjZT7nhrjUP/+4vTSbc24k7eBC4wEcR0lyO/NGr0vf0ZbKn0LzcpQzpYWhgo3xruU65
gA5kdsxo0ClhrX88xzhr1QwzqBaak7iZHBXCzDAVhq3ZiABuRJXZvQXmkb4gx90oECbLnXwjYqP2
pV32n5Zcbg+B+K2a6zlTm5lf5V3iX1+mqtxUR+E0dsuQvMHt3TNKTPdwty0aCgwJY077JwjMjH+i
XTOsqTkybygNUcdbsvqyjjXD1dvOl3AsZOyJu4oABKaJFTZGmfqm+zI6KJFgpI+o9jtkCWdrKhy1
7aMCDcUe2oQ1favI7iNeGCmEckaDnClK+jeKgGoN0/K4JhS0ktPXrlUuce03obH8cYpN7WJd9FDt
T8U9X6FNLcjoodC84+fXUiXzpu5OA53PoY4BbOenhfc2v+g+lE88DIuypFh1NYP5gKS7X1qwEkgI
zrqIAVPw6oX5jwOpSTiyB4NzAsd8i16sIh2MSEJXPM498acnzyJDpq9s8jr5wi89CzOayJLOk7y9
Xf9Arhnr+/GEwr+L9A8zhsvvxtdpYb+6mAh+tHUSaw8WMHg39Qo+zyzTd7OBDQOCKevSyg5NpSys
cb8h6b0LwggD4E/tjT6zzfWgnq1+Js/VFVY7TKyKVml0OGDkBeULoMaJ4fi06/NteJKoPtrZTjwc
LGWnbKmFuRd3N+JeMv4Ilx34lcaBp+g9h6ejrWAsyVmpDacbXym8a5VUuaN6WuLDiKVlJBpF2j0R
OjtAwROdwB/kPMVL75JvxoPfJ+CSuOFR21nEBWMMeVIVsAgME+ueDdQOtEz0qJRGsaaBB5AJ4f07
xH00vOjMcE44lJ9FXSVAC1VWwpDMiDDO2nvzq1vKeEY2IKsl6MNHeH9PMeHH06Gq5TP8hQ5yrul3
XMoer5DRWAX9+saUfxCAs2ET7jXC2ay7zUhEfD3PZk2L+stDR8q5xoeCZ2W2hBlhqaKUGNjm1P3N
sdI1tJ7DkW12ZYwbOwqchnt4Xb9fHQ7fIvjaOY3nheBycFdLiAXMa9lyv10cRmHTrMz0nvpGB+9E
TchiO/GT2sawbQx0xPwb60pA4Fgu1fwRgbI4v5Ep/+hyKo+7g8NBgLv/s1YCFLfExqscG3vokMuu
lm4XNBE/oOzQyypuYqncxj0w3WP1vvF+MI05ttsVnkzQBS+M4RYqWGA+JYHIfRZmqx2lKHNMQt12
dl/qWweq3mdHMYFSYV3HkqTi06kkJJeNIietSw5RGXDi0v6Z+pe/1Gl52LytEKvuUrnmjInDA2sY
gCZeBV5YzevMkQZcRuEBFYfvO9oYQhYsIzAJx9jjzvluND9eALKyQe/TfwNsNEy8vn2OLZVsjKYP
/HV7P3fIkSJ9ytHx/4XNrlllrVD1kQvV48HQ8/C8u2VYX21asqo1P6Ge8vhK0AFGsQ0Okxkk6gaf
STvmjP/fm+RIYAKWVCkPVqBu/HMyXpGhxszSRrjDepoZH+k88iNSXT0RxjPz842LzMLOnadp9zTi
ssIerh5WuodxacrFpaAMnnqG6QkJOq5Or41PDRGrxm8uWgV4v4AVvAB84oRaS559FZtpr3umvQP0
SQno5tlGnEujAaxHaYUR5zDpVpICxXQszBT3Cl5grhjiusHhmPciPCnMGrKFZgUZW2770RXovFCb
iELE+POgxQqmHdnd9jTk4yviyxPwOZBfUq9wCYQTB+KFidvWEsei2mmvyRbLP33LnIpwLONtQx2R
jxnsmbf4YsY0u7yg6jznaKJF9wWncvsm6nQH1b/e+H2vei4+bWBldHGyB4M3LxHfoP+65TFeeJI0
ATZ4ZrKApJYtOEzIaCEfS2lnQxK1/iVRJYatcX9oK241pg0bUI3SXwTZapCqwPBE6E9YefsiGidB
/77RnQ6/DUATNp6tKFpiFezSOmWnuzK2POm6i1puly6esKVrpmygQsJaTJXbjRer2/UfmRPPTKyd
5UHK4FhR9fZl4X61jsdjQUOXQ3JwXqO8OP3A8vDl6KaS6fukGrrVAYpgW3u3oOthIwP4mip5IPzl
nOJ5Tklc2ZAXjdgGJ5ACzWi0fB1K7E5As/cEFdUHs+4fh7dDFMKaRLAycOlqfAyIGRyxjH4NxkRW
nA2FTKO4WRO1D9huF3UPkW7MBZf3gwCoJhITxTEYExJYJ9xZRNIdGTr7Is0xuRdKnE0tMAoArqfL
5pcRtpcxbz9ZKYQm04KKJVTV++fdqwFuT59s05UpMtZEgLfWWvwMjx08OyU8/3NYZpOcAAbLldfD
Nv8ccsgN5PNmXWMpWN/GrFygDKF3GzPMq2F3b+8c1+Q07bgWB2hCjPd+QJgo+nbEBnPGndB2KRa6
V+LNiKjbzXhQOwrC4UxOapaPBSLjIhD3urtArT/uqAp+nzXXWFP+l6ZmEiOQQSjGB7b4DiJbw/eJ
XdVncmpbfv72UB/z4FuIYRi2anKmZszvlpGUeTrhdGG9NNsht430FZ8d0G3uZuwS57aWxpesKzx6
hDIn7CEhjm7H9YrFv2Su93sn18+iZPixDrnaX2zcUsBl4GZnkycLkTR/6O1f4spOvXS4EW2N8WKT
b5XcTxe2fOi2Tfbwj0zKH+uGP7Vjd6C9AcWHYch1s3kxyP5VVr3yiOA2DqKk1zsxW1IqbyNnmjAs
nj+ve8fbyLfp41w9GK/sAhfqlhL6ELImItOPAKWsFyda331MssC6ROxW0iebquvTem3hWtLPSF06
YfUkV09jWE5Q75hb0rge8vgBMmLPrvqJNRLR+FhHSAOxXEH+KJ+u7DM/6dzXsoPCv7pivPmQWDYI
UNxNmlPc1rstZt5bF5aN0rk/JJSBPPzxxyCMZldDpOSsFraPrnwW6v2Hxi7Jtmj9Mv4jj0XBeJ/p
7x6P6InJwcDbj6xB0voT9xAIyknTLK04mjjkXMzX8ENAyVDePvraWhACMHppLKxSwvN8tiV8VYL6
MQ0ZOpQy4yBm1tqmbHneCYZf02qRBsJ2I0LyKZdKP2a5O5jdj0oqFILTx5goyK3szZB3wje4cSK9
mesOefP6M7Nok3k3zUlLGcUfkUJqW6xSQClqbIgYiF6YdeoVDZe1fgUJgE+5N1nBpaBH9aNLzwPL
AORZHBmSLTlVSX1FXDm5mE08phaNp0kgYo9lw068Lo2r4Uj19JOWMM/9ReZoSL7Bp0BwEN6vmXfY
OkI0s6dFPh5JFi8rmKUG20vdLNcV88zzR8anstIafNjvHgXGkMosLcCWCRP9POd+0zXB2czp6nUY
vCBgxek03/0SkVAuSMIvpn4wl7LN3x0sOWOWtVjiovmbpbodSJ76wRwzWC4XQhlL/vjAn33PGgKJ
2Z4LxJaZ0yM2na8au4AY1iBwU9+5krck/dtzd56jnnp1KufV6qXpFECIBAiwMfSlSIvmcrPIYAoi
yOGgXput97l0wEbw5G4c0UoNPf5c8K3r4UtebFpaZbHc24Cxy60oBPwdwq61aoOWxBNj1uXB/elM
GDS2/NLiymHemnKM1ir7g1RaRlQqasxfZHLm1EFKplF31K/MscEnhHk/XJFA/+arQx/7oSwGjque
4D/+FhtkbgfXXCXU0hYAJcgoRACjjAZG34noIypTOGp1QxH8+PGzVC6oCpjVKLUd/tA/M9Vudbl5
k+Qp8yrB0wKdq9RerZf+Fl6hcamGmqqFXQ+mh1fIns7rJCFHL9E1clHBezMSsBho0HrWl8/ZnQLZ
4JddQAOev5i0AG+pHRI6038Fc9iWxz1cvm24FCNzB+YPOMn5fzAMhqNxQWF72H0DBvudt1A7DAYb
aqk+p/zhDh2zT9VJosVqLQ0+Hk8FCMKWdZx0cDA4jUZUkEdwhPr8m8OQ0qJn+e9MfJSDXh9gX80K
qPW79MHmvz/AZP7VKNbji1NDMu868HnISITlcfI6HP2OdAaOOTo0O7N86cYajX8XCxBQnmdw9rTB
QSuvP2j0kWlyeNGOFk21UXEg46ka44FLQpoH9+LvJeZrKBBoht9nnlTDkKWMAzX5BeXU4KFda6qf
SzFImIIFLEW0acANwrCEYoamM4EZDt2yhVnUjGuh1JYMLQblVpcsIZywbk07mgrmo7IlkMppRUgk
Ra2qcrJC4ORL+Fbt7LhgmDFHuL2qPFuyxbVeeMxpcfzfLjuJ9bPXtzpzQxGJMH9gI0hnbyng565g
cjJBT3Vtl8JM5QBlt6kFOTnHSsHNRrW/4689ATjFdSaNN0tmTiRrKRBErF1C4HCGY1CUgbLbjyFl
6gJ3i9TTT/3yZoKpEU0ZqOy4ssqkXj9LjhJWuul6ykuRTFGegs01d4hbvsyGYIlpCGdwe/5UOhza
UNyz21JfRZDfI9S4v6bOWf5W0awBwQhRQdT6RYWpboTmxjYPojLXF59PrPmfmNvfAmX6e25Iq7rs
iWVnMPBI94VhUExBwyJ2Ri5T1LNAwQfo5EdBCSWNCR42Uz5tpqnu9F5qzjNCL3E/xUXtJ44v9W5t
b57zyrercg3/SmwL6o9k8vISsxkxlsXnDnKW6XlHw3kF6pcbsQfOnb0OI7iegwSXSfaBwpxldB5S
DsmDkdXkoLFdrRaLQWJz9aLFNEB8s/zzJqipBR3elPLxV05OwhEQgqEX9K2CkXNtTuApR9jPG2FV
M/AF7KybS5q08JRhPfio9AfGUPOLUz/9CVTJ713JZ10oR+B3W5S7G67Loh8SM2uoou4Jk+wR81UX
VaZ/a3zY4M1gkwKS8u4i6tnbVuRNERPDhvxaJv3f46U4TYdnOmY/m1A90TF/dlLYSCOKgBTGlJK6
G6f64ynTW0qdOg3HvFeqAqUbgi3fcxO9kzjnnd9EAC2fGt0mqL+Pd1H8FlT0uqUVL0AMZprQX292
KhBaLav4N+NaJSYK+q4U5yn9w408Z0PtNplTcHwTMsT4aZY5iFeRiG+aSOEWgNI/ylm84RZxVYha
ygxvDrs7OZVav8tu2iMc/pz6Ovzv4zeIo7eWBEuhCdJE+mfZnlA6kqv5mebcyPvs8CE6lKbRbgQg
gEGGLeaZfB8SqVfIWZI7x0rbytew9x6iYQATxe8ROexVgHvkry5tPXMBePaDd4yg3Ep+Hf036N0D
F+QBwRhzsi9X8lTpfYoEkk302P2qg7+Ht3Z/udejetasueg8Fu82Kpw/S1PhwuBtOT8YSIEhwHN0
G1dylYSKW8G79NDmjVJGLVB57PxsxTMStt/T1yKtmxJUK2pzG5df7I666nGixx49TnYmwI3iCcIc
CYCSGcwm+Auy9O02OKMHfJ42i3UR5+r3xO393QOK7jYFUpxlBBbQ4yhrhG7YzGYgLW5noMl6bOVs
0O94jvQGXUcAAysLkDfvbwtbdkIdN604OJnSWtWgC+1XcAJ6Ji79nimeS+7OaAAe31xCW7gCiwsX
wsDUxQdevtuwse93BRI6qIKwn1dauF/xP5Kmry1tmQdf0gpwMibd3HNV3qJNGgqvAs3ejZtQ8FMn
njxsnx01sgvKD1XWiFyB6iMHGZMwtJ7wcubhPB5zdYC7pzH50o8ajX1yOz4dEIxDaTZTJVbSRC1o
FY6cBul441ZkIhz37rTbVz+HNLHOtNqE+XTYWxwbZEnf9W6yx4T7ltHTMeA5PPRoeXyjwx0zziFu
/6ZQL6Mk4CvL87klUYfBmyUaxBTdTf5d5j33rLWPLALEW0DQUanwEu/B+wPm12heFE+bPQ5FYMn8
t+CRUH2GVhboOf60nAOegzz7wdgPCx8LHURxdU09uJq+RarUAEUverufrowBtFpg1MJ/ZfgQ+F2Q
krncgJ+Ri4y1sVm1LQEQSFphy8v1UZmg2/4ftLrDvrdZDRnkKGkGkNieP2zsL/TFzFqFYWYtbOIT
w5mmwLQJ6oTJrkwixc4BlxmG5mJZ5IUdE5pZeGMIUaRQPtbVXpTPAp1xWow+zWZK68+d0ve2bMO2
4Bng/AVJTUd5IRePJGTpAmztXU6MQGvEL8FFtYbWmUuDO94zdubXtbgVtW8JP99bmqqEIHTNaOmj
Opkk1+wM8cr3s/U9ywNHhUfcu0BI1odDvvHw8W1X8tq4IH2ll9JvaGtRAxz3YCpOnnRTmLD9cfqM
Cd02XbsNYtVVnXCpTsawmLdByVtOWc8ClbSEk1VIUCnsQzeJBUvxmyC+IVOoSvNJiz4Mlz+uDxnN
4oA3knL5wlqN3QyBzlH8ONa1dbpkMlrxQbxPIhRcfjFV0DlSdgwET1sP9yYx+0u8LDFUCy845gme
/9HQ8OoeZS9rs9xjspJbA0g/lrPlIgdsA9ggOaKuQM1x/6rGwwohB3MmAKtNhPYYpvV/u9SHlVi8
f/P/CPKmprXiu2Jot3m+jL319uy1ZjyF4BOcBYkGWGyKFvcDavwCJfqkPfjQ8J05rRTxMLUziRnA
wpd6zxmZdU0Cb8jCpVsWpz2VypkwmGXheEZZObeQlQyBrE5uubTSH2DI26kWdZLBn4AEfwSD+Cf6
/xaVoubqpylPz1knMle34NpDrhKl+1d9osIuhOQLgHec9VK21lDK8O0bM8hKCJqQAf4jv0iTYFB9
+dswATNQE9J7bR8nuwk4EYZ/uQJ70dNCkvQdKz/dOVz9RBKx6wGm46eQuaWd4xlOxjfM+6QQdViv
TS3vN12oW4gprHbP8A25+5FomwdA2xOegIkEYKDTvhsw3avh3vE0JC3TPsysVnxMfFy57ehYFSx0
Z8BWozgBCAdppX7CtrECbsLPshgXRM33PWQWRKZZCfsEUCTXudtGdLrtl90kq0g7431fdYhUYo+a
uQNA+59GqtUsBTkNU3eENwoUkmymAlaex2FR/YuaIcf8JrV14xBzWdbFWBdonZYuZC0dEUyNIo6B
t1LtUBCZ7ruodcZbXPnnXurqOqDvOyMQkfdCNw1B9YMDjL45Ckkcx4iEzJLAsapyf+Ic1xUCcIqh
nU3h9xPV99y5oBb0/3Ntr/6fysM4O93gE8AL6f1jwzS6DQj1xOaqn9FqEKXCm+5GPjldQyFOzhA9
sxTD5x4YDN8yjaOqV4kwSoZsADZmQ7w+NMfKZd02/ONNO+6xMkdkfWXSlRvUhvHY9p15OiMJNgU8
WBGjTYIWS4HL1N9Tvp+qjxswsjHo7YPpq1Tr5ED0v0rvMhw2ezFX8iqSVISKvCiSZFJAzV47JtHa
gzLzR6s9uacLHSLKHosoSNJbJSmKpbN9DNB8EfpVE5hi6LI0A0ioPqYMPfXO7V2euAwHX+f8PD+u
HHmNzGlh+mlIy0j1Ggtme+uOaPy44m//lW7ctweVQPna7CmDc/2qLDA3cMykAsiuqjOdDjgBgbtA
5laWtjBESMtB4cXmCQd0s/aBkoDXw/y9OtkYp7dpMFYJyTEVjo0I0jnH9XMlIsbOcm04xEhXw02N
qtx+DiO/I+1bmy8lHpJ+BB7h0d+8YFIu/Sh5tWm/UeDq9kP/Z2Hh16H7gx2cWhauA+s+GrNDkNRt
tbPTm7EjsXP4JU3dEy82Jdlgu0CprGdGPFvIcgkZyoWIXtA/j+iqpA9pxXvQvoyOOJe1GK7Px1Vz
O0TRvlq7AM9HnIi9aKwu3a+7W3EjkG35WfS6QjUELbJ3tXglawnm5Zi3dQtzttahPF2Chl87+YT1
NPuAw64BEWL+WejrglcZayUPbhGZqvtFOhsQjESIY6fJFJokrw6QmKn6HpxVBhpxnZZ17HiCbvcc
rAsZQnc+/rjVamSjifAyxgj+m9JfL7IAmH9kSbfzRFTj/4y5azZB08JKk2kqSRJTMZTNTEmAn3+k
K/Tb5yMOQw9IVhKGRalXHFaANOVFl/lXUttJz0qt/NWdS5tDKntQPtoKJKRkltgENcjCWDd7Oa2c
o9fQqMTYxFMrHnPGzjdDigEHxTGTAnHwiI3q4LqTDi0qASDfcYJ7peTBV5zTgUKAQlnU2a5oThlo
VOzIRX1XsVKYSSMwnsIQOQ5NNccBx/wbghYNYtMTZFOljjVrMfser1+jv0zrA+ih22sp7L1rkFNn
pnjmon46ItDePqhbqUw013l7TavpUak64OAa/K1VCmaJukWxDHhDe4BgOs3rPTN61vyGYfAcdr3M
sXz8fHdGRGiYFA5Xajbag7IpL0S9CbEmdXNJsD9vuo31Yid7LMvI71TwJBJ9SBCWXr9U+U/rknEq
zkj+wRUDlSu8AKAg/9en3EshyS8gQ/HjWMJWIfma8m7Dnm3a6K9/us+WnY6z3W/74knWcSV8+1KA
Eu4XZo3z0KMlOc1JgqIdRPxozh881nq5QQlszkaNHl7e6Zu/9VMdrkcz4ywdd7upse78M0y0fyJP
iJZz0gYgKrxDw9QqBbWGWH/poYLaf+e4iV/SkBRYlg2T4YAf11Ljdd7tfF5Pg1HrHsw0Gyqhjmym
YBGbw9aaO31GLTesHJ68EauYjjqQc8qvoQavhzMH2z4yzNwjvrqic7NLbRvXmAJfL0DCfXk5qseG
NxIkYPUBEXAxYA5I8ySn8hxkCErL9f1NA+WU5cHrpfy9ZWvsqeddD5y8C5gyFGnOJYKJ3wRULGve
AxzN7ufr3JtxcGS8imZdqnuxhW6KZqw+ToJFxXvO5uUDFP7+VioK7OFotrvTE0fFyc6GnHgDuejb
q1EW3eniZpVbvViC6TVQKUR4W2N9RqcalyEw79Cqre1jNhnZoT5FZuGTNbBYkmHDcgoqWZD944hv
Ct7LXh50BGKRAJpSjhIzW5Tk4TXjdTI8HglVlEUXSjU+f2sbevyLsV7TeGl2DfD/PaHy59UQ1n8+
K1Pw6NYNzfFTOc8ay6COTaxxSevyDPS8HOCbQFg80ZGdv8B2AeZ8IoF4HrbexnaZD96ctLuY+lab
+lImmc4uzqmRj0BH7wTXWK8J1stCLrKmH6CoUKO9ZP3Ar0AltuSig9KPAyfLXheepyhVdxfqcZUi
4hHZ41jHWPICrRI4SHBhcZJhBBxoaSSWWWtdZbIfthXNuY2sc5dZ8lHcBDp6GpEKDyWHNR5qORBI
8NNmkldjqeddrmnJJOxDREAVZmDT1VP0Tj0bm2MX9Tbch/s76JMTP/rAxDbW2jifsaFpqF6vavjY
nX6RZ8gFGsFvYlLF//bGyAdrC74jGpqgHgN9i0+M5S193qfhgOPh3ZMQHfuqwJQyeGHbkzOVN7Ri
QPCQXE4YJMVfb3DS5WDuymlMz11gNE6lwa0iOfF24xrzjdblwryKcabzllXhTGWJE94yftZ0dek/
+gVIOtsPGTuFNTjfbOrkhunMqoX8mEOrW0jjzRxlzXyKC471DeoqBLvIwt2vZ4qoAHv524ab1rey
q9aHpwZPF2mXK//jOhjs0h91UCY2Rwcdv17++Hr6hA785L7MQpyqBXNEj0VtC0DsOdrSoOB4KS10
2Y0fg0tGsH6x1pj+RsYxlwjcTVr+eLkOh53AiuY/cANMgekmSSB8i2r6o1Oa3FmH1NNSybcWiQnF
MilYuaqQhW+fJwEkgzv2T0opJmcdMe2PG9UA6QskIP0xZ1eduFml63F2LbmKKPCL6T8IHjmkR2pV
jdYSsQDu0/O2SE32sNSgw4K/inP6af8eQUTGMbfKRCB3HSgu+MINOXhUMnV4/aHgLciqCpoPJ19u
AIqYwk4zARw6GzK3NICdQUv8/7x70vu6RmGn1+gIqTAFrzC+x3mYEAZ92sMHTG5323kEBq8CCa15
TILtvhjPNKMxA0aZJs8U7qoKzB5135kTFIdCHNYvXivbWnhmyDHFLzaEswnlkQoKoe4OQbCYFfuE
j8CC6jKXcVGYW/zxaCH6kqG/TFZxj+FiuNK33xtsDpGk+3ZjejY3pRgdHL0mZxMIKVjG0gtb/bCO
XzDEYhLRlUntXPMJEgPHKg31WlfGcIUksjQ1WagflnYYejvR2SpvMH+9vJwEz9J3Hd+q29qfWYye
C/0pYNemJJJm+Eg1R92/7d8YBUlUuLz3cxf5kXgMS5xc5jUUo4cWHL4G6Zy7Lo0BC9VIxmhEhxtr
XkiT/xnpnr32VnxCZNw+7z3/8g+7qR38O89wHhkXfklBksoseB85mh7ajV6aM7wYcmbr0JacMD+c
Gk3qadDoVQUxQW/ZUFH6EyRwwsGC5HFMQ6A1jC7FK/9HZ7qqq1JN7PsStur8fkRWYG/74YHNZEU7
x8XrEu4UESb15DZvNX+iP3sxBR/jz2K+kVSTvh0uLST0ZJTlrkjAc/xxVKAQ69EheuA9EKYZC3bR
5zbhYtNcKCpUt9ef5la4TWjlvq5w2xdqwccn0mTpSE2GviWgYqAxSQ9BSOQHTTdb3xnFcii3oUd8
tLRjmF6cG3lgj38nysGsBXZjzlBI7dgKhrexEJ50byNSz4f7lV+bFhPyPJ+ELDDW2xlKwwVMUcTT
UCLDYhgzuTAAgALd1NmHPHaPxCiYvK1sI9+mAjtjnEnicblksG8E1lFErTYcmqk38RTmRwbaGIsi
+4Y6OyUKjT/n917+pNlQp0y7zhvHbwEavlcPTFHN37XwVGz0ZHDykIInex4iEcQFV57EuySlhfAe
kJCWETiN8bu8ZL2Fz8T2UmZOOd0kV0pD/nIkWix1pYdCfMv3sgUp6BlAKEjEhmVJ2tKSAaLqrtYp
RPTgPKDddpqj0ZK+gRZ7ClqNGgb/0O4wLQ6kyXdUpyS1d4NoSuY+xfhzD6Mxjq0jKK0qbxkFpRyp
mxtUpFUMJ8LqawDx65hRQ/JOPn3RUBDOUpcgNUGkV0lKMdBvrrbF9aFPlEDQJzmhUGoH2Ly3iMv+
GUc6zHfEbFwnvCJkoIXE4YElwivCQoNNqMlszFudc+OMHfmXC5owludmMQYC7W7AsCW15pqztqaL
+I9lxn1ppo4LpznjxOin4c+x/MtUuYaNXM6laDSKl3RWOjM5d/3rKtZ1+QL6N0PVP+l0gptnxVfE
YRLrZhnvkIfEdnPpb8vLBQ445UxuJNg3pc7VSF5e+4a5tQ5AY4TftYQBkbkrtHMBbwsCjGa9OWd3
o0PNqfXad/geZ1mNJX6SOeMyPY2a0feAQOGf11A2l0cQaJM8nmM3solfEN+D1Zd3fiJkA58edaXq
Rg3vy05/9EuWpyYt/LX7NBIau3uFVvHuIUFbNJvuw6c2fZcbYAjd7koDWCNFpV7ttscX8sY+FN+z
GfQe7veDtMLoTkd4uMG+7mELemLvp/IRgSyp1KVmVh9KGNBRUlN3+8V/WgAlMxDLEuNSGoQJgHrC
3YeIAG+sdFPL+Ol3DRxGvdh0Iy/2qhnDfohix0iAaIQPed5Ei7hbDZOhsPMbf4SxSrrukK65G6YB
Pu6eloIYPEEMZRcnekKnwGzhnwpIim80bou349ChPtT2Vhte/XtsLg4EKLQ2BjZ/vw6MwxhGQw4i
cJxWAc3dh5rYr7nJL6e8Koy7dPw7jbbGuOcv28kLJdZ4/Qo4EcwgsZTMlWmB/J7EOwqRw/wPeHnL
kPJ/gHQlFnVMkBH/khwxlEkxw9AE1mYUwxCF6pCZ2yACdE3+vNiNvvQPB/MOLSooFBTClRvRyrx/
2gKIx6GLeXbWbGMFZMxFqI5WkPIfFqvpJP9eID9vp+AtVB9D8A3reBwbw0rgrQHLCCB12VvcouHO
VJceWkM5IXg9gV0rrMaP0gy2TaR43S7nf2mOYamXZjj2zQuAW6K8gBBvrTy9pwZWlQZFzbLDoaBr
Fzw8VM4wRJmL+h/2Z9O2S7UaPa9FpfMVYX22SbmjXWXE74ejWb4dCesilVzaZHz4lOZ5rTwFMwAR
MVG80RXNS8/zy8zcd6kJRmCC4osSzYDvly+b9ZNZOGW37KN7EEjuVEFmiZ1ACCtB9d684P16vjp5
hxfW4XVMpbqGjrBMqMezZwHD0HjP5PiZ3NnrIboikWYI9hSZWGRNNpQRkGLi+jncvgRxvD+OcvZp
lwhSHteRT/nGbJaB8UXr6Gb10ShEuAIXeyM4S4Ax/Ew7qCq1Vm73+a3sMdJ1oCrafeoyOgRZdPMg
8Ek1th6Korw6ZwqH9hjc2779iNKnuHBvE2Khq0cGuM50yGasLLzw4exI2G0n7INnoDBjyXR1QQmU
arcHkXua0D1OlYceO+EJ3zVTrST8P+FS4jVBREZZ+GqDWkkJGznePCaSpZDkGBtJrlvqqigm1QLd
/mwNTHpWksUnNf/aCdeyF0WjVNwrdqJ2pRSRt6Zg9iTCBBVXVh7uF5tUwxBV3L8tkrL2cqOgHfzR
v26DXesaP9CfF6yZzIBblHEKZtERyt6lo6gaPAC8+S0/uFxaAU2EX6ButrWNw4XvKahBCIIbb3/Q
GUm+93qJWKI630r2UoTySQGQ0IJncB2MeHLXkWuWhxK8k9tSOkyxbZLZ0bw8U58DOar81cSAVDGN
CqSQjR23EQBAIRoI0hUZ485J4q1PyEWTQgy6MI3e48siMML5c83UenukiIwmZ0LOe8MOgAGZuT2b
fUDYsMowHdZBd+y9rE7LWFEAh0fDrlJM89ZOWboO7hCjhdHV+wBR0VmJKY8POrZNgsa155Q/p/U1
72lF4Hxe97b+jzhsKR7bXTxhgxAfr0R+TWM+hqxHjiHQIIw8w0CpDoiF1/KYyjW/1jLsWoIAQXTC
WwmdmUfVJnGUSw92cckG+1zI60BqbsB9LBk4imq0gQpxecy8WbBwpO4dTg0zHVEt6T62tKXARZDH
l9xtB/mggHMtFac3NVbMylBj6h9PdwmxF/Qv3I6UtaSZMa3sFomsdGAd3B7yCuNh4evweq4CUjJv
mJzyVkOjtDL9t1vW0GDBWNLfRL0xdx8P8qvYmUrpobbnOqpjsTu5D+87Z4wXAGwEYc8b5F6qfAzx
1yyg87OMPYJz/vciAkZEkxFJYHOdeX+JB3WI6Nx9bpkfjhMaqearvhmJOHTEm5U9/O0uotj0A6BT
lV5dDfsAZd1E0XPh1PWY6XZhZb0ePI3sMTwPw9vHcYbgJg7f7+8r0AYJNVXqz/+vOYOZRorGxPCn
GdZqTYKCqDRWMaTLAacTuOzGS2ADTzwMYDEzKheN84dmp1vd0n3KuIuGRuvJ9v6QQBNih+MG1UeE
SgkUYVhHFWhiUHlfWmgxEZPaxlLLmAjfboN+uw+Vb4hQ5uDuJZAXWBNgfL0AlW68wigpo62kdcVX
OIlArKBNJqfXssn7H97YPSTrCftdrVnRr4Eqkp+VUg0X1vVPSCRdnB31H2S0fzXJ7S/Laf3Edbcr
qu2zAqnO7Q56eJXQunt4tOGc5g0u+f2E4bSe7EKk7wwvtzWYyeLmzvFs1QqoMK1vNNq2wm9mIOC1
gOnf0qq324/7+3UFL41GccXmZPTwx5bVu3hZi6aHtM3begXngH+1cX7jV4BvZq/Xgvloljo8/UE/
VTV6No1neHJ1jxynjuHjVlt91xlzaNyNcfrmihzkDJlKCwxhpvB2GGBfBGyBXyMMkcjixQoDOZS4
79CdZvE7EK+ihtZaVaV5krqsrv7UPM2Wy7lt/WGkaiy8G3kQO1cM01pFXD2QcL4z8/EgbsbUBfXt
Ye2d0rA9ok0PFuy6S0DmCpCFhl9QtmSzF5HDFjzmxjtiLnK5SI/CQQCNNSVNSQtXNS3oPJHUx6Fu
buAg5G+dtTrFOcN2w1c4KTtj5EA6853dnv0Rf77JLXJ/fbKHN2aDYONHdQYXPkM2FC8F55FrPSsy
s+G1SnyA8C2+0LDphumxQbS1dEs/Z6EqSuugNXoclDqOK5FHsFnQ/WIaJQLsuostNIdGs+m3cg8v
i6heQupjDk5SR4mE3ac6w/uJnypJpl1Gj1XHPMP15lnZf/i83XEQZSgfEAzJovDoXKJYmbvCcJB3
cXNnKo+xj8cDTHZT00QtWTmFNC/Z/W05rAHs4P5/wyGmkdtDfQJpdnF/SsrkmU//xaN0dj5b3is9
yO0fXpeVlVw3/pQjrpf9mQ1gsE12tpSjkvQ4aZSb883HiKtGcAwik8ktwIKiO6yGdRegRYeLCvnj
E56sJw8r1Hw80c4IdXJvDJa1u9jRq/e37+rWrAbyDzKfv2ezyYJiQ1VWzS0yghhESJo3Gy5m29VE
n6r73XbKBX/Lahl6lAvRc0L5hqmkebOKCwDbUWruc8Ymt+dyJVJ4rwU2aByzyXjkX9JFJ89EyPhJ
EVVRPoeeGYcRf4gpJFcAibUaR3gGlv/dLNodROx5mPh3LJCQ1LjKMeom5u+ua0gbqmw1wcHoQcOw
PwQYgvwTY4WgWQM/fwou5RETldKpjqj4g74hmT0I2C8P4b+ve1t4DqPoZ/Z05hpDMpb0wO5bo9OA
5o8gJDVVdtxTV+Et84nVjr6gNx+PvJ6rTQK0nPKO5AOs19ccWNsEFDiGcE4W4WuPupc2JgK9i84u
9mJgU1uw0AAE9xl2dM2ShNuqgaBe/VWkUcfXWEjEdRPKUGDLlyDILsQh98HqPs265MzaYVgjtNGw
tlO2r1udnhzh3BZhNauJs93Wn8uzIcr0O2m1ug5XS90vLVCj41uG+3JGoCHQmEBBKvuHK93g7Hww
8gzvZ6n0Rwv3dgWcS0yz8bW+6YoaXS5DKBj2TiWChIHOQM0n5KjRguI2tYYf6FlVT0/29FZPexHi
EwgGo8bRLimilELFznTvPQDo5xarQg2hjQdUojxHx4pHbOufcD+MxWK8G0DkppRm3kkq746cmMJ1
xiAoa+deaW1eZQ7/4r8DxIVhmWpGYdMYyPcsumJCRfSSfMXPACKDvUKhZKAyqJFO3n9unfHvsGzB
Nqd5I7NvjONzdR9A60F30FaadXfpUzJfzXyZ4eXv1gjpmrtNDM4XL4Stww01E59KNKaTPIIeoJLi
itYUfDnGyok43j2YfxPTEpqAdy258Krub/tRip/sXMtgX+ZYdls2LWEbMQURbqxmypDNJtFHOrHO
W6GSAwL7EqdsL/fWqYhmla63EWE7p1BYBTJUBSAUBaP63sgJog4jCTQhDFkeS2bjBebfarky5zso
X/+2U0QFtOvUINLjSBbnd2Li52bFlspDRsdXZgvfHNAP/Ya21skhfuhK6XB97rsS0c8CgH73x6Kv
ELDvghu8SF6Y1DSHveNf78g5pvmvU16Rq+9LapY6MJKqaTzkjyWojslx+DGB1zBvtw9HHeVCtPA+
jCD1v13uTR6sWJDhOOAIIGQmJVqsvOKAbPr8T6P6sctL/NbmaudxLbbkcyODwQPRYO/8mmO9YTCO
Bv3GFj97Bpgn9Sswr8ULYAtjR6HwXI9IGh6u4QAUTGegb39i2K9KeFIjqiEpUL+UZYudQgO0z3MT
bmaCzLKqfuL+yCTZqisrxNDcNMf78OpKrH8i4TzvUqNL9SdZRapbzjaJzUDh5S+YqEfy54hXT5G5
++dtV4QIiGuXNr3+btm5G/qwkHj6GNf56cpxYxgMcsRigMDfyKWCNEuHX2k6SXGN1RVoOoezXHsQ
6+TcLTyE7gi9PQoerl30IYw8IWSYDOfsXD6dKocygd55rjwVQmdMTzoG9N2QV7BSnweZsqaR9+In
F1D1EWgbznHBJFEJNUE1kuT3/kt+aXEFGEJN94qDtPJpIdurhy7Tn6lrl1bE0WZS18cRijv5kxwC
Pd4si52bijcct68cZAALioFuKHESnz7ZcTw0jnoutu0irn9codxn+XIVGRe6GKJGVnyEylz6b+5o
GxK7uJi03BumYKDW9gQ/b+uW02g4VJkzdIEXsx9cum0an72sIYbCj6emMXRimKLKOC0KznP3doJO
sF+POWN4E8F6aTO4QOMptofxxhs719KpCvyhEYAVQLRGf7UMFowBBsKe1s7kRtsWSScokU5bPM3c
OTeUXS4twyv9z3y+aoy9jVYQarZeH10XzylwPFzkM9mZl1ZlmsDyenucWDK9RwbIPsArhvw3mzvC
O1jlt7xEiNMkVianWHVbdPNSoYM+pQ1bl3gVGqxjoCPMcJgQaShCxKKKAX4NSjLB5Oq3SZ1FF74S
CuHdnnhuN45ngwsQ7Rfm/GcMZ1mdy+MEB7TMUSyD5S0/uRvcDwpRoadz5+SCZK6EYbECp323s2Gl
KbUlX9yYG/IOKL23lmzLz33CC7axf+mRVTyzxsrudAYGiUs2sLSvO3czUrlon3mbDkoVOwdC7LfA
RI7l7bK5OrUd53ALTWis/Z2PCQk0bUlkgm2bIyk6QDU7vJSVyYsos0JWwRID9cYx5CQ2vKIOeXBn
3mPUolQdrXrGVEtL7g+tY+hZnx0LXlx8oEYO8iNx6/EgnhExIBgEK9xI6f9yND2cJm2fUlsEZX2P
Y7zc2e0khFhzvpgqTOuReWCX6n+EYPwrZXH6P3Nj4uXN+hBGWSl6ZD9ycGfaDnZkZ3E2urr66xE+
oYTu9IRVB2qiUMo0oUcCSQ3NFIY4XeiX+GcB0khIjkWQeu9lNLUUefL4fzabuhRrCyKi2btFK+8/
/COG0/WY7/xIqIOFWzNlNNohpOobgbeCWpqX1FL3btRVaHr3S7Fx00f+QQ/oqK1J7TWv8zpyVz8+
+3vTExo04usHA/RSN8gKVWEVGynDOqMpwCGZ3rMHlqcjGSzwdEBBHOxMEIlKGw1NVqpX5hjOBjPM
hbPKNGu43d2KKTJ74+CQzHqjmQab7PllYlvGN578GqqzLnLAlAf3vhF/7vVVPYeL1hRenpJ/RD8f
FZrCjk3HTIjluGYDpd2qF61H7F2uyHB7eQhqksXm787OK7cmI94T2Ys94sv7qrL7arn4y/+I9Rdn
9FzI1ZVccFskc0C5fEczHD53zgDSdCuk0apB2eNZGpw7ict5tjdKwA1QoDzTN8zZUDkDc5SOaEyT
WGOUaN3Dnv+DdX55CqRlLRNSLKtvvNyzFossu8vOGiYVfmO/xZVSx5ktv5smVJIYii4tECZIXQme
NJhVaGZafV4JeMs+CZDCqgWGPvIsMCXEdtxvehW/12YchO32NsvmYPmRqubjN09pEyqVOgSTtWqa
++hlnxKzFrocbUAvowpCTThX3Om0whLS/Q1w1aPLmzaaHe/YqOg6lDKsdG9wJs6ri4Cc0b1PQo7P
btFjEU0M8TtoONgseAEnLqcP4dspzRl3pEkSvcKROkCeFCIK+YyHqwm/TE2wEC2boWShEQsTISSF
iDwZCFTlGssNwczfQ8kBmLNyxJlaU9FoLhWbD25WI+WeoW6/6UUqi9SaebAVL3j1/BpJ4fAiDWJM
GHdd3JyNe9eoV4+owAxCx6UftQrbtjy7MlBYDFT6KQwNySCaaOiCa2Gdrcr6cv5PKGAPSzodG/bX
BwexV9lD9iIHKuvrIC20SlnLDA5B0GTJK+J+tvb6ieE+u1Fx8vXilUbTLqHQp36UIiXCM+ikMrzg
41EvcNA/vwBSS4ntNfFeDXjAJm9+j2Em7/IvruM/2BwHT9juLbs+ig4Q1URie+csoWL1gu8hRzmJ
vq9h4lG6+hUnM8T/Dl2Xt4S1pKsCdLjX8TgVC/mbdll7YB9XZCOENt/Z0nzKVF0zE1z4mSBem5XF
XOtPOa8hGSU41eF/lVznBp8WTB0JIi8ll+Rb1Yr+8V3CTg7cMRYMZvCqZQjBWxlbATBg7W0EMAH/
yYmLJajczEqaC3tAIi6rpvPOePxhq2YXZa35hnqrxLLY2NY0bdbe23bVr+F6mvs2aXhndGiJVqMM
yKByF+kj5IugM3D9mR9RyhWrkBqEr3N3pWtkevoRaXoUliZ5knqX+0QgzD9bSu8Lfg7rxjXnfzj8
UnjzW9mMN/tdSBWjWwBpsmzRWcg0HzdDoFDsGwyotkDhE5TsXtDqFNDxoAPeGnKPzT66KtltkfkG
o27hyoslroL0Ze83ozmBDhwh3QdifT+AtXSA4cZhMS6WdhelRHId7uSxikZursILBQD2eG5Ah5g/
7/THMwKV5GyL0s1rFwfRYGsWZ1FZXdb6gzilzGJk5QFMF7tdraF/8zPMOMOkYJekE8ff2QWWoqKu
L43m26F36JaaquvkYut+Air2Y8Z/bqfMn+8mIAwvfqnYBrMQENP3Ox8X+z2d5O9ovu8/+zkxt7C6
W2hxhxmRLe1jX3xq3pUE64kDB6UlyTZnCRKErVpwGrcCDnfeWnwivnu8ZqjjRvX2MhNCjTBehpUT
8uxfZxrTOLhmrhGBl7Rz8OQa92tCcvqa1SKNQqKcGNuBOSPN7Uchud8iubP2LD8akGOn+Zpwq/Ix
8a5ZgX9cGWW85aIZySI4Qq+vM65W9k3ROBfdd4yk67PasXAJc5EIYwRAINx+Z7auXycNX4HdvWdH
3N9zEwDVLtX8jNYmkHtDRQoPSCdnUkDdsOnG6heAlUf0KoRmP+7uHRPEUZYTI3FH8gb7qrvuNUVy
LA67Ha/50dPU8i8wOPZsoZAMJv3Gh8ESoAD6Ck6GAaXjSZa65VcJYzoEdT0TWiyeVZ7hXR+o2uzD
yT6mnWOZ5+32SUP4dObqo61+JIw+nFccbW6i4eHrzjmqk5iCSoZ9fqFzPPySWvR5gkjUDFVkBNbj
AOBS2t2t3Y4cAC3G0BDD9rPDRuL2cgPkIRvf8KN2tfVRTcxmwuG7+tc4O1dMuj+2IBXJ/u2OHyQB
4NI51ZSVPDwFbpntX++nJw54guyr9SxMgjvAIk7uvVT6lolNSRXhFujCbxt92uP/DAYfCfWlOwFt
43KxCpS0UNv9v2PT01aV/RK1FZ3/5br2ooF9NWUiYkQs+7NCbCXW/KrRCg74+orKFqy8vIXRtZJu
nwLuWjOYBaRNA+0eOIHmS8IJ//jnojEW2pnWSg11FdB8/vFzC3CoY1nz6UErVUEWzvqWlwideeW1
48vR+IpZALLwxFvB+V79gk+gjfOuEwRjyUVnMtq/cMmi+in5GmqX/J3sg0Z1nSfd2IWcBZyFv/BX
wwpDLPRfxjedZjuvaMT80x6qotU3r4H1A13YgL+7MMl9WOcfwytosONrxwsRG7/6VHzs9f38bRnc
S0ED4/Ta71GdSNDmM28sfyXwMBIiL7md6GzNKakMUrumikpDKiuso/GHxoF1JCfgv02+9g4CTspL
10ANldZxVLqWRmiF6CRlzA8XmdvvX/6QMy13M1zU+G/l5A9WijbE1e4wJgaL5haUaTAjPgf69TJO
hTEyxamt4TXxuG4mWmxY/dp/TohdNHCBYOlOiQUMWMi98wQxJA5PvU6eSo1pJ/JSgUi3WO47FHvc
fuAekVK/xsGTPix6T5fISIXdmEoPRWldVfhq95fHcOruGVskWNFymEYsMU35Yk+QcBseLNEWQLjI
UxEjD8UGdmxVYncR7h0fIebR6GMyQUv3em6ENtcB5MIAT2XOhrgxzZ22CSHitNh7zCewIr3ZnkNR
PC2qfcVx4+0Y4fgvUbt1BQviGR7txPe/ZsWE0GC/TBMkUUmEv8AJ8YFQ0bmjuHX16rfXlI1WQZmG
j/5LjOkHus+1Fo02ntqmEqn7T51p7kwBo4ZOIq9rDmxmZRbTjPGMO4bA7kxMmPi7PN62YjDuR8TM
Wkjki27LLZpqAu2+hbNgtpHBF3aWuKoMT0NyOLGjBkMjBY3HLmWfdJS4JTyGN/rzAEAIVUIMwd3q
apEj2VicS0hJrBBqeb4o3PyPmPaXE/eh/CoYN7y6SgPR6MPpsl1mYAYBilDu0xqcT1qr2KOWMZET
ELsrfyzVB/14JyoqUfhfhSbBy++6X7BHAnqlgjTIKBnr2+ZM3MGS1EBZHyNr+n1g1DxCSNHaa8Ip
dRllytnXl1abgcHAsyuDP+fnbNw61Q812THUBocibzouNMl+uuZ7Jd+MdbuVHRBATRkU6SPY3d03
hqMftAvJoe5u3ln5Reg2+PMgHUZ26YYqV+psoZEKd/MLqUvZ2lFzXMNI4WqK+XexQ6LcgYWP1wmL
tkfulHu/FQHTqmepVcMwE1HcmAos+LJoaNnsz/cxj4oFdSFmnMZZowLUVMTpGr+/LP8ud3DcPmGj
siK1i/kXEgS80SOWWswjyEItVCn0OMYnYRHfcmGx1ikSxnS4wJP4Ny0IqEe8i737PmFfUq3l8r/r
S6Q+GYkC4IiwftjO24Ep/t51uEb3fkZTEZss9VlDsXV8/6auTjRB20X/eMPBraN9BcAuGvWA2QNf
RJdFhrQmxR4N67RAF3f5jcwBsXikO2YSrLaIUADo6/XSefpr8xxYbp5BYFTZIg+m5xMpN+6xFba0
BTHSd1N1zDRKgpH6t5cpm+SKyM7MD7WiEpoq99LaYhaJJ2jKWFJeau3zcPN3GksXuX3CtdsTpk8E
ra3NNjqrPcVRA3TROuGGXXiZZgkw1aEXlr1sjTpUZViHajtmtVc0WPZ8wSaLM7drJzp8gDy+TQzR
mnV0zBe1fo17yGIrcbNgQEIP8MQDaf1ssRaE0MsaHpHzBjQUmhw6IP+pctvvAGAcSNyCoRd7158/
woQXQSvC/+6YX5jdRM6i6lgmDt76OXwoaR4v9W8MLgSx0PW1/nTrVS6YjzmkLbrxWLBK0PHnqrfR
EnRhpce36b8auWuiCxC4972sN7GLYeoEVTyviWo7yrlXAunoW85XKtS4VDGVyxejbmKTRfZPtvp9
ER1+TOyLZEG5PnsVo2uc7B/9zcLKh0TU5XJ8wD8omQf2zompSgO/zJ0osVWx1M6X52cmEEVst7VR
CfMocbZQoR5nqSgAPWrQOYD7Uf27tr1PF1UmhMFbm/EN42KiN35vAuu6wfo5psUXT/6Jvx6b07K7
q951hrNUZbElL16lHS9g0DqYM9CRxzjK0+Scv3pDHaVRU8QS3j7s/tswCgCNe/vku2paWclrqF5U
XTp2sPV/3wMESBSg4eopCnxMMQQom07dvp2qU1xu9dmBCrtWEE0e33NX6IlKz2Kux5ECDHjLm9H8
lcpmen6Z1W6crWvwyozZdYX+BHoWbpJZrsj/zyVqJFUpQtrBmNHSnCBmxx+kg1MrRDj0KW3eMB2K
InGsbLBS7vyZpUSBuc6SDpqilLXJEJ3YIrc1YfUB5DtnGPM3ewFyuAJuKpliHm4vfGwYSibCeq2k
shFJV/rB8zRGMvw67Hmubp2MjuQndHk0mh/Qb5UXgC39R8DXPLvWgkyutkC4su7sS7XgiB5CrULj
VpO/C8lcFO2ThO16KRsHzh31pB0N1D679VOlHwmRkZwiiBgDjb4FqLoF1cTTtE6FwbPZ8sW0SMcp
PIKiQ2LphHXxOQFtp24vsmIvdyXnR0kLT9WAFw4469qolhDBQxAQ+dh58gaUyf2zaZSVzPTL2VIu
xNRyvAgqyA+88Z6mV8TKcW+Na3SNhwbOK9CrhC8eiXk+8L0GT5ntClgXI/Z8n2S2P4nJJgIwxkFa
oB+n01cENagpYOocHs66Bw81UMUJa+WPQwvxd+gl9hNQJFo2Qjyw1oIHexFejjNwQyRhyr/MeDG4
U2JsSDxk/23N8ETxs3BoCxOOWpbDHXZjbFb6bmZ4SSsRBis6JFNcr6RxgyUMd5rYDbl3CIIecIGu
eUtM/xzkR/BT0ja22DZbJ6A26O8CL2P+EvAHMTvDHz7niKXB6sPNpjpJ7S5pms/APPasVicuM2Zu
mYRHolMqzmmmZ3U2QUfSJ0OIA0B+KI1ViPXtrTinY++nnqSf7qmdSUhqVbMW7qg1ulo5w9/A1mWF
+cftXB37RKq7PRrQiT+kxSXC36bPEWnIgYr1AghTmWt8+YfYJ4SvUVMopOYMBe+v3slxJJzJQUVX
v9Y5eb2AMulUzwuqqBiy0vkiIsz7B8rbDqcZazA5SMv1fcsYR5oRQGmAmytO1KK59aGDu7zOD5Qe
Lwu+yOG2vtQ+x7cTLGnH1FPWk3K5SsvBIkcreCBlJRe02J4R/c7au79YWHMoogb9xr6LYDB0ndRv
NoRTlKxnM+o7evny4hMMwq3ZQH3v4rHX6xf6kwIcJfyjI0j1O7Z0NUyQC54sIa8UMk3mJLidZauO
7OWlRx3KKQPkvW9OYLPknG1NSAMhZRlLRa8YRXFC4yR+pH5tRSLBd8Sl6BkBahxhi+OA8GTT8gke
kTzAYYMUxvtMRZHrQqMoQ/bVMZ/mpJMPbi8cTluie0jjcPHojmHNEhDjmNuOHu5OZnaMb5eOOcux
MhKmP+d3rW4DK+cErYLKHMR9HyyWVx7SX2SnSJa9IrgEAOPSCditunnEdCuo+1QyDbxLa6p2GzL4
0mtcg4RKIG9jANFv/6kprH8mwXPZ8keZVrlKcnEx8XosmdIJmyRqehs/0H0l7TP4s0FqB+OWZ+9v
cN0FL+dARG0M26hd7lWQrqZf5IZAuNuHXqjCE/k2VkbtXHXUkaFv+63d5sNi6668Vq0O+XJK7DT5
oYnhgR/nz4pxjGylbpcQnYu4c1CL64m1G6JNXl1DVUzOGni3EnGVeZkdcybJ2XyfcGqQ6XOoMgOT
oK8F/ZiNESbE48SRftQxgcoIidXQEG7nPb7nvWdpdosz1enLOjw29M9/zT0eMjNXhKVJ0xba0UWf
/wf5DhMi/AlCXsbmHgpXKi1kJKzJDQsWSCArzumBKxtBHiPwcD4WRkZFKh689ADpm9oIxqTRcdPe
kMYltU3IFu2ZFZtyekmmZ9cftQULxLN2Y8Ik6sU/C8JG/ktjk3czfucw5E5SGs55OGSBiJPTQMoi
LT6sh7LVFAOsexdUvpHnrKoeVgL1Jt8Jhousrag8xiRTHkaX3go8msvfz3wvP++fbVL5huCnu92u
XoonbN0npihJ0VLDKSbUS4GnMPE7Ae5IuK/Su+Vsof+4NbW8ky46WK9aQRVeiOZ+3fAJthi3VISf
GvUUDVBdYekrBTx7xW58KdhR4T5iIcGMbPtxrUIjwaAwn2fTKCJQ/8oJey16SppE7XlK9QPgYRii
D+4szB5IGrqDhZpX5w25G+sajLw98yeSFKuvWsW1aBoj8C010+91+gnRW8/qj+HWNa874zVlWhiI
1XsUcz0OObmVucD/y3bUG9OgKu7zQyAoVjvuXsoTOe/+ylwpvAq4KcvuAKIQwJkDPpDL2r/pGD44
ldvHt3wPJ1E4LmJDch84XvLcFA+EVfklxUgJsKCKestKLT6fbtZcuZcUzHN+N/GZSEcuzxHeR4kh
dGMuxHX4zGQm7uFV7ddLCbzt8dqYsuTKLw+OzezHZB/U03leCgio+qY1F8PN6+cz7voDqGgQh8O+
pxcc9aPoBcI6KBCb4gia5O+vD5WrVAioiPgeFBBc27b27jF5eSYYYAvgXzL61/B8ZGpfFW1MfH96
rfhxsT8l19vNq+5H8OTGEOBHDOScQmPGD6RaCaysqLHmRsFogOB3TJ3lqXxUwMCIE00KTDUdCcj+
imGHvhnzlHEg4MGrZEyNacw/d4TnhTr3NAyqk2LcPizeFeO+sTHvmEq8j3bJbUPtAjKCZiuVX0p0
9N5uXFQ8qZWbmcW4qfevJqSJluBACo0MgMtaipzSrz6SXQFwtnnUHf8ajgYTjOs5bZuB7TZ6vgN0
lf3cwP/7P5hylFRnv4oSW78UAnoALWMjSjp3WJ+r+R0Sc5NkHY1CoNqUyZ3NyFe4aHULzU3qURxi
uB/lfv4HL01RAtkLf4iptMqfJ0PpJjSkRCRMepXATC6PfnFgsKq3+G8hap+qEDeR3KPilwWkHXmi
WXOu+fgC79YyZSuJ4Y/Iez99K1A0Ne7dfdDhKZhWn1lteOQKuxyh2g+VMRJ4K4qGiuPgYgZD14fA
UjFsMFaj34MjtzAfNBLnYd2KKOXobAlvmxycR1c0SuJD3Da2z5VHM68fw8vicNQ5/aHzPpOsY81k
yqnVXke7KQCfPS37TaQlwiYE5CC7BZaso427mhdhQ5OtI98M3vvz41XYGgxVRBDgJmrKPBQcz6jA
gkjxksQS5SgdFCpUpN/1aGEZ4CNBRayzw1mXD7O6uZokFYmnZ27MhrObyjljxq+wSRrEWcUqNmVj
xFWaGgNhRMx/lQmP9B4LwX7LAek9YvYfgfVfohD3K3rsd00eaW+AGQlxKcQDqHGcRhO9axldH6vD
cz/WjMhLVboRDVqGC0jV7mappc5641ycz9ekwzVmX9a1fYgGyiYNSbePevQ7d/vMwetVhyPjGrrp
JOrwF6FnhbYEC0bY+VmRjBnS99qLuLZIGCPUln27IL84cavfeRAHcAqEIFMTN/wx1ti8MVnje2zk
QfbwIHewyuyBmnTYldzvH8f2qK3a7msDc5gYMGhPZK41iwnSBMXOdRIthfeVC3bBlIlv3u8Oz8gR
VDnONjO469c8Ck5CVdIbdABr7+vpaasEmkrygEWzGbybgd5isJGYmgreU1bvj4Km46vvalNTU0wQ
iWINi2ismWN1xu7VzSwNaC11T3ABnP07NA1M1CzfFWapmyUZp0KHb0dRwazA2xJ9P7QYRI612UTc
aD0gPvDt0tuxQdq+zJ4AolV5hjuIkVoaIWFOqAvWgWUhbcFHMmrT7LSzsByEyc759GjIYqKmK8JF
90+rfSMiIbAQd2cpiKYe8dRwi9YWn9b/oV3phjrvgXcT48feDg3pysUfo6FT67ZdUDf4Pdml+AmR
Lua0idX8kWVVcRcuu00DIzCmGCPq8uwMN3Od7KCwKser6eNRkW9VmEbcgttRoa7iu4hb8tQhlnMs
gSzzQU2AMZhcXVTWrm/2MKd2pavzbPayxSr7tDjV9txQ0zXpZH43vURiM/AL8w+YxLMgbH3SJdS5
wzpKMZKjTZrXv2uH8rlfWpADLgqWlnSpARPQU4LglvGfxtMspGsNDHSP1545G9dDe6UTT2/DyoCW
HZgxrre8s5qE2zPo9996rmwhEucVk03LGeBARoVS5oXKbmYFPtjKdhgyDjGkp7UoMI9i0VXdCTti
m8M24CuxOmqvf5YGgpoWNfdFaL+bRRz5oOl9V8tfceaPbhPzkZLPRFQCnA8+4uXFcgKR29RAIwV8
nobBlQ5AMm60tfiLbeHJTem7r340BSowiUVwFdLhy1r79G2qi95PZEgG2yFUNBeLzqeWo6xFqvbK
4RdUjrqqRlkouety4SoTUnf4TK5TEe3g/y+Xf3ojJwtYmrg1EmkIeChyHNJq32yV0iPMZHAIthlJ
KpJW8ZmB5gUdry7W9aLUGpCDuwQI/bpr/IWYYsJsgsGnGNv/vxTic4QwgWUpYc61suHklVSK1wlh
ooufhvaQWLSlPhcin5RZlNC8jlROxXfiOouXUOz2UvFLTSuCJsa6/pvBOJ1OA6X0SxTtI0iGJ4zl
6X+YSN4EubEVebBGgtUX9KiRk3+rIG3FdBustHVSI10dm+1kltINSaUq4MJ67ZxlJUcwZVNG44tN
wOue2KuAMSQmOz45/Caiz2RP1LoP1rzKvdm9UVaoZ6ClicIJv6I7hYuE/72DlhN4/+EwksS/V2Gl
cg+whbcg1qCCCaIrQzh0Q9IOucB3Ysk322X0IlnNU9tPD1yvg2k0t1QHseJJPmpf6upUdBJNbvRH
9h64eDYzH2EvQvUXUj2oWIffq9CdRq6Lk/43fqHwmhmKLQzYIY1UQ1s0gWoVsPBQ6FfqB3UVipb9
uehZW6212O4d541kAGiRjzRa3cIUozlwZnUJjjqHD4eoES9F7uq84yupqlCmmoJJxhhSPNcPK500
+I2VQddxbVS+r4PwRunMsZ2AQ+RChUUjKXnbMRn0uSF0EPe1ccHAh/jY6yRKM7SXHvPUq1YADMf7
68nqyh1NvfUDfgHodfFm+7CfUgOHwpdOZ7Dl69HFeVvCpb3GhhJ8TYeb2gJAxyO10c1CyHzPiiGH
73QbvltNFFhe+8RXaa8j6Vw1eChKLI+W9mIZFK2PbvVvp8SkN8ZVb7q9ebt+B7UeGNXS68NB8MHd
Rr27IpHBxF/wTWWUzgzxiPelYxVGkIyjlh6rYhjNM6/bxwvkgih3qVc95Ik2J6Y0QyKDOYliPEIx
cib+sIPOAIYhfedWfkTtTXaE/s66RaAXtTDsesrqv5CNWu7wjfL6V71AcG6uiolTuj+T8Gz+Wywa
5Y0D64P/Yd+VZrH8ccWfCIQaOsIR4YWW6HtZur5bVJso5t65A2gxpdunVvvk2YsqsM023iD7CD2c
LVuFADFU1Z6cyQYtUhpqq/OmuU1eXRPoHHxo0HSDb4z7HE7LPG243U+9cUfHFoeVd8+bGgEF1jNq
lSGq8qGMBvF+aytQWfn/z7SkDDH05Wfr/dnUr3GBaIYIBGi13IbziVIjC4oRFqY/E2XG+3j8DmwT
ra3gy+H+19o+CNpaILqSD5udXvTtgCeXVltpvTRxwV15Ja4DYMVlg4SxcVoEAA2VNkt3czr3Ji9n
pPZ/bkJ5B01XrX1eiBeNga3geHBu30zAfpXD+AmXr96vSdonyYfad/dCXkUyTVCCXTZpjsYQu7Tt
5Jacui2M2kYySTmDKEp+E4FIx++AmsQ+APCpR6mDAF/iFjzLcph4oBXriZNZcFP07rVH76N6Q8Sv
P0llnBh8BSfWh9MjFkPve6wtox1xvFLlVrUsAxD+tUYX5vyn02PEWG2oqaapvbA0gO5A8CL8cOau
JuWaiCDRObjCXX8eMgHccAfQpmjYeT2GHaCYR4FWQKF1B1+I+6mJVX/Ex3E2RecVPX7nLYmnUHWb
MBOCoD5zquTQkR1hE3UF8DKrvYbIl12YFKTiaqEOZWaZHIXkad3oa0O0SGFZAHWeHeP4LnovvPYO
dacuy0lkvY9DzLJlcITJPihTscAOVgUjSoshQGNlf8QDqpkNJ+M3+/kg8njUgtSYre4YfuNlSWey
SCS6cVwmhFv6Q60Ne89Zb5qU+BeOiWWNbe6B5inQZlmKgRNpvsw+EZ4CLfCc0VKAT4qfpQ6HtBjw
cUX6thfPwg84PD2I7u3qu1ohp5TpZoK6yLVepi3gQalIShp3jK/SCOy7tpM1EOBiIQ7eyULUtPpS
0PRZAPP7+rZswk1YL/kASMwAJ0ZT4Gm0j7MizkeVE/FbnvJvHT/CjXsALLquXc7CYC1ERMayEEQM
0dd+Nq9cjYNBKUupbfnja1+Zs3QOQq7oxBUTwoNtj0E59orDIOj+mGXZPf2shjBZ6KnNxmgcSFJQ
/E4sqrdwx0ppjrJzt5+jodjvE5J4S55Jzfw2Ml2yS4IeyFc/Sr4UR8dJpqF1HL5ULxH2EOooUewn
tTH2GtgMaMR4+lTDlAwW4+X9ryHMZsT2wzKHNBNKmk5/4CGIb7AiHr1ex5P+UkZ927PZqLAIpF80
CzHiT2LiXst1+go8Cw5Xr+0Vek957soSkXulu0zEmN8RdzgUJ+aR1BqutrD5nCi6CK8DXtBVEYOg
zyAPy5T+GKM6+97Lo6VCUTJfRX1wmr15y89inPHN72nIKiDzCxBh+y4N1XJhaP5rYe0y1KFwrwYA
wyxmzOJWbm8qi1noR5dfyahLStBiiy3ifcIvPc6sMlg3rOiwpESxNoCxvwa+6DFgvpjby7TXA7XE
c4NoLbo/cULIncjBks9G0IqXcYfHcnuQB+slsthHpS4ZpuxupK5HZTvLUZPMCbDsHQ3jvOo9gOfI
CLG+5UUF2oRFLXZS4LXzKu4xJNxMLvqMdx7b4hDVQPcFG4+xQNMX6ZCeMIrzNijSEhgPIF9ECC47
sYr63MocnV4pxiLjg0BKREeaNDufFKQQkEfpnAdveqRyj/LHzSu4oH89ZAeInsj+nGf1w3FasK96
qAaGsJpgzcQWCePk9lFbNPvFU8H8/a+9hpBOj3tcY5eA1C8SEdE9NDJC3g3dAUYZHT14C9MmGe+e
I3qB0vkGuLHtBVZ2T9jXX9LkZ74uQKa/nHH7QkjoZRP9hU2Nu7EpU3ceJwIe9bjTcbD22KaanDKG
IvKp1G3dASWfSXTfNXNMVPa3r+KSlr5tpeYEQ+cTxeO/2d01mxcMJJSJpaBzz3VpEq+/SaM9D1dm
xoTusPeIIXQjMJO5GpddilPL7jeIylsfUDkX9xqLkJ+OrfhEWXQ9t4D64fK2dsibRvNEYChK4lha
z1MyyBsjOLR2eT4AOEfjjAtkUpjBz8vi8lCg5KgKs3TGGcUvONtTk8+hvX2mombZxmz+NvzdtqXY
iulEBLCDGRJajisaRoSdWcRX75pC3is/bdYAVjEZH3NNQudyrdCcv6bvvs1PGzHwGNkl5kBYtnzv
rgBZ5rxzIttpZJ9th7lHCnJaO403UmBBNubrXHI/TytKax9fqDKNh82O7tZeLvBYbq4clu5WfACK
paJ2l3tKqAmWLeZXyD+MVyMdjXZuYqaK4OVg0UuOsyXv5x6Yp4posUxa2cznOSrXeDLP3RXWn6n3
C6zF6WngzCLQ2aN4zKKTCCvOlHYZH6TO/XVlUuoK3KRYmYvgqepNIyT7QAAI7OXYjc4/lxBR/7UR
hrwTlealwhwpveEEV+y3l9xolMPFMDd6/87ufgId8Pg1hruByFJvbpnr+wUECCwWZQ/aNih6xEde
q50eALR67QrR4CMoXf5Z0rYCTp5ChBU1xIL5CfxVrdWlZau+WAnN2UJ23REVb4dlM1YMhjsDtyDZ
cWpLKWflaqgQQKjSYiwTw3e04PArOJlbN5I5+Tb2MufDG9mL72JZVqS0mJDewlbpx+kMQRhxXhDA
qDygNT4BwmAO+rHxBZ/KNlu8VEWRurKQUN/hwfYYsSFRpXE3dwi7acCdjVI2WpEXXbJnvECLRpQZ
IyRT8e1jRvkRM/lCNj1fY9XqMzMf50FrvhDDyetsGrvYsUEOsiSkSCNau9tfLBRSY5fuxSykH1m0
XSwyQemITB2eKPdkg3t4fEZuPFYWPYeYqYfq96bUGebeO2Qo9XEp8/b0VCJxdZZRW3HDM9p6OvPX
rTJWfblgdZZkkv11gE4sfgE/89wNXpx0FzsTxSlzuPLS8ru6rSVMkQtYfZNCGq9adf0kOk2Z3ahu
a53Af4/k+qOMQEVJMLsTUMsiirpqd2rtISinS304EicthOWRQsAS47wxRKhuPG3L7RR2jeEvUYHP
na8FsAP6C36iemVM5jrDOwFoU+G62Bg4bxPLLP/momPqWUYa3YPRmh7cOBbmHDrm6s3UcIKW3Ky+
J9IA0aX5jyxqMMm7KYmO2wPW4amWpXOpnYS6eNauNa1R983cV0JLEQOWDrRh1EZev9Tl0JdrRrfu
toSjKjEzYMk/jri1CSdAgpxHaJpsSCGfjbNUtNAMND9UBVSnetKRiybv5gLg666JgHFAMCFUymi0
XXm5f/a/QMMCAsm8gdGARqow1K64cxGsRz//suC34d9EKQArY30OhHgtA2n7ZW91BjlTXHBWqS8A
/JHws5LGEJbcf+tHwV3vvyZPDLYyTu6XVvGtXLgbe7Nh5nxp0WG81N6Vd2Tn0NiX7nCXy/cotF4t
6ZOlv2aJbP+ft+0gVLAMV2BxAKbaTVZeJ1boKhfMdX4napp2S6q6X+phZbLjCcxMmCr9Ffv7Vya1
3m8XQqRMYf0mdlRQzcDlGFdt0Y9i1ARks8vcDAOYW1XQraAnlbyo3Ta4f0aRA7/EgU6cbrvOtSB3
7EyygjS2Z3/+BsE5IIKvY3IfFMjNWWXven7qhQPLfMBlChX13droFbmgT7MVXJm0tl566i7LML3y
zkkXkJYK+h35A2w0x0RnCj8UHsXSdXbVwKIckpL/TQaAKCfuEp73gJLVzDfC1dm7MeZ5lIB4nNSg
DYGmuQsaJyYex8KwWct9joSwQlf/XA/Bk5nFLlRRWbzmcWiQhpr9GiQcfO6oCNui61wxIGi1BACi
KH8rLtysx2C956jhoPhPWphFqKugn3J1B7/lxlJgVhT5EfclZuQHCLvK2DgJYExK2OcyPrbruFe9
YgbI/eoUvHVPvPvzGV67lh122DqXRFdiNEyTu6XIKLT1kYdx0sbyFp42B14Xifg4rhkenjtWzV2U
9mhHNH+MQUkKWW8FssZwFMgtYR865UHFYNthEz5Ns0xHR9qCCJQ6ZuDVdrQRTpT6O7rLB1W9lGRh
JPn+ZWObuikzNrLwFwOZm8Q5s5rOm04AisqPmNa5X0J6KyW6HwHl6/Q1IluUL9t4zuFu8YVCrurf
BeiUiTi6mr9GRlqvrFzq+iX8vJq5NUnkHAuRYqD8nvoaWRftWGEW1XFXURUqshoOyv1lZO7w5wjk
pyFokTZsJUqU8yltuHsmqwOKiDFvJ5h2kf4Xu6KLQ+jMdCKnL9Gk+KSbKck8kzNnBWFqTSKjNu7Y
cq3vqE8sjkxkRqoWkUG3DCGhkh54ju2EMGCptdpdLS5fDuoOmvHTNcM7eJ09ELZJY7p7TFcFMGpT
uSmQXgJQCvohE8TmZ1ll+EnS8i9z4yukazfPk3VfM32ltb5Gzt7nTW/X+m1+j4fFbAVzT3kOawll
x2VHy+wMhz7VYp5Vpf2WFXTN17Jf3lb+LjiISsV2cM1KmBfc+bjgb4RcRKS+h7+T7AkvB1MDy7fE
Wou/fc08y4xh9JzuOo7XUMQBdZPPzPH6cAruNu6ovf2Ht5h2HnMpShwza77m1nZpqHq4v5vQf0WQ
RbU1w8odpXPpJN5VGuiiNNKuielPK6aspUPjJrqIiIvLaIU1pHILDp4+yf0o2p90jCDUmT5ZlSxi
7oo/lk0tOi+JJtfPZ9rLzllbvQUbNhZc9XT6raJBQbwzA2tzhTYGepWjMO1KwyNHM33CJELz4ivL
vlQdjDGgkkpv8upVmrRv2kCnfIPJRlhyJnnbXMUIljp/nRXTkgSsGDWg6muJiy9+x4cxCVfZ488M
XBKmF5ngigPZ/kFfAw8G7h7ONCdiD3mapSYoZTdlrybmdORLzEU42kTVOh52VPivau6cPPMkYu7u
zUN9m8fCItAO/CFc0pXlo7jy4CC++5lfnL85bPZpE4H3E0aum3tfA+rLYbSOU27dmFCDtCfs7ocC
sIerrJNk+gLGzMYn8+igb/Ebsbx6uqL+qwg2oKZ3rhStPHdJBv/BR/VnJAVEgrznTIwG9S/gDoqC
ZRf6pL307hOqcj0QKPPQ8iTgqD5o/7pouDfNIaCTYAuv/ow6Yu+OCfWZ09xZUaG2GV1Hqr8CufXn
B+FlySlpZCv1SU39W3HYAfNevEudCXLdjWRxJlN/aXIO3Wj2i/QEEW5CIsIrXQh8NeUbu5dcg2Uq
gAwFMeVzaShF/e8cOtAYv9r7znqod/DZITskHfWJhR1s+1rIL5WXZ4VieoHm8UNbyBp66q/dbUo5
S+Ea2GS/oZ21+fHWxd6gQOtvZfEeLtS+y0A1dDi5ZTmpizQHa2Nn0je7o42xQY8jm3DDRLTAbf7n
0k6DEN11sXakSRqueVJV3ieT8NTJoYDVeJV+BiXvHrbgv5dAllufkjzirVLkxZ8akbOLSdYqKyW/
Uiax8/I+L/VSEUlr988HB116H85a/Thhofh781y6F/WniZYRBL6J+2/7ihWEmC7k15hww96XOijG
suJcL0/TxirX3DLiuYiiyH9iQxm0iECCiO1b/6BWt4RGTF6jqf6gJb66L5BwYHbHgz6sG+s1xMbw
UCISRU4RPwwgSi3s1uKCGTC2hyqjKF/6i6GqU+sSCDAnHZVWm3xbTqg3ofvMvd/s0FSGVhozwdwH
WbQhiA8BnKerOFx4Q861SW2XwY8hFHi6kEn1RWvy7ahWrCbyP4v5DkPajj2UVktJRTVB9Rn5nynp
aca5vjZi8couwZqL6zOpI3BVwOBdazSixgXWGu3iFf2qoFMhGRYcdc6KEyswLTn0xMvX0No+p/iw
ExsDiyntCWVL2sXQjkOQoIAHSNnorJX7jGxwSS0mXREe36bDKSBhDSdKJ1ozoOkWz75jy9Bzxm8l
RICpSnJJdcJPJNkw+onNtjm5+5XQzWzW0jk4qh7TpV+MHVUDbtblKVzmI38g5Gjg7wZfuBxCVMjz
sz7o7ixEopO8g/yDtcjhDphV6oHFXEhfRM2QAMZGyn9Rqxlii4wGrD85sdygIymKk60IGyfZO3F9
2epben93qYYjY+wTCAsb7ULdfJF2iq4M8Nojqfo5R5wOhzJaWgXrT/+x3ALMdveWOp4+TN+SgAFg
+iEUXE0Tc4g/3mNLw5eZw8FwlVyU+tqvGAXGQTshcANJpgtFnrQxjRMyhxowBeII73Y3tfFP1YYy
3nAmZ8XOxjDhl6MkM84+zv5tgHSl69DJXrdcSj4EcKXmv3RF+kuLN2r/pssVrzJvWIg+3G18YMJp
v8RIjT9nZzG0lAnTSDAxu999YL/E3FT/aDxXdaVxMfdOT1A9PW7EYzqZC4yvnHHoXlh8r9rPwfxd
lF1Rgut3OV2qsVjydQeMRcbzuLSW/kBeXOlfGN7EQMTb5HqPkfLoznBO7mRedyGzY6+CDp1QGCkR
X0P1VsO82u5JMzm/mO6Hb7RO9hJk7LsIGzyUjKmrAqyYnF3+dPvdHQQU/zAzMTdlpiIpi0oC5Xz9
AMkffkRF7umOcMs/QSyT97YoVswnav7hV/tmAzuJt1PylZx5Eiqncqz5yEo5PKCGyQuHq6pNnIiz
S7xRd2AMowUEC/a0uhbHSsYgedLUFvlJCeO6D2J6Xy/GpPJQPKidzm7W7uFbuGn8DNK4Zby0Tj6P
FD3ZKyL/5DC/sM4d4PrcLny0p+NWk4fPyk9+t2+q6zWtgI3+KilDUlvfLVJ5AJEh89exmNcX46y2
BshM8Bs0WWi8pXj5dtTewrLAY/f3DySJwz3tsM7zWTECU/+EMIjQB9qEJODhAHMuKebTuMydHChT
K2QSZqB4YoaG71h3Xa9Z5ZI4Ym5jYWFOfNy1NZv9uMZZ8u4UYikb6vjCS8Xc2OV59B8iioq9mTcd
tQj+XUxzz8wtLCjFN/2eC/vssRh+OZlEv5K6SXOS0ruLa0SC331ypSD3EAWfWG6nvqL7MishQuBC
JmCYIIEVtWMLoB2ZQ2XgBEFh5CvSPCpJOFnvXj/utyYRzY7EdFvr8XPUHU2d307ndPCps1l+8aoa
Xra94qWKaWFXaCJ7Pe9YK+E++ySzasJRZ1UO7LaYJNqNFSFW5JinmOj6Oq7FZWr9Yoduyr6Xac+7
E91IhtGv0rms4JAjEHJuO4qifcwwnA2dAYjujpST8cAX0pNmqycYrXuBIR9lXoUnJ3e8vHMoleOT
G/hXLNLJrU99Qjp6pxR/c2Svm8syIHoY5KfvDWTi4RqfpW5Rm4cV5BNe48G90+gZB6RiP2E23LF/
5+zZ2u/kG2SvHt0vpOtWYhVOjP0M/RUfWDWo6p83zTL63a3T1mjjcudbnymNghIa4m/qSHgYwLhh
qeIopv95bfNshHy/d9N3e2PMyvIfbbs2mbf85BUIbas77Vu41JkOHe8eb4hki+H8nyrTVwVSAmZu
YhCXvaULvzOJzTbCNySV0kTHAIIL1R9JxRGBtfI8wapYW7xRr7OqPw2hJ7ZFDy2h94y6uGMTLO4G
jWZjHErMyqvJ8Ps/4uVDFDKqsOEzt6aPiZyvg/qrKkevjY0aJflq344zUZiNcblsAB8xAAbVa3bc
yjVGlsSZSkxxcRmEV3X1x/LjkwYuLYWe4tU2oMftCd54QZPD/IwCCNOo3wB91k9hy5Q90oo8x8uy
q5iXa5grupRyOulAxne3ZSwMyvLJwq1EnPj3GoaZaWLSUIX5YJ1E24KYOfU5vYbVPo72a89/Szni
TGVSoHtEXnvO+CxHw5EnBS/+gIwroEPvUczFdVfsXTklrhSAt84T0hHjKzpfcIGtAodJNIs803c0
H7zYevaf6CblV1/KlzHoEfhXJxNj+COoJW6rLZDTcpyYmZu4r2ShL5Y2vFaaXXrzjAZwlXqdc/D6
0knCnw9utbY7vlT4LbFRctGW+AO4gUzqnGCqr+gEueLa/xWJgsjOEsKes8YX3ezZVLWoI15ZDyuC
3UB2Hv/BwAoRcLLltpwe6yw8hWjfL9tJuFW78Z/VeE+MFl3A3XRq9MN4bsnLgQcyidKf6n4vx2NO
JbB0V9XTdpjmwwqOqFPbqZCWJt6hfc84TuocA+8b0I2eiEzDQc41iCHkucFdcN1Hlo41ZTdV4A22
ucEmCHm/ZhUSuyfQ3X4QGdsn/7eR31jBHsfzhTXes07WK2Rv2moCsT9faXI+79jQB8C1Va3IywNV
negg0wNkMWrtGI7dYVeeOPwILspZZ4l4vGgpXYKWk8d4hPociIyN2PZ7WRXhex1qtQ8grHQlObTE
atJaWuNbJMSutLjOkkI1qRv/Su1R0BkTPBgbKD2Zbdiub2bQ1jMh0uIINvjUVn24qMk0oVUZkbDU
frzmE9JEV2DlRqmjuIBRd+y3CjY4tsKiaA9m7uCqbNZ/Fik1+KvpqHiQwqewcXdDQrqCQ9twXBbh
pE6GYfbujhhuAx9KzxxAXLPIOvScfFuA6cVQ6R8zDemqjkfjQiGaDCl09TGV5Tgi+qAQSdLXAiRl
iIKsVs+W1Jt57LIvwcLr7BCN3fGjOPO/2OahKDwMFf2VAQMxX2mzU4OikFZH/Xi29kFCc0xGnph0
QHHJ8oGfpHYh0kxcuGO0GuO30Hf4RP+l9RyFp3Cio6MXrD59qB0a8upsbh58SieIITHXZZuma/T6
f7WrLSRe/eT49lM3iMwkoYs3SXIYfU0cLDzaM0xX2uoOqR0FVOzWKeZ6j6uL33q/g7pmeyBFjGI4
fgu2TkbF9SdEnDyV3Qz1GescSQbL1280cv1AbDhH75QXTGaQ3zR7E/VK2usrdLReMmYsh+X9UaPx
A3dbg3RLdHgLe1bQgAiXqQaJKFarkeYq7MI87tpvtLXg3VCX+iykRr0IAHw7cH1ewAkJIiGr5LiH
3SVvLhvd+pNEKETvpidvbun3O2BGMDg+xe5PMRx5f5IMw6GJHitgiENBgmTu1s/vXT7SHyczRgS0
ibKuMu8ZdlND/Fq5HZg7IY+iSK0/nATAl/iKxWQR4uGHbmlqeKtfrSQt0CJphQu1Rxs3fE1yW5tP
SLjOBMAcl7MSFfJtGDSeXBUI9kOVbPo3X3rgbvN30yzSB5bmabLNtRMQahHklDuxE/7zG2HLA1P3
NefJxx/mhf+s18Y1mwHEfK2H10jFjOlZ10AKGvK/CgJc5PnLerVwcqKKVuDN8NaEqBQXKZihEpkH
+0NanputqNakkaHBdBd4dlQ0ara0kQPKTB30tg7mwyCh9UJy4g6OAG3gOe/nyJPsn+2ohBEFUpDY
qj2WZBW4DG3pLZbFMANqAhQYDzPd/RQpmuB+fe0ki6A27JmkbcsMfjonAVFVjE9mM/M4pdHuz5R7
RIRqORAZxMWDRiDZBv5QJcxZL0NohMu3j1x1Rq0KWs7YimfGAfZ1+VUMnzphaMFN87ZdFmFtdXJ3
buFjV/251Nu12Bj5cFp3kXPyy0IjFWY5HW75ZL5U2nfP401SqYyV3MDx/H46qSswsMKx7kpEgKkU
5Dvp2WECEZyb9pvBaxH2w5lQ2AvjAudqHNVG6qDcTwONTcXFWnNBmGpebWqLdZ4y4bHMIaRJBmLz
ogVS4rtgAOixww0I3/kI6Sqir8/aZEqcDg9dsmwAyQgGPFb6yj6SRf9plbA+jwq0aj/eYZuTXcAT
0XAFU6NKoZsKNlqn9X1+hWoaLPPoX4wHjOf8tutUYrpemayDn2cDKs/dhKGMif0Nr9YLloSUtLWp
4CeJKiRlJsfezfNj1v6FxLTt5jfrtQ38+JvhxmnINvYmYTkzGSncwpvOoqToRuiCG8SCDAAODJt5
Ndz8U6pOoPfBc2ZIEdjhw+3xbYp8aWAVTP3xrCo4cxh8enAc4AO5QAlcJUj4DrrIQHhujNwytrpA
T2DesNHbkPf/LRMegaRMIZS+3WVI+2s4fR8Tant71OnUqCiYr83GEXAGxJfEzijKvOxkkEbUujPs
XWG3vAvN5b8gabKPBjAFaTPx9XxXEULvyonXPsvPqD70QBZO9YYCN44UFT17qzNLUUMKH2A8rlpb
eujc2/kqgPWpdyCKnzdw8qLDb0IAP3cWcMbZierdVk28K2dlUUnt6+V3ycDGr+aT2pIchsSxCWRp
oEimfJC765gdjs4uHE6WYMVPP7OTR3gEuoqSi/Dg8h0Zi4J2FsO4pRAgg0qyIMO2IW/RwN+WiGdg
SVOARTTN5IsFJi6B/aPnzAxz1hZQUjeCNMhdUN878OmaZrzJ1mVYfTGqAvVwupnZSMzM+XpIFw4q
/oTZNA+I1yTYt4vEahpZOuRlP04SZ+D7mCI1Xz2sHy2KBMTUQXwebFrxD3YxYvuMSIm9ww1Ohjjp
YcNiXda+TzWsb7KxKmDjyJ+rNFCo11A7cRAg8dmFL086qzGNq7Tqf/e9HBI8uKzyYCYITEHWCttL
BhvibodG6AUjaO6GihEcWIXddaLDD8dZOLhjyUaaL7Oz/3G4F0Uy7lRlidZL94hHK9h2c37EVNyB
6iIExAvF6Q2+o82uxtCr8KMCQLa2YahK7xs56xydDZQDd32kAK7EzvHYbW3marThUHWFl2giZKYK
kTmD8wwzAw/jcU2NXWg5Zol8GreMdCkcPHfqIO2ojMSDppogbIxiRFvfqpCtxgL6vKgtIfqxKCsm
eSktxEbTRqIZGtuJQ8oeZ6RIGDG8x5QODpcY9NpVZbJxH5IAZwzDoQB5M8RgSnPAiEe3Bwg60HVY
YrgKZHd4TnzQtXaaRjf3vakPEG0jVKD0pHtpw24tCKaoGnBvq0lQn/cYTr8kTBb0yJdgOdyP5Gq0
AJimf1xabQWMJhBQ6lqJJDk59rvmGFlUPp6X0T0UYYLTwM9Ago0idvcbMYghkXwo9Hq4LwVebhOC
RTuHVX8eXW9fm7C0eepOuPUwnJCf3D54CRuO6/L7t+wA2NTfAnzZmKhC4zDf8nzUJzZk4gMnOjwM
KjQk3C+RxZOheOixCF6iXLQo/xG9UNYRZ1woPSkv0h9tjJemf7RcZHk778x3tbrJ5WH2jXydGZAP
CfZkQBECg+p9km44sINtUyQti8YvBceY2gyn5/7eEfnruHiMsOPLcW8CmBQ2Oam/QrnReFGCh2Jy
OibUnM5jnN/lPOTNiXYZmrUoV/BvajmGZLue0HrbUPR0NzTX6KvY7su0I376dOVT3E1X5gpSVn0r
lO2Hc9Xhq3o/R2cKJTWJKXLoUjSDt+BhQokGKWJ/XPQw0skJgRblKleL9LzLx5+ZGdl+W1/uAZ0F
xl60RqsY/wAkH/D8FCQaqFJAaHFCYFMx2OATwJADXuWsEMRnZQYjBIY1ZFxvE6hlyYs0Wj3TyYhq
4R19f4idDqyr0F4vvfG6I9YDVTNDR5tyVtZq/HvRfy0PiaEBpVXift8PwLjoV6CEtxVGRaB6tjEG
JNG5QCcvIk8oWTycbfFkwL6w+/gDlE9U/hFIXI0Oxo7sd2wEnWorTQhC/T+hqsTArkyM0PE9jUed
wU9mWC7VVpdxg1jYIqpN3eKXifaHILzMQnXuYQINYjO4E3fttm8a3L/nh4uSzC3R9S6/ku4TJ6DE
J8uTVI8SdNzY9CjLKu9s5z3Zxcd9I31MJbiO3+dv8Qy5npDShvOl/AksY82NvNf2qHQSvxDGy5Tb
/hhIZzoed03as3oZ7KK4hHCXAq8y5qNs8dlm+bv7QTDo+Q63K6D0R3cfl0/gjnIZQi9n620/9Vx1
FkSE+Os0TCSX1apR7Xd5+Gn64xWsRKtjeZ89oJYUOa9icitfiPTJ3j/tPoVvq3ZwbLCJvCBHk5sf
W8kGMSqemttxWwWzu4IcJ1CF0mNwpa0g1GOIwBSLP1utv7JIh1EiFMJAQTGlh/lLkEhIH5JyJvXe
/xQMMlL0gqBfpfyC4BSAraPpYkIrqHSSmYzAe988FJQaDIf0BKQXN4Z2RiaAfy5peFmCHPGu2Jcx
bt8OEG9i5jiIRwhIYrieRbFT611BSiQkWXaCWmYr0TauxM8TbNY8qdnEqxnnuY1wbq9bFbZhAw99
Rp9CczZ+JZdH/6YcepnGsEPzKleK1V8jLz2D7Jnyc/q9XKG82zsR3FyT8RM7tCtI18opunPLpmRx
S31YAWzKkeXf1NNNpzoC6lv7Ko10TiwyjZ9ZXI/Xr0KUYbVTzr/gSoC7aC293FcLW1erncco9KKy
Uprs+0CvdFsk4TRlsNJgPR+pdVemA2GUa/CFPVfJYslq1l81MDG+reJoHpHlicLAPvkTNjo4u1BY
LV639NqEIs+fyucPfnq981TN4qkNSZkFLfEkORpQUGOFyyrvsEGSpJ/fK8O3IL1a/Q+1vVlqJw13
qW3PcG1XOqRTurNHe4nvORfYfAnTL9NC+YIkZwNLupBjtF7RvK+bLgJ+63g/nJiRvPKx0N4t8ukc
ZBkvA4jXXhZQ+GUn/lSgP9bm2Qwuetv9mDcOKAMfqIRJntE9DIiuvpIjW0N8hYk2V9c+wSpI79mP
R3+cMkRRCwEKxOf/gn0pD5zrRR68tWoyIp1fCkUZArQBPabkWysytLHQBRO52sXX0ZVxJpNYHX0C
e6OlKKOeV1G/7PryV2sFVzWNg/JzZMVOTHGDTJpmfsSsTl8k68lnQUYRCmHKMccC1FmXbizzOTWa
o+hD4w6dosTaIdRqTnr+rEdTGsysMf9P/yJD40rmRlJQncTXX2C4lU4bXpAubt0/XftyW+Vu2Tme
Wi7RyR5uDqsfdvTz3fNsSReOKxy4YlGImXb4nrs+YHeD6NQwvNr7mz7+80rZaY1+TAfWcn/7TX8u
ZaZJnLRPV/qWorxIzyOdFw5AePC67bNjPMcI8UDragNpmleXG6jk1FloFH3AcA3ROfkqGOsMadfM
Gx2K1IW0nYI2VRME6rgBII3q5/tqPZRcye6Ou6tdanSfoqgyfG3efibn0hGcIZi6LZY6MEWQNwg8
yZ/7YluJMZHS/QUxTw5T4ojOgbLOS/UdPF3lN+/d43pQKjFHNdzpyY2dqmGhE9J3t9TX9PMsODMI
ceOexwSUu8fJDjaGqIIgLUP3mf0zjvfsXu6/6pmV64g9vPARgbEnrSyN3qnkwq1yI/tvSvQg9QgV
pUDtTNe6lhSn06RXbYOt8U4245XiRJMbxDSc0DChsJWzQ00Cwvwaf3KaW84wfFXc5aCbUurACGzM
lX7PvFOYHxkWYZHdAXYhbjqHPDzISSMDjdjaR/CW9VywLLQLfbIP2NVB4xu5flkwghJhzXOLAbpB
hSIwN9bfuFiyINsicE3HmRnnZ4A1UqJXSBMDZ4F/9yBA3ZsSXRVIgibGTdeZ6Z1qQ0uoHRuNSDXC
oAAFiy7Kf7talBP51IymY5RSnul1ggKyfdg1AbKx6oii/dRWSpslMM8nw7U46H74RWUf9t8yEphC
SflPejObNifJi7Wgs2epbW2rv7cy7p6ltp/aNn1fH1YjDDXfrvibCCvEmG874/ZmJwGlhcDUAwlG
W+MNB3XjIAX/PjOlcxg7Gef06va0Wni0eUFi5pvLeN++uoVWDIYigpeVAyNYEBCc76a49t+nSAMJ
Fhto9MxcwtCcj8iyNk9wskreN+5ceKwQMI4kzd4MHf69f8hm1aMg4hPLyVKOzqBjJV3zpqsurFI8
6HeEzE0ev6YGyY0nOnlJawq6ircSaKkvXTkUAzxeRqfUi/M0KlmGoxSviiN8FK6qXypQeojA1ebA
Dk3VJwDkQeMHWghmE4fVQ06d2KVY8i2Pmj63VyMFOwMBls0qEAuRmWUWTDg72EhGNQK90DxWJ+Ug
1H85A8DrwvbKEdh1YddOLzrac+wpZzYpPaSyQGuY0+4POowAYMKRvltLWhflaCnxOp49098Ko6Vt
ECBC/MZqx5CiYPW1xygnVZXwaZQ0JqXFl9nztktF2eIEk2h5ONnWcduvn0f3+z+aiHZMrksLChlK
VUpEjvDtsOxXsxbSBAz09q1JPK8x4jsxtbDa1Sjzf0SfRqSlSB2Jlc+1r8U+4p5s4vfkrP7fBcgR
9XCJRLjdECSHQROrtCrmBBvUrcsLmDCwdf5iaPUNAZG4etgie9GqsclPMErmp3iSdeea6/MpTL/7
9EiBDX+IpsR7sK7D/mCPm5gDP+Za56JBp9yw9Fr9cYg3WCdE0XtiGqtdUZNPZUbXf900d66m+2XN
oW5lmrbUfZ7awiay4gFC/KMbWbmUtpZyiqtV2EwObXttBdv4OKV7iHizxqlMqA73blP7vDZ6VhMR
5OfMUmTRiTEyJmmcvhwKi0oIt5GPLY7xOLuBvMZCn6YZFXTHJXn9hWgpDqMwoin0ticU913un75X
7Z51WFmuhzpOVxYGxcc9I2JprT/tyh3vJvbHfBXHlPDTI9OgU90S2KIHwTObcQnB7WJZ8TcKl5cC
tMkpPLLDPF6sblwgM76GnNZOcfqK77b9y7/RzQJotuObwd0kfW1RRVBfamBvXpc2pmUAMosTy8R2
+xJj6D2tT9GijjnVbJSSNr4la0CXK3hmDzZNRY3SgjF5BhFZbb+R5xH/lOjKtGJvhqVcTYZWrqDQ
6ztlGGV0Otcak+uLjRPRcAh3r40ltrqz6MD7cieinkz/BgremOMJQmAaqAhHNq/cX9iTX/c6WGAm
JNpIQu8T2HAGpHCco0bP7d9rdCNtNh7BSciO+IUa1qlTrZ1jJpK+btn9mIqE/nenUUGroxJ1rgAx
Emr76RLhviWX/TDkj+C7BEljD86Zx4gzoQlkMZiX9Sd3yERm8AsOrT22GlXtJyIAJ2J9LPf7C78W
HvaL6prkyYJmBo5QoWs+SkMsas2tfUzdAEbfF9hkTTO/9pU01FHjis8pZKM7AfjyCRvffQOBzZpP
CvDK5+BwHLOfpLfmwpXcyJZvNNWTsAY1AsoC2USAxVsLspiTIqo9TUsS8FyYcswVlOCM3ZAvhUrl
6Zaj97YMkdZ0AaxIpCZskBEvlitWzsxOw3S9d4KDk+dUodW6aEPzDIrYgXb3pQWsExXv+dvKbUim
e3QmqLjnvtrB+3pBFBdxRD1HxWuTkECly8VT1I8AH1wU83Q/EGyIaihJlSflF4ybR/lqYy3ahdjk
HefXBAUg0a4kw5u6HW5SbdaaxTbhCdWaTZsX77zCxl6eLqO8bOxz0j0f7E7oFEj/9RQjQUNs/rBS
lkOdFYVwaqi9HGxBOwngF2jb6H8SWJm3r3zQp3j8bxyrA/CLnO0pnxmNApMMKfxsk0DhgioT2vH6
Ti7/z4uriU+V0PHlhbFkQ13VPi3i40rTLF2mZVor/nMbGoooGpZoZ5zF+MrKdqQHd7La2gGI4ltR
IFVg1/wvp3RJ1TuDeUS2a24cqYYR5tSsGZqV4BScmtaXTYHoveorpbiONtnSPUVCEtq8n6X6Bh+q
CV9kxaUvlOKOv04FZfv6M3vrvgHG4Q6ySrQYnR2DArBaMnXkYLBLHy0DcJVwXk6mxd7LSmok5Iho
p8ib5fyWFJHJz4VVBE+V3V8IfqHS7qoAtQB861wPhRd659sfounKtz3LqBrRKDNG9v+wsgM/HfC9
KitSR6XMsZG7RexW3fqBJCgsAZfmafAXUg0IDUfPfQIUtqC9VAOF8qaZ2YE8m+F7OgvH270E+/VA
v6RoySF7HRFQrAA6gsyATNxtYW9TXoxDQTfE7JAzWI5UlQxNyI7ypbaT3sLl2CrbJdYRKUqMAhoc
uOmEOsntfrttun7SH2/91Wy68E7+spt7NFT2sr/PUvGfuCkkkX2fSADWUgQE38HdCEZXp5CtGARD
Ll3IjHp085L0uR9UT9V9qphm9u0ZaNo5MBrayaZawoEra3SpYx2JLeuxv7HiHnZcuCLNbLQCO4im
7sYvz81hzow8LfUhIoB8Ufpt3ppd93zHxZo4QDdOHW2x4jGSL5lmJEbRZwp8M5iNCreJvXms1giK
mJPOW9gjFqq9reA9pURPOP6Rlt6IYbf2T9Id++yZC0wbGwQrDvBmBFGIsyrXmX1NjsxI8wPeO27C
4qBcftU95SHl1T/WMIV+qttjyo3BQwcQ9B9gE3cW8LuvuSFg/rwIGxIJ2y/lEumMCFy2y75mwQFG
UKxUF8StM63OrH5KgFChJCG0+Mua/prK8Y0zVkn1hjLVHq89/MmoM6fPD+JhMgZ4FjU2MWRGCDqe
7BErqdTXQpALQy48Fjerlu8sKi1vNakf+2G0CLzd9MP7MwyIB14xKO2qOvjHnaGqKsFgukOEVhyf
z1FEybUoboY6UISMhYcdeccrGUeEgY3Kk3tPqNDPb/+a15kUMMH+PXSthmNcQnrotmR6l6HQ1f40
P93YIZxM2H3LuDU2BTGakPHDBw/mhSaWk6NyhHJxJlkYO4oQjLD2CdE8MByGZgWx/dSpdq3Oh2LV
6kiXX7cf38yww0B4lyRVof5IxJQ6xoWfHtnOasRD5TN136SBie91bkxqnXa6mm/BAi1q+w/+WGSy
yQc5gD8BXlQchFQATxO1SDtHG+duagYlWDOZRk0CiYZ9pUqhGpKIDjT/1BJ16UJY78/NxqOmnamS
gjr9bMOmzTtk8nOn7B6EtLCnyACReKLV73xHU+BiUTFHb3xEt41eWlrOMQLCuKb9mRe3l6WmuaV0
AMOVjqEFj0uiNNoKqCx0RaMaPKNTDXS++PG8ikVkM3OwC/3nREFAIsZ8UvjoAtBoYThlGgTHyKwC
5itjoHr0Xt7NFSceLoFpC6hJgXzYqoYaiSj2s/mQmruIxzJPMsiQnhucgxtoN5TY7AtAuzex+BNK
gcTxrteztqkioO8L2w58CxeXyNbIih3zFOFGV4I5DEZAq/fv6HA8ESIGAL0x1ly8c6gWy0VkZ5rH
kiCfgbb1PYCQ48lNTPJcM62BpidNE6hCPDigb9J+NQMfltd45ADAOCTeOBl5Q+9kOWX2KCeYc3Y2
qXXQrZ/jiJAF9puGWa+1IuozR+LxjWN5yI9DadZ388ca0kCJHrS8AwA0nrTpPLjW3R+CqiVYfD4H
0F1SBIUozINciX7BiPjxIcLcBpIIUGQm7Td6VtBHHmqyw5u8PvzlX8fjurlFHKL6wsLsRAbEkE2t
VVvjsR678WE+XRAj2T3q307QGayNoTgvUuzV4uJ+3wTZn+vE7SYScgTEOyJE8L8+E5oxuAKzEMMj
O3EoJQ8oju8GFliDjTAyK075r1zRgUihbG5FRAHcjGSg10y9VA7fSXdUQFr+uNEEWuM0ykeKvLD7
0FgAq/S7975pOHLq+kV4q9qwe4aUuYFpKIcJKVA2tNgmNWlLB/2n/Spk8Xnj4xYydCq6QN0bZq8y
4YoO7JCr39XGKDWKFxOE6bRX8IPkfKPHGIi5L081yYAg2vVw2HCtvTVCkeWKD8Aj6os12CB55sYQ
xDBmDMw6EbroTymhai01VqkN3+pLHCmMcx4ash8dc9XrSsuwCmM+mZdsBrF8q1Szo/4LfmRKuAdp
QaQoLMmem/r7FcHGNbe0eymWNnQGt6h9j+gF9TXRFFVEZI1lWVb8fMD4a/0g45NaRgm/RK+T+AV3
mEJ5w/msMbZ0Yq2gojp8w8ZTim1YKou5EJzjez5TsoSqJqLAGnIL4ced58p3tjt1z2xOHTTG1HTh
6rYFhsuzBMm3d4hMHkFpJLTmFeg0wAs3EEa9EZ9FuGycWFkqFOJgKeSZDVlPDnrsaEv6bLXdBCgG
vrnUia585gxHzJ4rSfX2h1DZLKyDjtei4S5qxbN/wMxJdSD+JalXaDKt8M/l8GXDkpbIj76Fz4dx
ArKmiPQWslfIRSkb+wbcMJjr0oLOmMeLPyo55dWaiLQRYODGn/6Mzf2a4LqC3ElNTbfZpnmhyw56
ANKKdppqV4WWfl9PJLKpivj90FiwPo6Ye7HiyrW7CNqKKtJ8abeW164IDPomTWF3Y6FIcX2fvqqm
kK7L1SddUg3cTwKNWgmD+tDGqbB20D0P9FMk0s42M4L9w7cGvcyKjv84lWtE5yRkJ9GzDOR9J+pU
gNSYCfDJfTi8rPJ/7LcK/zW95bO9RisnspD1K9+hzOaqdix/BBLdIoiSS/n67EUEL9b3ONWHpoW5
2KfKyvFtpyYgtkF6/xGYOI3Z7JYOmXkLFS9kGxxxAktTm48XZuBwFmnsN20DSAXeJVBM6dUAMmya
kseOiOgJoIxq7iU6W+ICV6I5uRca1chP7TxR6BwX38CxXkUkwaXPmxunnqCTFWZjpbvwpZ7F/QmS
b7Aefvl7ojQWKkbUetNLYtYzD+a5WNt52SaYqo0zYtYZy+pd6B7VDUUN9w/Dnjm1tIz9QAzdmYO5
Df9BUlFvVpeRwJKIdS0k4blKE64hEbDDCxrrUm8VNlDNaQGrfUL3so0BoY9Oy0V0aQAnTJ9wY2x5
veOswWBfWKdWQL9bCaw9RjJEVeotmwb7NekDgUYMMFHG2WwSatRWaX1iPqA9qx2EmfDUa7ezDn1D
sq+IcciBhWBallxFhBoz1HHM7T+HzIcr/+joBMiV5qNwQn643bcYoGTEJWMM4ahvlfNsTtPKK/0T
oomJHdNmjnj7E2caQkcYyDRbCqsnuYpnzPI21qyjE9AmqvKioZTqfPiIWEgymb0ZlfmEJs47gNoY
ITFFjMkgvbXcrCPeRJbrCaPBFj0PEISYveoIbwxE1fSbfGRQcOII8eiytWn9sck/yXHU7QCfh4Za
RXsVF837yE0umYOGFO+p9vhQVf/d+1oZiRZozzo76P4u+ECisyNTebBK0TgYW8feUwM2gLkXfzT5
ok1t1R3VvHv6IEeepY1rMsYGIr24fjm+4w10onFTtxl7givNIBZnir0yCShmlY2MW2R1pJnQyLKx
uTvdifW+MMdGWm+vY7t957Fm0aSrskQW+dOsvXYxK0plY4aYzZNy45FDBFaKBEM45tdGE50XyXR4
NimPkDNr7sjGa91aPBih3WO81FMN65MoYPyuH6LsciLNGyiDLb2T+2/xcd3RR3zQH8LnCFcipNW0
xnJEf7fRYBf/1XN6jUqsuVA9eHD+gtDElqqqjpNF2dKnpx0NUzChW+JNWSTRKmxx2ckms1G00a+g
tY1nNfFzT2PXv5TLd8+ERqndSB0UZXWAw4Alckc/tlNlIA5qFfnkC9gOztrbCOK9d8+FbzQxw4zY
MpprGE+3IQHb+otWpD6zuZxqCSufh6+JPZflLAhrkHoBY7jLaUJDal75nHNjLKskVPwPS90P1zFy
hvj2kqD8/Ki9QCdZ7j72efsPBdGIWyTPvGWnyOPupWVI7njwa3c/ySpu/xlUJYOwCT0a6wJrqgqq
0Bk1Z1oiTb29lDW4RNeGw1fzB374IRiIgVyc9FNa9J8PUWguaZ5mXUGJBH2Dux6CWGCfSMcFOmgy
8aO4QtBwnlBp9b4zFz8q56+o8mKKNA2wG9YRT/AXbnyX7KeiO9Kv/nJutRM7wBuXLhXQZUWE8Qno
Hm5EqM6VgYgVhAuFd0qV5Kr/NTp524Ct6dfa5jbjAved/p2Q1zpySXJIU4WelePR8tdDWgDl7ggU
GkQSneCb5j5FNQc60vET5wfIv5cvZPy8VBJCxUIQcanOXyLhxES4UYa2wMIv+ODUuva5ASSQsgfy
R/i/iRbuC6pIVBtCfWdlpPE/x88kMrh9AZynVgooQZeM5B7PpkWXRZjRdkYtlpUGGmPEUDwgAjEH
ProbY1upmg0bhRQqDVY5/XUVBz8kL1+mEEjl4C2XM/qEnv62+3S9FiQ2yTP27hDoiTvF84uLgGBE
rMXnTzNnIk28afC9xPK+DS/EoTujPt9IzqMAuocVKqyXPjMdF4zIBfOVeefNwKc+Ecg/e89nEsww
CcoOHPbOqCH1YI6nAfpPGqBYiDSymxxWlsYafqsllmXdxEhrqkczb9big/HCHO2HVrSEiaen5L7u
lSgerOi9nZtqW4/MgiRuLWb7JzsThBGnaLWMC5KEHHZWaxLELK0OC7zXSYR8q5NPhddeNtXJgChh
P30Dcc0vstmyzJ9mQLYWcAS1m0GsYwFDGF6FzYtu23/5Cye2rUp/dOo48iCWgOnvr+EtEuTeIFRl
N40XzXqgSZqt45cgN8GUcAh+uBJuB/6QhdhnybSWb2WNBB3GFi82b3R4BxIliM7LaLWFIyGsEedF
++0V5kG47h+5vRbfrHWtNlyvXgtvZ0Eq4UeeZzTO6AuAR4yskxC/1eAn2cRQpRkVF2jvgsHrT90L
4yOvvNZg2jaEQOGAie5lWLMSDMhANntazbLJCQ3qR+H9NwRy4QPgTLjUNKNVzvzS4stNmXqgI8t4
U7j2KvQjXwknQKMPQH/WxEMAlRPLNfMxhT6qAQ5aFo+3cubxHaEZak7goMhNEyqDaOtDnvI/6JFt
UsAD852ALXHhfYfZ97/Ov+G4rrii02/C06nkecLT2fV6fKN3FxtDogHUkLcrf0iW6faMremGyCW6
oMAmL2W+k89abzvPv15Ru/9jbouhGrElLBDzwWpY8Iv4hsGurRQFrJd+zClC3KOCZyTQypOlNZER
RPhRJuDQaadRtval4tcD5zi54ap0BEm6mmlmFLWMekD6/sSivJTBf7QDa4eM2y8cSuMs4xZ4sho8
GFLhLIhrBFKRdtRu4Zj1Pqne70lnvtKSjHqa7AHs86aZ8QCY6AzdGbpBZHgslctThId8deaDfzh/
rD6Ywf7eCjE97a1bObm3tMWesOuEDsvHIVNScI3qDciE/2E/Y3Ptirfm1Lq5qzYa3KeigVXxON2B
D3WDslgtzEWH0XMGutVS/RKUhcfHTjmgwEVBFVzs/iYz6MuYYEfbbTDPtLKSplAf+G7xWyxsp7VO
CpDuKb5e2zAzQXeIOL6Zy4FVyJokjcz2jlf1q3EmQV+TCUcL0XuyHVD4HQE25TPleum8yZmbzmEd
jhzZDbLsA16KxnVqfcnLOjPWQxinhW0ElSOMO/UUosDmGVZvZ16yoEZ9g8igdst+1L3qz476XSnj
1FrIRIU6mr2vSpcL+7vEwX+uYVArE4/3pYEeApFXw8vgWX8n5U1mfvuQzJEOpmPrVZ6jF2G/byti
pTpwcVT1DFyMJUZqLZ1SkiHuuiVDYVHUuaZxTxIL/k61BrwQ7PfqX1ZL2fgyY613ZNFSLRrB/qmm
QDmpqa50L8kKYjbhmmk7p7k9JtmHgsO40xbVYc0O8ypmiMHu/P+7ZO49M397UQHC7lYaTNiL15rS
1PuDQIEts7bedUVLznYjclwFnsSarXTpe0oW48iglM09Q6WRuqoJAIWNrHpYB35Bu4h/e24DQlC/
p7IMg8F2DPcVabE49kjjb4ZFanj3Llj60cUbPV7ZD4HHb2b1Ow+sdvZ8oDqbIHnxFDrJo+/zg/F8
Pq9348TJPe5rnPXjrH6pI+T2hrnFDrThbC33KuXlJJHcZydAwwD24uEN/YP35NbNieLt2jJnwiHA
lHTtNHp8cZFxO0z6lRmA2rkD8CxZUooXMrtKVLOzW71lVn1YiZPkUcYRyd5FPxJWGPJBo1abpxmW
ZxnCQ9WGA6NSBqghN6M7vSXwj5Y3xuhqf/h56CICTeAJjNesI9h3nhyvk06SmsLTaHShPbHc2X3L
FfIgSkq9v65dCjIDDBMV7xxZ7TAwpFzBKUB+BY4Qy+iE4WrU0j6BGe+FuUfs4pDELE+wG+0iqP9g
7od4XLbY4UFe7GxM56Gjx7v/5cqFjvdRdeljCZHG5JAobd3Kewr8yeVtaHkax65YeNtY+TnIeM2S
suEc082Fo+51TK+YQHPGfDWDxwwxC0RoiINcKXMOZg2+ypjvJzmsL7h49HGZTwE6SD449OBclfK6
pEA1FSX0njYNkOL3qHTY2NF65Wv5gCenk4vvrI+mAK209nalQpStWJqZqmaLtspXcGY7yuHD6d+c
VUQ3zbZB6adsEVCXVCnOrEHI2xL3Ts7kMTVRUdH6yovyx5IGtzst3A5vl3BKKPb3neYx8Nj6UErt
t2FAn/kb4X2FnVF758s3TsU8h3hFJXgwXUD1vOjDmbgFddAvMMidA7QFmzpYHVtyhS6rrqhdfGeP
sKFwehK+brGx6InlHodkR5eXODFKr2pesp7UQ2ySXbrC11pFEAT/vU6EG8YzGVUQKpFyGLfkE6sY
0MFug+SINszO4LuUj/ZeGYlCMbodxfsDaw801aUUe+tTU5DnwIfMvVK8Ni65Yj6f1gLwhNDdrWAD
ReKJ9zOeUFnb0fumJVKX8/2JYGjGR2LkwQ6y84p1Bfia/elAptfguNPUFDzt7cKcW7YQS1t+uGQ3
5q87AZrsDBoRsKCqyfLK3SxcrCzn7W4XPyq7nbut8L5mraoKDqiirqspHu7MBS9K9uPcKF7EGUXE
d5lkjd3wnG6GD0JaCO51GBI5R7WPboCgXSW+pFNeLblSH/BYJC0IV9vY1TeNiHvSkXSYBzwN6enm
KIkiHMZFhEmVuCeLnWL08xEPa/t4gJgladPT57biXTKN+zcvFDezX9lkf5JMKxWq3OLFyq0BXmkt
kdx/xzRC6+PhFsGxw7m13eZYqUmroXfJKhrMrstfbeOwCZHqUdMc/tUd8jpdfop5IgEzX6jmegDW
QiQ72LjgPQSUxfHMCBoqMkNQZMjCWhaoxBurR/QFCcFH0t1lWyAYNqHrv18sSHER6mCWkgp0FDHJ
Z1AvDBpzap2tSVfscPCyIUA9eauTZJp2ZgLc0PXAckwO9sOstNJKyegMJxVZZ/plR9q0Vv43aWHY
9LJdpz4Nbkk7QXWRCs3/8gKpSdKGhcR9ZaW4n6s6UDNgkzNoduraU6xv20tNYDR4vMqWBttYe1Kq
RdlXvoWlQuTyKZZyHPinv/AQMXz4cbaJ+m7oS0O6yQ1Js8KKp3FIiTeLyod1joL3geRmknSFfZ8l
0OCR9tmelo+qHINoC1wEtYpr2tvusHSD9kHtbLnz18+KLCxZTnOT12+8dr5MF6OgokfvDdAfzZhD
nHp0toIq4oaVBPvuCbTioP1YqD4e+BNepAeKa00WjrY1pAFUINezGnjecgr8hzx0WzKV1IsLSJL9
5dKSvMDQ82mgrs9zJjv5MIrITI2RvP0fPva7A+DsatHzHWEum1m3Cw1qY/pUYlFTT6NRtDkSq/5P
Eq8W7Egl51TiSPMHbcgb9A2EdVjS50jVKqJBZ1VJ5EDczTCVKBNKtHBTVxEIB5THEGvXJLe2LumK
/cuW19cFA91sjMUhDjvWhY2FYrJR1f8wwwg6uqjL2broDMev0NOYpDUiVxkq73CyRjGQlah1Otb8
5aQ8PGHLJjZwjtNgJmCTpVfMSFjj5bOfCPRV9QdWutvotrWG997nVe7mzkFZf8yAUVNxaQv8ZFVR
aDPlgvC24RHGJOQNtJxxBNrIsqwpBHv1LYdy9g/j6Hqcbji3TC+P10B+neWUuCwaoNeqhYwxbPeR
DiQ68oowUD3d6sKRGxWBuFzcYssnxDQUCnZ3zxOimbadYR0JXd8JYv4/zNS1+KL7lG2opGBvVaQ7
sgPLNLmCA9dTsTbf8bmQxVvqMzvcDGmqX0KhTcu6fnUjLOYrDwAPMLud7j/LMCj9cfaj9A/R/VaR
y5JQ8J5Ba3XYsB5Vwty/Hxrx8xpB3X/rGvnL3UiA4nS+8mVbHO/71RH2Hk3xiGwZ2fvF2wt68ao9
YoNaDHzNv5NafXsnJcQNUqx2Bv9jZbe1tA5TmPlLiZuH03zbNjKmfP9o3jSMYLugeP5op/00vfqJ
etuYP4DSow/ZV4tUxKZQGBEKtBISo6IUNSrOAwImNmKwucQMvodj6Huir7mhai1AwRoTe7zaUd5J
Omwz5edgbFaMZC6xqi3bwMDEu1msV2zQYFPx+2vbFLx6QuxyjC+pnJQyCE3w5/aGnu2G/CZI+F8X
2O0ujSNrn7/nwBEVVmFBIYjQ4QE+4IuyTRw2zokFAzOSkC6hj+KGnzgVmFpQtXTgqDRrVrFaV4PL
RLkO335WkIcpWq07ti6SmwkOFs0+8HiI5Cc4W0RHN/DGJJ0WfRW7SrDWA4nnS7QKhhuaQpx9JH2I
7r6JtYNa5e/6Yl+4QH1Jh5Ju/Fm7t+Sk3bYvwiYNDw6hBAH7AgrsQi8blwMcKE6CJr07mRGs2RzR
TVvHsZDzzkQE36SvtUVX8x4HQ2IbUVXf8h0dOJB1jye9mmBmZmDixsuIIvQ1jidiaJN1MMiSHko8
kM2tXQoZ6fiP+o3q1yxxqbSO3fUFGtNSY4Sf9CJoYm/k0UeEzIePR+sEq6B918KnHonwCurdDSuI
9WgMIvNN9dbhOouW99Vdgd9Sh10AYhasjNFHAlzmMOVj7RCh9QUGrR1GqBoUFWKwn6aZwO+ONd5l
CHQzxXeNqSxrG0F2t2eeXcPTfAkOvHUKZ5evyhaarq2C8MfMjnn5El5EQiGjkibqLqoNCmDy3OC7
2wwBLUekb+5P8/oh34M0QV4N80W79Erfv3FGTCQfWJL1mXcPNtfweUcFkrHUoij4xiJcUkKHrpRd
AxqD+kDMmev5cZZ/WHgL6jxhmuLVC1+hynwqu4cjNjiSh1C2i0YHL/NytMrMFG3QHvW3FsdOILhW
XDdB1SQ5y6TppG8bMHeP7KIk0oDqILrbYUk2ORSZ7MUdkKTNASZMm0XK1x/6bPpPmakbVvQOgmwu
ADiILoCkKxLe4UiVGr6rCKpx+1ZcWI/Cljj020wgbiJUuI5YHR0knL1kJtkdFi/OpBgQ/U4aWLsx
bX3yuKcAttItccBNZryEohXxibDHpRN7knZ/a1zk9K761brfeq77xD/xCX5faBMfSBKDSZf/MT24
2SDpJvl1cI9nJD6NA/gzQiDqtkFBswr/agHnj1K+0RAoFv1yfrH0d7xjwMziaNgQBXUl3/tr7abq
RIWYP7ESjx4UoSxwjgjdpNtVm8vO3DyUKk43ddnvhSXaRFO8rY2TfrRzc5PNqJy2+2cCszvkF0vv
U7Hxeb+o5dJnVqOuUH2b2Iv2LaMjBOD62QVRVJr+9Wr/szfFZFE9gN1+i3sWJzHZpWYn6Ows2sEE
Q3M6WgynC0VM66LQUxm36YYX4n2GIQsQOLPI2/3B5vW/NT5tSW+w9AAWLzc7NPM237+KiutSlvOI
JLDK0EnIUuy4DF4jqeZvuLTipUC92Jgp3TQt1mh4oPt7hH9UulU3OC930QZj6u4C8WCbm+8aDD+5
MBSFI6dCI02neB8+gLSWu2yQUQmTaKnXsKXaQV8eLxMK6yeayEeZvRX9eahjWiB1o90AiISK620X
453Hb6g24nMH56BCXT4Zg+XhEd9LCiCCtIslptOvftLduTqEJCiSYbLo5D5BJ3dYrsbVdeAbKMAd
l+I2Lh3KPAfDmkPngS4NmvWpffxC7Rf/KcIOuEw5aQBlk2UfPATAJkIQNC3LOS7/QR1GixQxoGMH
vcrQUDD/MskXaFbpOPBMrc75jOS9UivuK29LmvOnpHF3QVAhQjUlGfKtiIgMFu3UBRkqAuzRwLO4
fSYqMOoAumvyz6JWLcOV9+4A1+syF4j01gk/AhxGAnfGaLywtPr4iRH8R0ju8eEHl6VGgpIhMR3l
ac1B51LtuVTqj2cUNhIsucY5UsQ6+dW4l7+N2hFc4Yif34Euu+JI+CCp1lSMJ9fPOZOicORnrlLA
qPfCB9UUkASnnMo8blNMsQT0v8RqSK10stwfXqbRSR0/e2dXOU/5s+opr0K7oJxdnHNTNCl9yilT
x2AHdF9aqX+zS3gVkElH63JeA9veEHthOjAYu1OZyg90nMiuf5Hvqw9l0VH+3nyxHKMvuZFtMUuX
mawDrqTduxLMTG9VSq7kCSu5lxMu7GHdMfFD9T2SDI34qlh8zx5il1ETQI6g/AijY8dBu321dxCl
jB9U1gI4pO/K8r8ZeOBvoApcKNXeuUaxQyre5GXTzlJjJIsRrZSzSrSQ+C0LaKyXh1DQOtpdvmrt
iJCCBizXyrYnzVtDtOAqHxtUSnk6dRYYAoOMeIlnj+1PTHA/mBL/r7eKY0M0ry6Tge5rZ/ikigx+
JOvtzLuE3E9iMX90baZkDW6fB82+kAWYo0u40oe1XAL5MchKlwxXcDnRQi/TI7G75+Ds25WXaFd9
OiTidqbQe5czo8pFYpBcvzKJ4RnsCF5UxncejPGWsKnEc6gR9mradMNseFZ3yQg5N7SRvN7xxOpl
51Vct++HmGBypy7eVOMhILWK2CHCdXntDOCKOjsSDEDP+JEQiTb5oms/FZ2w2DAB1fuhHwyUdT5J
C2fZjJkY4+wrcNbo2tx3+k/c//5dPur1bzJlZndeDfD6Me8C8H6oreXKXjM2g3wZuVoOrpM4ygsa
fdAmgeHa6mmXdalZrRjoP7beL+2f6GlT9MTCLmqCmIAf+mejWXNlj2nceSHTYEoIGM6kwk2pDJZY
TwaFyIC/ukCIneULuN1kenwcIPBlKJaLzF/Blt6c7Sgm7ACbN86QZC9bzskCssiomTsgBhj4uTFe
c8ZeDkqNudjWqxzaKATYNMGoRXyGmdH3RVcGPlhmawjGcWzGPLMHKJqXmKuCwWuGg2VHngb0zf3z
osu68dce649VqSPscB0QYM3ptpg9BHMRJiwGsmMUYC7fwI34zJXd3+i0t7ytyBx2SvQoYoHx6yMG
//V7Tw0xO1Z6rdW4bgOIRyifPbTnAmmhEVBdAW1IzvBynS761cdgBPFEohjbCQuADTCzNJ0rj/CL
7dd7W0CJzbj6OR5cQ1FZPGX9mTBQy4i0+jpzQzNrKjssp0j6S+PYotDqGLA2hvakZsBIu5Y9oZC3
mNwe/eso0CeaDTra2m06fOAuCWD2JzWoxF4DyRkTYx3e+MoKK3bxvLPXt3hmAXKjq1ZdUKw7yz/Q
kKwtBxgzgSM43TZbhYnTaJJfddkvuHrOWGmgvFJ0o9PfLk3JidkOzClI7x/WLb7hTb+CE3yGj4dW
wnuQ/plgsX83duFgrgwBoJKN9zY8jiDZYltrEcc/tyupwlHi/674So1YAqqlZCYYG1R2qtB0fLhX
oUcDg8PSpVNaTmAu4XW3LQRpVaNk5r44QQmILlsyPS7f9Shp9qv8S0ukjL0oAsaCK5yVQW9KqsUW
hHRbzX+r02z5NrabNlweMcvr07rCAss9htW/2I28onwp4MdKLvNV27GbhyVaHAfanhNLopwgAIS1
p+1Pc5zoXzl7HBpu26UjUn1RUf3YxLdSmrvEcwarBE8eNnoLDqMtqguKFkRSgqg/9S1/y7YV1xa4
pUNp7cmNTLGby6pMYtBCs+nei2bSEJ3AFvJ/lGDe3Mi1E8tshRQlN6ta6jquzbXNoOBgy25qkHaz
o3x6I141y97quwTFaZFaXi2GRd1SS7voFZ+KXMjjnf6ROBeRNj2PUCLQ+i6Y9q6AC6uTF8GrdauB
56HRWYQAOvu3nOT/4sXxaEayiiptipy5PcQeOTWaH54lYa6PAg9LPthU+Yzz/DCKgQ9/W9uE4tM8
FurMhy8t2re7RTgouX69SaeWzHHcKWDZsVMmk+KTqZnYWReEx95mkUnU1DBmaciAIfd0AaxQ7Ivg
5G2Azc1ApLgTajV70kh9yUjj/8Ph9b4Rpxt413wqs847Mh6RyP2xK/4C6h9ku1JQSIgi9a52GHdW
pzrEXnz9YvuHfAbWCAKdVUxF3cb0Xn6ZgpsTGmGR6UQ8PDZgxIZURy3zxlip0I/tp0socmbYLmzd
5cOJIUX1eQ54x/pCDXpF8t0Bkl3n+QN4Ju0CgvDzsnO2UnmqvmT6ADIJtnBeM6wAfR1liGOdn5n7
5/8O4Y5dadLCdb+yoFQNGlhBJTZZ9uGB85l9fO+aJNkjtfLVKIZGtseyJvnnmBtYxjXdVeOKjBdd
7zAOOZeRJlysBWSFkInk0jo2I79UiWTP4aLzo2m2IwzWD6TXZRevmwOREsZY5gmF1DlprVNjjq0d
pKe26+PGyLp2H7GI+MRsx4WQFqmGvq2BOsTwnHeW+tJ+bb9vuzGVt5ZrxaavlWu7wom+GLbbp4WQ
HCO8KsvFaF27kLWijPbG+aKeWQ8XgWlc5f73YkrJGav2wIcEMFKHRRNitIpZic6jNi7aHS0eHpkn
eXWLCjlpHaERRJdle+tvUH0fIZY+NOYIRX6dxxPmhl7EQn5GKEkIcMl9+o0yV6v4pFf8+kZJhTk/
XpwMnVfmMY0C2m4bdQDA+45CS5V3gaph6AHHiUe8lrLGfnjPlx40Tc7UXFe7rCXvEd9Yx69QTIWC
pmUJrJtvBUoUmDwn5ALygUqWVyoAt6hLr0Jqf2lczpoHs+8g8C1vvN3dHtzeWurImWB9xvvqS/eH
nO5H7XpDUCraPiI6cMnTaOI5cTWK7pbuHqixfTq53Ikg2FsGn5TVYeQgBOq6msez2YwS/KiiKJum
99FrRGNX+LrvMIsD8eEX+Gbipuj0Y/G4Nu+y8CytNu9j2g0rQadJsjD5vlDW0ztv5IzGyPrusLGh
Mlq09XmdsTxdIsy2Wlw7SfPvsIswa+8srvJiuH3LRx46TgaDlyWKUEvDzB+pQNGibknVnsKsWdaE
K4dvTm1Xm7lpfcYi4DYqVX7DTdCQesdUNH07YUzau96sP1IT6xnYnA2BKllNTyqER2kCjJWluKZg
2lxcW6jxQOSAW5cWuKun/tBhNFbQcdqtpaIKaKZi6nu+GlzPIY7Np8p3YfCCfvbT9Zx5wTaejp10
SHj+XPBJlrkxra10LV0BhXLqft6uGFtfcuo6slYgJOfB3nJehXLDvzY9BOaV4LlUlP3hUjK33PIN
Z68pQBprOH3d0wINIUPegEUzyX7jc49mF+Enu/s6YKmA41eTK4IjRqFZiSsrqzldMdJfnRKJdXCx
bYj7j0Zp7reLMe9FLCaIjiBtGNQbO5RYudgZMGa/fP+XHC2WMwO3i+9uyd2Gh9on1SO0oZSFqnLI
XWZchbJ2/9OgOvsBfB2yEwaC+sKdbRUmHpOZ8sDnq3ZFKV0KzS3GbXXGkd8iJxjKapIekEq4ilO7
ElI3TTlv40g3WCsom6nrN1a5Dy68Xnm5REu9FtacCtkycbr3NiOIi9EhSJOnk5ewEdL15lzO47Ac
1EbnPYGffJb0UcpRmlvGhrdgIqNOBVyqKtukhB3pZKWbpOTnkiKgJcU4/hYD+VzXsMmmFGBIT3t5
oAuOj5Ig/xS8K3ZfcY7i1YiIdV5f1QKDzZyjVf6eG7GirTbHtx39nQOwV0yNNzNNODmJL5wSCzSD
To8b0OXq+aQBD3TjWlvhRz/5ESTp20Iz9gva7y3gqkK4bi7gNH7cSP7kXmbrPtAk4aMCLNJXiR5D
fkRLh5jmNe33RAHtlgJcqhUtRXZo2RgsoEjo47gGkkfMPqpf/0nYGiiNmuZZcWxcBx9z+cxoMn1E
04IdlMzeUVdAsw7lvLMHMIwOkWqdQ+d3ZWBogrkOansUNg3dIGtva6GJpr8rWz7KWNeuRepFkfIn
+pu9DNjK8R45IwLjdYv2ViuAW1SZIUjrH6UheuulxdvsuffykiBVqh7vEWIpZuCYy3tfjx9YBwQ9
iHQ8xaCLiGAAEg2iaqy6Lgqn+ypc04syJ/nu/e7po82tvw45JxOsgCAo0T5r0YFTFBC+a+DVlpZo
ecxuvE/2XpGhOMvF0yNwTqrvY/RgMliQ4AdZKHJG8bivfxoI46E4+tWsttRW2lnX67ViFU8QG+G6
0nS+9RQN2nFaAVyPxF780YlYL90E0T/N8kq3/5r169KPOV/TMkXllfJv7ug41FkstWTWcCfYLTeo
DtBpGwBHhYn4uqhBLLwWgQTl1WDx8FDwpP2ksJJhLmdXF4l2+G+Uyxy1MzjF5uK9y6EdHYnCupuX
p7AnuWNIsUnrqwhC/EIHSl6Am/ArPca+VVOz/NEepuTAAKX/fKbdfB2s13jfzqBFiRB6kRX5v5ZY
CeU/KF4lB4LFqvHZz6X28XUltyUPeFltjavrk9Y4+Ar0A9nLQpyNzoAGcKldb0Rfxn21Vy64q0nE
uHkFvXvY/1+j5So8cFmqZKyCt8f8iCgDP0j3RTkWAz8ii4prOxN0te4qCWvnX0QSWE6Fd5wSIs0R
Q7kvLHrxdV5foHfZgNYezp8ESOjonF4MsELrxC6ylNqboETvrQ/EEaCiJt5aou0HICewVb/hJxHi
6nKwBF+8KwZZ6oBymsyhaRI8IWXqCw9mXaDR1WWsPfsuTyTMZGl9oIo8fg3bBuUY2f8s8Ij15GzS
+OcL3hNVaHIou8a6pa0sokk5l3yy+1kerzvwyU6N11He3eORhyvbWHqkrzyel4GJpXtJAWqvBgn9
nquKG7E0tmany3enDm9glbyBORVcIkr8/FDWE3kxmwTPv6E3Lf6bSLUU6xJH5M+HkGOrkvB6jGNm
95K2tRE1J2kG5rX3K8pLAAkTKZdLG1YaY1H5rJfansx/uR1xk1YauWKcVPxrxYyqMDe/Xg45jewa
49gnxcjuEQkIpGoHHEEOnaFg1i5TYUJK78OYkzrzo2nVi0C5x7vyJnl5wHPauW38CrCjdWhItT/0
OXvTkIaAEv/VToRRvHi6DRNwThEsfsOzK5AvklJ5uRzHWpIb6p5ews7U47cX7bBzbPk5DJ3+aApT
TkuHUCYp57s08SS4mJz87tLIbHrF7gYtRYt5k42akVBtex9SX3JpSRNI7BGpOybgragFE8ATun4m
VktCQ5tGzNGhUgB7opnghBUaOh54orsZ7Xc4OjorvkN0MdLON4WWgEGIWJZQjyWu56hU60gN0VEj
QGMVJKQkL37PUVGTMbvYbDuYwBrO03XaULiYGnLwkGDhOEpzLMFbeB/Uu5I+GbZ4cpQTt6H3B/7C
KlZXM42II7iLXviVVaNh4tXr+j48RCzIYFB1/pcD2cBFYrYz4WZ1DZnOoTfC2bowDG45qAzzeh8f
Geim4iJai59EvlMeIDbGj4SgQAgNBBcIPPwX8NCqHEz0XGHNFsiNydE+kUaw4MRjb31q/+TdQ4cf
NjswDgb25t66ib22AgJ0mI2HgHouYMQ0GfbqUTQAsCG0CzSbnEPTNzWB97UnNvDgKNUxrXNkm/ob
6vv6giiCOmM0MnJMo4llItof09pOLf/3046Am0M2IT9rnlqQ/a55//6FhGjY7hZjpRypnMIHSS1A
EEQ5hdx5dHpK8yP2Y//V0hCtaifZEHIF4sM4P7gJxVhJc3fRHa8E2oPJ5UibaMOaZRLpcJrFkDA8
JLuVjWafdWDRyZxL/aDDN+jiO9dgc+JM0vmRf5F+VHsNUqso10tbXB68CxFa2xNoIV6EhLAzSD92
OwBgncnDsNfLMWk7Pbpn607TLHk3F8DvFJpVEM72QvciIgtFwlH5obIy28sBA9PI8QJHu5yjFDjh
t36612O0/E+u6pc5OOhLolBk15lBigQ3zyAGSErSObCGo3AQ/J9y9V1IICohWt3MZ+d9z1gjD8DA
Wccdv48Wwe28LCzhJowwn1EQWoQGoZEInscmHz76HHaE7AfAzNKWrvQisF4xmSyiuZ9gCMmu/yol
AIKKOX0ArFIgaY+lhm6NXJQABEb3aE0of1AFqOOPpkUaKBnrZyA/Rf6d2k0xnfrLutLJ9mopHd6t
7Bu0zbKjn0AFTnMA7UCEKL/l+mhF9Z65OqzESgdv5Nfl5YYxDKYp40mNTt06JGYfhHBME2O6+pcx
eVs8tx4EqvrEVPYf5UdTaH3xwe15jKZUqrSH36mNUsghLfByIFHqIgfiIunUuC2taFDvI6Je8QtG
Q46Dl9E1ppk0Cp5ZYuO6+R8kR2mMXLUTpbUlMGvOiBdhfmVm4xawgZkUMQdouHduckrhe/m2p8sI
FbLgV1iwBL02y0kJGfNLocwoDc88txn6BcIGe2A4lLyuymMUlqagm30dfMaDMMTwlPIlqCE1yHIC
S0FWGh/amSIsSPOh1L42aX+lSzeokBkTe/wtHnNC3wZsHZCm6mbyfrhy/RNNjI3BQ+rbcS+Pg9Dh
86qWAe8NVr3wBSopiunEyd3WMae6FteT1NvsVCtunQSubdfbPxbl4Kp3ZijAFWKb4SruFyY57g8D
4mrveePB8VbtD5Fwt/HZs9CeTTGEPD8KUyHNqp04ox6zT1I4RkFIFR6bfx+D/OzOqbxMLDrO8YpG
myuBoV1428L4imXRLvcF8R8865KmVqiIfe2AXIY5Q65dXwmpUJmpycb7xUwMEYRHnrF5fqnhDFxG
Xnx4SMpO0LB/RkpqfgVbB5NinUUg72Z6YzqojS8k4A9ChTM0LuMlJzMXgOYb2R6SAphacYcwSrng
0oLxJjqkSNp71dQnd4a7MkwhgyqmA0hi3t33iORos6STrjLQ5elk36lz1EU17VYO6PWAH+/a+6Mk
xRZX+MkQkQLkcr/w+GaLlI+Ta/Z0/pR4lVi7MUGhttYmJ9aNn8JOaz2q8OmNQRtIIfSpOtWSnjog
xE4tSpgolcJV4ZxvyMHJKt7nGXZ5GG3VcaNGpAkkOabFi9zprNf9kNqCzQeL4bFenKwUWXg/YEQJ
IlXwslrLrlNREOGxijgcthIBqsM0wxQPsEVHstZBE49U9sc8upp77zGMbSleSV/IiIC2/o7q84HM
Rf1sMT+drA0s1vp/0C7d7wD1p2rKdwH2imWrABsfjI5HanC6BZEHxJPGoDQWf9mNhBaGPHuo9BHh
UZU5GoD8vaLLtK9CVNB3e5P+WxJfp6FZukTrPxXtZpxaMU/79m6gCtIbYTDrEadX8S03UkjPmaHW
gjD1jySjw6YilW2ddD8Rtxkpog3K+oVGALZR4N01/uEuRty6yq7sKMCR0XAo03eI+72ODrEsk/DV
7hgnw3HU0o2saJJnn/sLdlYNI5iHWq1e2fQ1Y4WeQ2dRbisCDta864MREvGw8QnRCc7AaJ80wVMe
7QWH7gmPI7MYdSXdWDBY0pd3VrMenCysZl13qqmeBjYexb7TtBVCvZw0eX4s69Ikwml0zwhnboIQ
c1DrYhyZYA6x7dXwILKp5Jx9ZZZMk7o/xX+4weuntrbucxprPrvDZnIEtUfIYexNvz644MUFq5IE
kJnQY+w+79HOuRFqngamqw2Cdz6FBLNs/n2TJFUuie75gRAscsklqGrOYqIxAV6jaGq8r9jhnJV7
/ACTIluzEZs8eailQiWQpeoTnMMSY8qqe9kyCP/5MC0Gfwu96EiLoc8AgaHyj8CviowgekC9LfPd
PyYy2mrjMGh2c39FHcO6UC4Q4jPGkJpNIjfsXX1EE9EkyxMeRdB1atVDy1rCbloxbQ9TWyyVvuKS
+dFB00gvfMOIQ6hn4ydc2s8GHyTLVMQEhe/QB5QElV4biWDB2AolHxUokpHv2N4A3ka6zDHMR/t6
gHmr0wgEIcbsFHYsHqJiA41pgAA88kOp3RqS+0M5rzIFJqkKy4yaVdr8D1XHID8QD47SELHzC6rE
i+NYx+smFvmy8m3EH6iRwSK4GWR14qsIJRzpA6LUMGQiv4EU+5vErdC6XdOl1vyE/IacEwfaCEjf
EdfKWqv0rsPG16X06GhBuQnYcnqfqbtDaDkabcFUZzEVxzY1y1ICAJ4Ti4IElnCaxVNAquuBGqgo
HT3W76Sr7O9uxDI+9zwjxS8nBAfAUz2qgrzkbYt5DBZihNdQ5UkPAVpL1heaynfxwU1hDnlMt7Rl
dij3nNOzcOOTcoRTx3yfpWfPlBsfYGy3zWoxLOSWUlQBVmfpVM3z3jR2x+SA/7WPyRGjYLg4+0W5
8CnXrTCqGgqfvnHf4Ckr8SbyWcM4MUfiTXK5u+S/Gk1f+iulL4jJbwqimdD0V4Kc0o9huyc1nOFx
E4YwRVmgdXbBEhS4mO+668559lXcomwKR+rKnLieBubbUByJ7yB4qQXjb/nb7pWxpf6NKbx7E6pY
x1vYBXYzvD+aSipUnNIelLaxH0sc0G+xvHCuVFSyyYQRCO6nCA9614lXZwdbjeCvjKe6ibU8Hwiu
QC2hfhyUTd0Ek/w9fwcnvxoy4LeGjDOFpQHc1JzYwRfVCZBWrAcVLdwDLzCTViTq1BPJrznMd/Qp
gL8bbuqxK/I7AuotmzlNZ08KCi8ocawkmBpvgpWS5jmizB47NI7oxyIyadLeFrR4yQOnEcsey7k4
EZP8Whz5iDRW64CF0cnd7zzft6miU+gyIDD7XPbQj2DVOaxidk/Lir2gzFeRJYdBlnouE/dmjdv3
S+c1aKYqIEYAM3IkNUBIE+w+1J/XVVqfC0R89HCwJdzaBAXKxSViK/Jj3XMs58RmfRS8EgF5/eDY
3F7WYG/DYqmPa6yW1yM1NxgeMZYD3HKvqUa0X71n9p9gGhHmZMv7BHG0JvCwuunHAzlEc7d8Shr7
tSdR2O3cn3SJqx/qucSXhDZydErOtvyBcX1c8SZ0rVhfJVVxVkyF7jIsX3YwKoSWe2aNt19LOqax
SvCVZQExsWKjqn++KC+NgGl2CBOhzHcPeZvh0HIriwMOXhCGl8QwGjyasD1dPX98iJdnu7wEC9cf
0WixUSaJgXcRZ25Iu8QclXlMZ5JOEtTTV9ZZj3sQ13D+6ESa464VPlu2buzfi2SKCxmr3QWGgjlc
GjjdX6S3i+FUD/4mH4j7LRd+XoCl6Bng/F8ynqWUYbn9yoXLRQwr+40cxAbClf/X9gysQM13luem
GvM6UY9ae7qZK0FJjOQqkQPoHVve4adwte4867NW/kBE8JEgsCWM8qb2qMirpI3AmcRvhGyj16yt
S1Tew2W7bEoTKEDuts7G8Er5ZYoY9BWqlWvlCplD1pdRx2AoFXfKbMNtx4h4PTBVsfQHIfi4sgu1
Bn0NNpJcJxYv6qAuE0fmnCItgAjZo0nupIFRRMlo6yOGl87Mb428hD/AXmEaPD3MNrSzPknjGL1h
yMxf+YcUSf2avtdFVKra6KlcKDt8FZEwp9wrBFVRvJgQ9onuEimZu0oml5aEz2ndQlJvmrkUmiqS
ZYS1uRjUf87C11b+9b3NjInBbkePVqUJBpuM4W8ujfOP9TRfeHGOclt/7MvhWE0Yg1TThmxBh3m/
yAt7xLo1kzF5PUEWKQ4aPtGXNtx5YVLHPaY24DQacy7dmzLRY50eDjt+9cOq0ZfDHMWA2TNzrykY
bEauvzO4/uSshEI95H1n0yvY2jy5s6tDYfXYiMoTlWuyxjlLwB4405bncPtp5H8prwYFuHeukV3z
APoBVHs16tmg6tjQip32HI+lLPd7AIAeUjauknUSMjHdPoCwXzrIhxwKWV8Fflzq+yTDMxukftT8
4l6JhvZjc1fsMirKFc1kw0rN1A+XKX0O/5/gJ7uimBVEmzC7jWAYqoHbrwf3DKWYvlLBGYniH3zV
RswbApwPkkQ6xHih05imd3AvVrtnyGaobU4YGStAS1XnC1IH9z1fjH/jmgSF5Gjht8jjBeAgdJsY
SWAS7Zr6sped3nsOMSU2/rbVa1jFAP5QzLzlckAZDE6KssgiVPdsM60HHy73zogZ6P8QL2W/iZbf
xubVotkAaMbnwI12QIvOamYatO8L8Px+6uxipiKgF+Vg+NPJrTFmSiR/MEY9V5rezsDoeVKuU+Xg
L7D5kAhTK0zTAxxwseAk8E1DBI1VM+NNjInwgdERR8qyDKxnIha4TTBbq+n7hRSbpr+mTtVB+2Ht
E1Rv2yczNdOaP8INye4mchaN3GhwIS5lhug6pNY4k2OPhotkITD+i/qgMRVo5ABHF+X+czRlUMSx
BYxkROJOCyKjnztzSXKBsXQ3VtmNGQWv+toI8F4Yzl2avyOaMTEhv6zyE0+CDRuka1LjnLxGO+hB
ONgdoy2Js2FjLX6cGvtmFAMSXqjp2T0aUknpPozYXuPwT7CkNwZyw8Mxlf33Fp67Ugg4FfAHndx7
aPTjX3N+b3vmZHAIojdWkIJIovsPM5vg8lVXREk2NxXH6TLuLtiU6+jf2EqjJyZvlyAE+ls0YW+m
F4kDmbWEMIjiS/9JhGbZNY3w9VCrlq7PvZoIbyerzaN4DeBPJWGpsZndGlznIVrY52W/ZCp4WSSk
xOAkzH8N7RCriQ93jlQ71W7P8/tebsVoMwSglewUbfaStzm8rXG2RX3XBo/PsiYp5K8okKDO0ptU
dOPlsRmMoTQkHKgXwPnVs4phvLlXRgxi/MhxbU6Vf1BjV3cVjIrtFAflOUSG1tU78gJppA/D1es3
pfQP++inLON1/cL84r8J8jiiU4pIOoq6sVAUrgFpzlIc3MZ/1GZAWUbNC6rPFW+MNJrwsvoD48cg
furd8Ggaz4fIrI5qrcUQ5OtjqCqpeQM4tMVw4Lx2tOuW7EpB1QIQDvZSdx2sZEsofiHlTa3ozwTP
z6scqhwqZS5lIPUBu1JyAwcucgmc8G4CD1IwnToscQ4yZCzNg9jSRO+/Rab5nWyibQaK6uGX761d
O8jlQmDO1Wu8u/vTmZqDrzOQIQK+UJku2jkjiwSOggcdgZGruapyS8GQ5Nl6WpwiSyUc5LBeJK4F
pu//9IPrzenP9/fYS9ofEIQErNmWqsMiLqwBmwh/hFHurktY+1HwxQKeFykhtsFu/4gBJKyOeId0
xsbD5B4H3IuRiyGlIS0asCZOyWTnz9jPfUpMRa4isnpWwad2jEK/EjNKay54qVXu13y+S+E9CIvB
BHVm2sJ2O8T/O594619tUCmO6aKpot9jnSDUlFI5GyCzMTHXwHsjJzzltiTwF5jej3h53ayOiMKK
QOrYweizCFkxeoy+3hbvCxtAeJBQ0tW3QehocUmKCR6MXf+fUhe9CAHt+RSAb0NaRlpuudfJfi9T
jycYtoJpRBfeuW9SozONDShzGom0FlniSAc50ZyaXwx59bcjSzb1x4+9dauACCK+57SlHSuQ1KI4
MXIdvFiwlOdVGXEWFXTJUlj4WAW0TBAFi9suxZ+v5uHSw0XHXTmYBQizL7piH4LUodpltCgj1iag
unOXYbfvObCJfftH1ev7XA8Qj6t3PSyB5thGgXXv+W5/U5a7HmpTRigqMVVT005MATjZnI5WT9go
pBii9m5d2F8xCuVJcyyP3aNI1iVf3OO6x866QF5fFJ4N6jw9I1GXYYIP3KasI2Wj8Ld+alFyPctu
aHFK6+sBKPQymkveGyEZDRHssu3TaS/Mj9yFU/dABEkPQ6zUlno2tLqT53YAnJhrWRfRuXdA+c7e
0ADQDtWjwXPA7xjJMA5gNbPKPKpXRl9XAzQINPWpntDqpFBTZMa/oLoasaI0504RatovJKan0eLA
hPOQ4MFfryBhazPeyvkgk5JgkcjAHdzn9XNmhi20vqu95b4JgfEB8ecjqPe27yiHcXDtXd/XQhG3
PFOpOCNb+mEFcXbvk7n/lpDMOgHTaiaxneU+fW7/y9IPrJLbyI/XUjVnUjZrCb1cSVDV9/3i/eGd
40hSG9Z2WrqUsXcuzJp0Jhc3j8EcwyUlfIei3ZCsuCyLVcTbQJ8rdLAfwF3BExl90XZJNOuCqrNQ
SyDmLYJyDhPwGxXmSbXjm+08xv3iGfV94VSlcV4u+UP9oDeEAHBFKovns1Yl/F/hT0liBDY0K5Zu
Jjj7HkhrDBCsPJ+2Nxvu4n0d4P0bnN6oFShBrcEgkvWdJNggpuw3CVagyzvaeFxGdYEEJjeUZYf9
a+nf5hbBpXAxiJiDVC8T4djH0Dk4TvJT/MGujBu+BNT9aDWYHwMfLPnPi2GojbxVfTkcSdI7yhhv
dpyE5gnztaJQhyGuaKILdCsXonKHn8cx0jfngDwIozdMhpm1xXToCvkT7rZM2+iSEFusEN6/J2FQ
znhammp9vvNgelUelUqVcSXLbSgLXJ9pBSczdM9R58depvQHaUH/h3gNpaDGP4vMaQxty6WzcNjp
qNEFt1OgdXnewgvtmHmegTFOcqwAo3LLi3o2eIkKyINoBWi3FqHnJ7L8FuTsAVCabIYIRtt4iDSr
eFR9PwzXdRoo0Sf619876IY1zqTrNIOJIOoTgajcNDRpJhFcozvzpts3wVfSih7nLJnIrfzep5O/
7Ep+UehwtTAJFFQQ7VNzwt0SbGvkKJ6mVXSVe7jHjK+j8iUC422knl1Sq0m7NC5JGAnOT7qDpeEu
2TeP0hLbJf/pRM/HGj89vWUTwnNYmM65BFCyOygqJlSZRbfaWrIPMOio15aUW9Rcajkur7EhPUs/
yFDxhbaqTWT3jT0/l6Q3ZTcqux1HCG8vtQpFVZ0jkHGedhUBh8x9ZDx1v7/KjIFaR8kAZNOksARM
f6+TUjuFXA4+ikZiflWO9ULBg0z+oK2+M6R7Rfn5id8Z4UZ7N4FAZORxAG32gJ868S07WVdylnkf
B8RtTkpe65GYj3PkGO6kEu0Li8T/9mgtPc2G8xMoJBd2gu0E60TwDc3dKW9PBq1hLClESabLGyd5
k/ajqBCs93QKs97T+aOv/9FPd1EcAJVWfjfJ/d/tCzx7R36p3HU1wdrgQ1YG9Y4y4ds1YpvvHNI2
f9mr3dpnnzE5l0uav6NxbMxD8aWMLTE818O7bNGhfbZVwMcgxE9aGvZwMVWW94EkgAlAPC4W96q+
f9axRuf9wWEUj75OXhjhSsvRx2h4dEf7ET9ZEBwi82JSgRxG/91I/dJynx80AXU+sBBaiTn5QWFL
EgILUfFNvUwreglwVkNtqglYs8euNuMe8ycXYNhVuCc248zKrmtSNhNgJn8mnsBEDmosjZxmKWzI
tz31gUOh4PjMW0keU4nx/AsuHnzYqIh2NZiXNYMozWvo9M1Kj/lOI+TyigUqYA33ofgTNBjKPrcM
q74YwoqiGOxvs5SMt05i4f/FWfu8O97oziyC2+JIOcaasBpcUXG2DdxRcTSoUC05f0siqvQ3t1Rj
7Kg5lJkYDsNJ3BDfuCp3b9fgkZMsBAHq6jQROdmE07fmjXIZLZxZmyZGU6dd/xt8Xdu1GTl0/HOj
eTr3R80YYIovOnkvVaGBRV9cQvNE5epB57wmdcUBjXV3rHDhZU9gEgd0H6tDM0yI5vQqLMjTid7v
iERL8RWQRXpoTFtbDDhTvzlR+4YG5oZuia/o92lPROlBJ1Wthx47xo3FF0R59qOhjccZObyEQeWo
tIMl9+jSYiKrcV4Xb4RZpWdCnGuwX3vl38jeDOUvSRKrLD3W9EmuSIvxbR0dQ4b4czIIGVpK2f6Z
9vsxH3o6lufOQ9UKdk71p2QONG388GD7ILFx3egfLNiWCl5oX3Hn6K0NUw67z3xEVrakISrFTro4
i5K5y0FSBJX9nZCkiGTApuffkW00TfUQ/hd4uV9eDPrk4I4u8iCFy6e1rLPZVrr61Sxondm0zCzy
8Dnry6UsHOnMLN6Gcd9sqUnUj9LRQxtBl9nNvBc52ygSUyCcvI6F1wo66fcFGCHY8qzu8wEZXpvx
nFSShEG4TWMKXl1TNHKPZ8DD5Wl1b26BzvKckxobnl45mImWqq+mRG3+s2BOzXhWORjp5iSK0ob5
JnViReFAr32SEQ22G3+rWvr3w+QHnL/Y5FPsGz+H+9fauImO5hnThUoviZjgg0ESi7JALIJ+2pq2
FFwc6fkImmNPSp81RmUbtIawL2MFSaVXPvOTjlW8tcvAk84N4i+1R0IP8RIBRH5KhH/v5bdz5DPh
oNdnHovZYSzsr+GieLoBUyIbsT+geooho3dfOe6I7oKQG0cHJP2hGmWZU9hpEtQd3FkrNFv0USti
Kts9dYlAW3x6d0vcNc2iZ1Z32+vwgVSm9iAuAA45o6imLFUC4rXCyjnWmt/agJbbutwYhdFAhM7H
lBYhNT8SteCDxvp1A6U5jjrkaAqYwsjxgG4kpEFbPy8HND/qpCJjsqN5UV3xklSNN/+iiMggYaSe
76Jnh7t9qgApx74Kk+XaPhrtCZs4mPR4muzye0Zz19AGyCeJluGdDXdzO0aA9JY8/f1NZVJSPL2P
G40chOK0dcJ06l3n7pPhWYZnhwHn6nrBa+my4ytXNU8j1Aqn9Nn+ogZLLxzHeZxZecZEeMgmTWTs
jIymDxBiP8udLLIDO2xtuy17DcbKCqIoDSr4yheTX6CpUEDPqQILuA32JrQ8w5WbkzC9r7Boh62k
ziAQQUxLzsV+sx9gQVbMVecfybxcSki5FeH47cTo4Fn4uiLqK3D8kGa3+A/sIp6pfPD3EGRxaYm/
71aPsB+qMB1hiHrdHau+tRHnhobIajI6pDOqYqUDiQZxDy0sDzqTb2syIb0X1uAda5GctOLAV4s2
mozldIVKz7Xd/QwiXWdr7q4qYKyaHFMCTZ9RLAOefXPYy7LMJ+c290CVGB29YB5XaNRUt0uuzg1v
QPKtJB5OkOAxdSLeg3SshBCMI6mhiDyRO3hh7WSD9ezFqcJwS2BM6uWVseeGTywbtMT9dgJUUqZ3
iXZvOqKcEsiRct0YX3riQMrmdgRhH6UIEkinuLmM7GSsReOjggS8zrTXSxiNnQDRSQMiq6w4MGrQ
jvX902pZliaMbmxfxyxd/ewlOC/i7FEMTzGo5I9JTSTSDnkgRWZbzg3xOkxFYMj0nVcZjixC/d29
j3ApZQ+kGFnP4K3KnwBXTy1Ie0MztG/lza6BoaB8bI8dFDih8dIF0hIQ3ufL4YNXfglBYSNR0eXE
sWAST71ruuFbW9IWVrK8iYATzI6MGRNKOHOJ6txr2f/GyaakfhqG5rNNEEaiBz9sUGv08Z/iwZrQ
6al3rwqDuk7gpt+DzWukCiY2hTiaV6vmZESN0Uz1Vpj9WaEfWKtWGXOl/a+rY+wmKJjYBxiSfduJ
bFR3NlUMjUkaPHEs3r0GQH27R3XwF5oY1pxsaUDY1t5d91hC5a2HgOu8FYNzvbu8Wp+Uj1c+6Ny0
Fut2/ojrdK06s4Gwc1RqOgdK++ZFbtdfkTqXPtcWmU3ox7mB8WTuZZV2tJWCxrtdpPFZM6gUcd6y
rOaJ6l5TUXEV1XRezp6pi2xA8hFWSvopJlTQmR5REv33s7D888C4HYcUFecQMyxgKSnhVOZxm0+b
Hfg4iXhF/iS8lZ5Us7W5iIRjc2VnbPBJbgNwcPgRlS6zOT7x4yzo3BN3fJu1cQUjF4RErp4JnXGk
cEKnLPd48m+soN9hE/ZfY+GO/GG8hWqbdxjQD4YHOuSwPsEflgBDKvlgujWNOCrgBIc5PJCmcJH9
AFb0NQqdcRyTVPfymySYiM4YTYh/qEMf5JLCZ+4KKZoPVE7kXLKeaiqmw4sl25GIXb5uRF9I19T7
LmbnfCQhF04rT7GPwKdps1tqi5NBryVp4bqn9RRzXqEA0VZVM0VhS8pbS3FAN6C88H6tqPcmIdpc
mRan0b0QfXuJEOebAW+M8H5PmP+G/hM7fi1J6O6FCEsJStYq72Du+B36GVp2Sx12TeVxH80BV3DD
qAEtt6r2YnJjI+iJDm5lXf/28hvCV8D7mVYWbQZRPW0nPY1fz/g28+ZjTzUKX7mSCRPJTK/vJdR4
pxKasPYZ5jm00jOdA8HMaomiDs3fLnEPqW1X0/KO3YNcK8kvsGVftileqe+o9hi6K9l06RavuQ5f
0R8KU2VmXH+vgClXojAZUrCzLssvlQ9YCHANxxjrmLsO2FimFfW+fIWte85hXHIOs3A6ndoHEQ1v
Z9+LLZw3SqXM9xtPw+kKvKB7OkhgFOQBSRqLhFxRix1Zw4CtjW2jaBs5H0r3DpBr1szm5X45ske7
5Bz4eABLAEtBvcHvJVY1jZEwIVkHEIlw1qWwD6Ir21mb7Dql/O+K/lXFz/ds1RaJyupMmZIEgJwf
dD1/E66G8a4ekdjH7q0N+Dl7hNK7uk/x/6Kh8i2t4fEInvDCJnf/MOdw0RcFc1kunFDvuCVXYlNC
KzuyJ4LLFwaqyNv0rarcpJBHRPaM0e4UsIZQG0uJKqaJ2dBysRbDSR0YGSR/xFeRO0WhUgzVCQOy
L6mIOS9IxqQomu0uXolzOhbOJ1krFEbnx33vMVRR5xv8EJJKHQZps6nS/OHezoqu/0aJYkJu9Z9R
AnZqYqK/IWS6rCXjeb3tzbzRaaHr7i2IDB1rzE9+LIEjbKEfpF23sD+XIk0bmThdprG8wZS88jB4
qpPHRYSTG+7MeqmIjPad8nRe9sGxVJS2iIiIKKDR0QX0yZ1+Bac52LYsdMjQXSPhBplGE/ZG5yV9
IV2FiKN8tf4At7f0o8eLltZ4VnLRhm5TPcb8ty5O32y78i5BE0pk7NoJqeCcKAhQGsi1VD5aObtZ
SnP2lyvlslLwxkxItn/csmYPYcc69SA8OUdeVIENL5X8tJH5R62ZfD0npz3juozCy2A2GTUwLrqP
CbtfK/R9CUMx4ca/O9V8MkgY12n5nNCOl7gldtqT5Wqn5ZaFHmm8abOkGCvN1NPrJ8gou71gByWI
SNL77IxUpR6D2RdSIgDjIUss/xpUOng6DlbTggyYHWqELkVvmBFZfmKnp9cDt/HexKSEvRXQ84fX
LTo+wy6iKeRsGASXdGHmWt5fOarElWR0Ob9tCC/pZxYsJ9ffISYJzZwB03jSywp+SQVtYoB5rZmv
+V75VUw7Q5Ckvvohbpset2y+r9YcLJ+fyZY94jX4TLIZyKaSU3Ab1B8PASBlb/KNrbtGIG0WrySz
nFwcYIghsUhwMSALK9b8mAXMa6Z8YA3GoLUTHnJmP1RsyxC2aEg7QyQlvI5Xn5Ep8k6zKQJpsktL
dKQHg64t4ZqgeyI3z+3rGb0hqzdqERfiYvSw3pO7hHrWjW6PxfG45jBLg8FDm4B0u4ZLkLTX+dk/
/WkkRCTcoZYZlSd69gxUtW+tuW0h3qxKrjD7wAeSTC5Kv9BWYcULmaWrirAU7pnL6RlpYnSm7WnO
kSdAeotuDuTykSMoZGCyr3YFBhj06erJB5/HIGAY2jzunCfr4Lbj2z12WLS342AxEc+IKlX1PF+s
5mWcHkYJhslQfZRMU36IIm8be3audRboLh9hFe0phbUcTibkEH+MoQlYBBPL9esG5zxGrBSdF5P+
58N0Un1hcYEqi6r2vbnmqGKRwP0r4QfTaatnsmxwUKNAi3BEHQX8loJmp7TkyhBoPATWXzeeImEZ
9z09HD93Ov/aLHBW/bN+dp9/Z18K9RvRaiPzEaAY1DXLf/cABLhV1AfBJuLZxUHpsn31nMNNjzpL
SN2pXlUlOZiAdPoZkQ2YzQ9p6JNTTKFUOJ/VsrAgtVRRW5dVrtGbiNmv7jTawcrFlFraa8mlHgB0
wuxeMRuV4SKFAibGaIdvjk1jNaIIPUyuPgtWc69ZHKra4zPYMDk8kCwKb18BFktU8Iyqik7qZDBY
l7ZctLWvpGWJkvN6X7T9xaZ5ifnSEi2oa3QuH4HIhaVusZ4RpFaKIsnt7iWmK5WARPdOIpdy7X/S
wtBqqVq1IgCJVa+ybUvDkbe5YIyb4AQR081xbcc4Btdb2o0e+deFTdAQn4KsvNxdkieeif92DKNk
HIzMfBkf0gloTYjhH2WXNc/6oLc3A2CKghkWj5PlgqJXZiav8Ro3M8Qzdj3eFiiyzwRENvIJNGQA
zHNNGkbL8QXtJGC/wbgk7JRK2Ru92WP27r9ET5TGFboB78ACPvJ7QtayKXYQWkY8TRMQxrODGZbp
fizGhvZlSBd4yU/3l0LWgjOmq2zEx313xUlN5GExhEIcdr0D8hQPYhZaZOsy1HOm6DJscaX4N2ki
WozR1BoxrRBbwymdoQky5j0jqAIJ/TE3aFVTX0123dUEqNgyXSMnMai3dm/TcnSC8yr8ll9FmhU5
qNyfO8LcucYid+a7XYNlfJkEpGFzfYe/2qF0243GQS3YGaYQyAP9AvQ24+TEXt+m3I98H4fB91sR
phwDpVFNLeVZssJfFNO2d+1ImjhAA3IkE0KZIM+I7gvwspqfSLK9YGwb4tTJswNofDx9oc88LJ30
w5XSyvqDHLMGrosSWYJ51PeJLu2EA7y7mwf/Jw/rw7ooDkV4lCEg35SxCaFGdMtQhisgJNEBTSAp
l0ccmhdxAYCyUTvP9Y+34vYRjQaFRlHjxK0LX/E/trZ51beIQEUMgwypzf5dIs7eP5JFBVpGTMRC
tHd3UTn4LT80mdD+b6GsOcAFOECNZvPjfdjEFfD8r1n/UlzTvAnaLbnI/tj2Xpay2FDRPl9XXaMq
VjTd11x3GoOrGmbGtzUXCe45Ty0+NXvwmrAempRQMnGxwHsj4CKn4qa+1H17cU1UWE/B5HD12Mh0
gZ+Z834MDX521jFKGybsT1IRtJlxoytTYrrEBpVrdXuw03T02SCbS9kN8TiZizspwMZISHZ4s33e
L4hktIyVv8idMMN/qznBayw9XIBxEdya5uzCtOdgzdv8kVeQE4WulxxVQcR1lYX85dijY4NILrzk
AxX5QQ/8wCN8NNcD1r8Vf9ZF/u3ykwSLqGxylUfdby/Z3j2/jy+/6E0J04KaEz3EQwRKdIHrieru
3UPQoZZoFvTPqNIQjXkrxKkgTqkJ/u6AccY/IGaViU+YsNbBluEpQu0EK0W4prY7uKi9ymwj68EP
vR0AQ6dy9dxZWI6iVoWCS1v82kSXPOSEPWYxP9oVuA3MbKOfORbO7QGP4laKNUQcCG2FTZwjJmaU
BRpGapuUi33ewFx3QM1U+ZF+tcvQDOzLGgWya8M+fG9BKPMDm3IISugEVY5r18thMiWZ7/yVRP5N
ZufBT+mSzxoHQKfia2+G4Rk4nmTMKR8ie8lecP1tgkI2CklbvwoIdr6HS88lHE+Wj7/yQSbOgQL7
HUAU9jc4nELMLsqXXGFQBiV02F2hgGMRsBjH2TlNzoJqGUHUOT/8UISg/3dcF32n4RmOi+3UZSBg
/l2QsuvImC7KsEnh3IEYMpfOi1tlNmnX/3WJufZQGZGs0ksP1Zqv2MoHcBv3DjIn8R2QkrNjEADA
WB0ft5w+nNMOvEgP/0/TF+tXZOK1gS4Ti2MkUuiLluvqit6SBmOYp3GOINzIgA89kMDn/PWEnX1y
kB7F/CYt9DTahbUGbIgBckvPYYp8u2TTXjj5AY2k0oPHI+S7StbnZjy39o5cuozvt0J4K/+lyq48
l9O0N+TY3zuRuPxsUTLqJKfh6ZtHB9MqP9DkiL4pP49gb7jxytdGCInXTqvm2JUX+1bQ57iNt41f
CEj6gzS4btlxZsrymD6qTlqS7WeOECBZXde3CwSzA1GvXJ8MP+1UG9+IZYl9f6WG3kBRwtbCy2DT
lppSD5CWa4wIW3fTs+5QUN7TLb0b29VT2w2dFs9QNxBUz3QF24LhwlX+LKwYoqBdR3U3SiuUIu7K
cBj8wIzvfjiWeejQ6xkp3fPO0wXQFeJztI3+h0KtOR7Z9yRB7bM5w0lDHDOtXBSgqQ07fAiIJ/FH
7MoNl0psQVgbLVMvwYxr5IcNQ7iyerFTak5FolbVBXiCjP+aZ02Ezzze3SvJxuoPwkuC2MOqKk+V
s7wjsh4QYLiJEp2HxWLj1ajNt4VCjE1g0WoTyCmesACKcTBctgwV609nxW32EBWszVkRgiWHjQZI
ogtawnOgCOUtduJIWFpcbAFPW+u92/6qKadXvSHvmSOIfzg/ayPM7/Too9SyJp+7p3lcbT8Ylq4M
YRlBqLBX+KuAoNZi1iWHsZiOLLV0uoeSZB9Qdh7AFDRSLmR7JEzeaIbOfjJYAHlgcd8VX0L9tIyg
HbejjveVujPhVpi8pLBGroi6PFKN26jrevN/GdhWbNkjfBeehIXSL49q9ff0weSwKW03lnsltyi4
ooNVNlgwV3ewVKgOZm78WHx+b+WelLCQnzx17OCyW2hbLgj3PPxPpNe1DghgjT0MXmV2f4pPixcg
pt+P/tGw/rpGVV5wtogaT/qYz51MnTEsQFWHExemwYmRY7AFmZ/Pnlz3CfuT5g+o5bhti/vP0Exu
w2LJPQJH2b1vX2u2qixJY0cuitEz+mjPw+rKZH8QkN+mpynLEwmGeqQvcACYV5H0Q4oInhcEBTCz
yja0sStiYQ9DT500jywjHFdLWYdkiDDgkBq47KFhh70byoDubP/z3WguOXn5wXjSLi/WEuUlpy7i
oTjR8spUyuDp2wqcRHpXg74R3J9yH7bvSnhUocHUxB4lYJT4IToG1LJYUkf1t7Sj3MqKUO9jlVm4
pViL9xoqcgPKJ7xXB+NIXqbAaLAqbmeqMjxEjPX0wQZdm4BqFUJ7/7GdTvycmvKRjbGYnIbRivoi
P5JfKEIxmIvLQ6BPKdVK9bzh5YiRrpweXXvhAiDfCHKEwyNvzfvuJm/XrwEFMpcN6zNgUTc20eNt
6f8TLxSX4Di9MlhX6Bw01rddIrNxWWrFRD1dEPZZ4BE7X2qOjkxOFIqCb+/jpH8v6BeznEav/GyL
AB6Q1UwkvwKr/yWsTxk3J06uAKTGF+zyjBVIWVHrUaingRX56aIAr4j5tLSuHmQ1O8IviW14g/Jd
kUot2bsPqS10ciAdFE9qY0mcoh61CoYTFL17xKxATrponMS3io/XscmG5rkIIeChMkvewZXP3wMK
Cseciy0UY9vm/6anCCa1miu8aHAqREXPNcdXQIp2mB1P9bcE4MUvGQI2MuVFJxnZoMqWZrki3igT
AWUfKTp/7DpizF/YPXoEwv4H5XBRRtmbo4svDR/Ph0ZkPJA0SpS0dW1xHtukknx9OiGF+iyRoz+R
PQ+dhT2dSaLuFjRgu84HdvTrDguhjiYQclWLMQo9eHSm8XN0BBg+27vIHQ8NY6APS76iTsF47VGN
sQZq1/CFNBbr028ItVYfiUI0o8i1mkXTvYv7PVzUWwWvxNZTjmliGFBV9x+7hDpXcOW3aAHwf7DT
Oio99M3jGFqIRWdRjIoR4VG2FNIemoN+aHQdVaekgJckmbpqm5rSMk6RoVeygRbplAxR4clTh1sr
g99+lssiUhhMtEUu86/q+afEEzdcV03eJ6d62OcE4Wd5GexDQghuZaTbGBKYpscxRLhD7xwSorQA
Fd2NcKFgXiG0BTZ4OQZ5yAbQRo70KM7MvYD1jKwwQhT1Xa58fWmPKqpkbzUcQx6KXTECp4m1YPZw
mTqoOQDQEF+qdV6H/yEIPdTxCxoXILAD2rWzH5RSmStC/+P1rdo/dlk9oT9Qgib0whWFYc7gLG6f
kvMkdQP9mC4rTSC5v2zYkWCODJd3XJBqYgMB7dMwB1ATi7n/xS8Q68ujNn/Q3PGiapjnleP02PaI
B8rTsXQfY+6yWVPCCXoemAme/jsXiwhnZzp+oF9jEVlIyB9IZekqaL+eg4bHnERWYU/Q9MbP2KdP
wPFdAaIQvMetpclLiQ92U3PM9solrAko1fAg4Kkn0ieoXNFzqjUdWjDTchaH1CSQWItfelg3BKXT
qjRvLhmQSrHbMgDiuxn7b/8CYdNVwxH24T1vqT6DItakb6GGfuLvyHLfpRr3CAmvHUkKcvlWBqhb
nR4chyb6Ha3qEMv34sOd8dT/sGk72CG7Oh7Swc/P4/WEkI4aMDGXRbDdOq40hANM+sJjYXcDjHKV
VLWWp8EerQPBA2mVm8e96HbliuUQDQK0ix8mTdnw02J8FO0sNNM9sCnvUftfYm7uvnHjGPZM+HeP
BqiwVobj39PyJrdTXwfssw1OBQgnjiAggB+uJs1Wid3erRpF1BxTky990azQBob6VYaSik4O8M95
U+2EFHF6/3vm5PyO031HJwzHgoEbo0tqcyTsHRYHxM0xe+247md4ivkL++i1Sp6bS3DtrOoPdXN3
AASa5G6QBVWdJETTjmcfP83tFqbApSmOaZnDnOEveCnnK8UdTeMLE36WanPxXoQs5/ACrJaAL9hp
1M+cyUn3YnVlBOzYgGCXb5lD/lTdeA+3Hb6mD/+gmF/Vzah3nKTT4NaU58NH4S6d45wrkIkLAmTy
MqkGd01G6qEiIDnY9a8pWL4VJXSe1gpZKGYfPJyUo9t/wI1DGdXijRWXOOQJyZFuKiB5NavHqEs2
l2RNnKn//DOOXTzcHSY4H0U+y8ycae3TGBC9a4RN0E2Vkd/De72a2s+Oo9VF7DW14rSutEwaFfgu
T56JNLXKJN8OnYEX11Wok9tPYmclKRtUU2YHnMVo3XmR2GUxA2qqNVGoP1Hgbf3shqLVOgrp0JvI
n+s4kZzzde5+qDKrs0EROA9zKXAsJ/4UmEiTt1yaqOyoECCYKyk09BIhDi/6Aew0iACDnq0EGha6
qCPLKTBRI2DX7gAqqh2EamEg3jR3dJbHii0nQa25J0z9eJf6ZVAGmaqUsfw96/2v9WXw5mDVKLB8
PvsXKGv6cVrCBmO/60hTcbNJ/eZPkzNofcvjJ5P/rQC9ZxjJtLpaVmLorRTi1XjiJZEVeZ2W/b2U
2kGmu66QB0pINnmXu/pwc7J5UIxyy9E3zBGrnhEeGYVnUcuJZguyig758lrtIkJaj5OHaMVAHNZY
pBmbiQK/EWAVX0e9U2as3MCBLWPZ7ARtODJMPUJtlJ678JuZ+DDr6Fo2Ovy73ojFy9K4jC1nFe4m
N/GcHWNHEmDmChd0hRs4JDmo0ukZTRiRhGD7Y67bDFTVfeoZ6R8UWKFCrIyVwSR5UO5lbxLLJDgC
LO5G52yCrBfEP8gRMs4mmOF/xKvWWcIGDRxVoC2nGYK6gWZqkSmiURXLADEU3fanVAqSk3jmLHTL
C9DMekWBjAmUMqDBPtLs/twPJeFkqaQJp0HxyNuis2dXJCbsnjZYOMtybAEdlPjNLqXChnSuHnrb
16fdI0xTZTj5WHOu871OQFfpQmDNatZd31zwxHQzE3cJp+lp4sjs+qHUKThbRsnwQbDoNrv4Yt7M
wldyEf84inzhZQSKDO+Ffu95hjInv+u4BcbMHsaoh2V42ej+tBXpd0C2ZNPvHLN8XvdjrZS/iVTi
KkS2ems4hbQCwUAdFGHNfzPb8zSc65LzZH30tUH7eCtX70KkfQekPwukVeMile9QUux+GHJWRp1k
kAS9vEOCTZn1fEmbHrP/A8WoKc0vv+RxO0zuBkp4IoLDNlkSAG108aw9JznqNxpCc2qii0AAlcI/
Ohjq1ogE7nmc74UegSE3t6lr4xh42YOM/P7obR7EdeYmBs8kNZl9+SbbrSUFoJoMJPIRszNo6NOX
2nhbYb7b5PKblIwrj5EQsc7lYHkUe6T5rHDHDWzebLjCqqETMt+0IiG+ekssTxiK2NCwI1lLviDQ
XUW4IcOYIYlBxle+tRp961XctZAkKsqYku9Ywu60h2N6EFtACOAG8a3aqZEZnaJEWL0kLOa31LuM
IhlQl9+UE8UWuVXHjwjE81Suo8vnU9mYvglQywYWuiGyIhJBmHhwj67jGFhveG850gb0/CVekjTF
DeRnaL2oeJYgD5+9kdE0997GPGMwIG1fTQGyRIhZ24F6CqkgaC2tQZ4kr1ELswxvnajcdDVu22sf
1gK8ZOPphI1sbfq7HrtZLsVOA9/PRJx2tGFfEbwlqN5ycGr5wbgw63QWEEUga7zTcfrfLNkhS9oJ
Ma6pw3k8eTJnoBre8l4bndhq73EiXmDU+qA6rCLwTHOPCtmkuMGF/KYXckrbsDY2nvX1F/DJVV/u
qt2eGUuFvQ+JderFHYBQWEiFwGYdbIE5ZT7I73pkkK13ME9t4dt0fCrHsKmhs/jp7FyC+JuUGAZG
OHOlXDRZ/RN95ewCUiveM0+jM6d5TaZiCH9tVH7TbPNXxavgPFqK4yQegcFo5Zo7v1xmbkvSh7WX
2CuqLfm7Z+16/ov1rFYED1i4gaTMyjherwp7U/5vzXu/2CYh2oD0mJf4oVfNtN91JegdSR2tDRNc
AhmwbwQWkyynlZX0TlExbkrYi2k/UQiqXnaTbJMX5u/ijSsbt7Yfvn0lGLWK85R+EtYVXh7fkQX8
WDwLsRqLWCfKqYJf3dcgkDoThVnlW0YZG55lWdnwNUDZKMZDrMEzZVWtS07HNipraycBFJPng6Yy
oeLT3ofD8Gm3IIEHeBukoH3PAgsd6jjQ4/Wrmw6eDvktnfiAXvEyt+Xf7ehWDKVXVZ+0VLD78Ro/
9aJtSWzxsUZyF5Wgd6UV1Rkx7okdF1Tf1gcLicuFuVpedIw0zODrp5VfXp1lwcSv+EuZRE1stQ0L
HDB5rstJ1Ch7zMcvUqMEVwqnAl8cdYdeMqFyi/aV+RbYUmBr/6oKJa5f+rUFbZGLyq7Ojx5S3Qce
Ves9LRGEUR/T+xbiQFX+J9lgdM3KU14fPU3MOFsFjiBhUf36Hcj+9r/Rvxn+QhdgNWsNfODRMVAM
e3T1Yy5PKOTpxcoeGWsv/XfcesfwEHxfVCC1q0hjfP56FXFW2drIvFlft9k7tdnD+RTUtlq0gxnr
DhsHvksIxtCY+IwX1oGtgxHMnKoOFGNkM5FzNQLGzin9FO8upP8vL6zjdtGtTUv4u13BZBKbh8cA
DowaH/ITUNCWNmndlDa48teyO6/yiMdKWd9QDFrdpJ21v8jVO3WXOb5nUYd+ow0Fm7oGCRPMbYbt
w6qtA9Z6aqdbtera9RWv8kGEqX70beiiTUzOzFWt14KD3DTHaS1KakAXGuFck4akMRyHC36FAGlm
HpjnvjdogLxv7KMUXEyk0Pfhr5zh7dyPQKVPJXyxPufKDdYBZHv4efsEUEh9m7P/LXwOJAPn/rQ+
kixyXjRhdogvAEJ3+6yirV5RQbvi5qkXFiI1ipGt6aeXL/jMk7G9ZRgf8oAbt1+j51qqbYWqNuzZ
hx00lHZOa0acKMtsgWlPbeChHKLpsK/ri4AiE83YmLPpjxMANklCqXAfg1HTCJHAxP+JoTo1Ecth
4bSzyxEUo8v+lAp8iJYBQnKqGyz9PfmjVda9TBGMLGqDpRyEOgalhXwMyzKhUHluOq5K8zFDPsRx
21XFAC9VXwuHlIw6200hruP42rgI1nQQu0HYPlgtXGZU40hylooSB1yhDLcZP2l02kaD2CGJqhN9
y6444jewp8zL7llm7Q6Q8U9g8JZtzVtYIO09pUXTs7mHlEsr35iTaY2DWldb4FLYSDcUL9BuSo/o
eyeAW+C6qVk8ClhFpGe/JAfWwYYW0eMmbGsjISgSoPcxh7pn3GGfVU0TWiv8WY7TYFPdoobho2c/
GixUA0ho0nVlf54nDGdKzFWEY/yw7+Wzvqgl/j2WE0O09k3f2mMUZyS8XJRDnN8CdGxM5b8F2Gju
zsnAdOMxNm3VP3+/HbIwvekKLMQjIYcgViMjms2EVTeiCJE14ke9s/Q6tL/h3lvkk1RdPzS+rqKe
IeoknT9KtoVs21XR9681bqz1Fki1kEzOZJ8I/mYhXdBpKWK9CBpXwuKBCqgPUowF9zh/IV4OLQey
s5MUYwyHqD6TyVf6hYLj5TZ/kxoxZUT9A9iYq9vVFy5BqU0/li6ufTIOxk25NOBgijo7lGf3Ecez
iU1Pttlm5nRu32fVoafVHHNbLlxWILGODfzRLkRe2PbtBOO5hrINQA6BjYcu7g/e/eLFQ3Fh6DIx
Kptc9iDx7ue7Pe2qt+aq8c7MWLh2bfXIAU6nRg/VQBK/pxadocq4JpVfQ/h9BAuFdSreSsH+hdf6
qmp4y2TLXMCoRZSW1nsKALjs++LaCKYklGDAMy0h0afymbHglJabJ5N+iwR7hjT8XpDrejdAJWv+
ZkFEbCmQF957A+A6O1Y0Qqjg7Ngt1fcZ5wXPgD6jNr2JEexip4g4+v8sPN8NzPZ7R0f8+gxvBF+2
kD1rC2Jn2vgf3JVLhHByhr8uPaU+qDWOnrNqVjV6Ax++et4/58uo8S+8CtdZBvMWffs3YjB3ta4Z
wykzusf7jxyXDsEsvsoNgGR8LoGF27axSJrkzPr8j6zewZvJVmiSVQ0UpPe7ZoqaT53C7hK7Sxgj
MJtyK1sQ2MeCgz9s9x/ty9JDGieJSOL3/gSS9i4AJyexjwWMsKYqzQuVC/BH98epeZV3mVZy4WNv
oG0kRgOEpfk/GNWvu95rTBYmhRk+WZCDdi2tSDEkjR2k13Ep9UyibF6F6Oj+Kf0gdXq86yW7mq8/
YAppM9XbIXbIZaZc7qggvgDf3bm2168gLvHxIFnvUsqetUCY2vv0hQDjG370KF4SaNwDWanfgZVC
EzVKI1uU3unthHEappLUyDxWKnYRPeSXaWbnVH1oAOQdh5HwAvShw2ae1FP0cgg6otmbgDlAJZAB
QGqstfC4t/S9xZBg0g9WLF0wYj4n1UqS/K3gx6iTixQXTmh4tCQEKvjbixpa0I2MxelHRskXp1ZL
d1cuiELVE5tR6+YJRAVdj9h0bogh5e/67YCLY/nZ5vcXPSj+kkfHz5HRGRkoT43+iBLVfSvsljxh
++uuKXiyDGQ3zq3WhcO+cSX5QbGw2CyN2ePL1RvJ/PnCVjRS99garX6JufKweVJgv3zeuZ6GslZI
VVOJ4gXFq6/x8JJGqdMkBzHjEaogKytoWz7rUqrsn0o1WC8iKy7vej58BT0IMKVBEUbxqrsjFHbo
Is90xEwyVRrl3W/nwgB/Y2FawR7OGyWYyJKgAAj+AilB9uCbLymRLQXP+gx+GWGFQYUTkMCSyoP4
S9JUvqGsLyWxUeH8kfw6bOR9HCO31+/a7FXPvjlRwNX2owLiLRC/1FqP4gCKuY3OHkbQgwC7pbX4
J40DmcA6qgDn/cS4tIIK0SV9JG2X6plQXS9lbuhyFsP7KC6Dz6VcIHz2uXhEPJCvYThvZ2LEZ9RZ
daX/BP3GRj5CR8ifc/r19IzDTox6mCP29kCD0PVqKGk2lLX3nBwdOSxkUUjQsYPXtjqvIS+5SgNx
rTVlBX9C5c3b13IxpucgR1N44zulE40Q7e+ObGqr0HwD3sqTDJb22nZfypcr3FTQN+uxPyj/aEML
1cDCVvUgk9vQ1BF3NphjdtreZYVv3tvcFTNuCGMlh0pyDhuS0K+g3ahABGJRZ0SVX59/x/AZK5w7
eCntigJnBFXVZIqf1lGolWs+X6rFsztdRdc0F9OB20SfBuEHCrf7x1i1yehnfKni6Z0bWrFW+aSE
LAFZ0DHZ6WWUsYlLt3Gk7dzb1SCKHhGwZY07EYA5Ii1j/DJPYQxmqHpBDjmXwtTxklCP1EMOlEpE
S55BtMcroQn58BLQr6l44fh+sc/8hagI6xPEKMaD0AZicMBezhVoyfOyTO/TsBVPOqj7btHxIvuB
nD4JwmVdGjx7Z3cRR6liGKJ4FKXAQklyF+EX9NiwuGcLfERq5AcE0badM9AUH0QyP3FEW9zl4GW3
V3QuktxjUsaNFkMMW5BrabgUeEeP3RwXS7Tb2u2ZfLc+4kcV7u85UTYatNhu1+T8GxBLj/vj/FRU
gMmsxQJXBk4tLtvyCwahM1Wtv2ntAjQRSh1HvXAXeJbmzONjWYBI3OwWTRfTd31Y0m8r/MfXxLt8
mzUi3w23MNXOk8TjyiWmRSxifkODKrAoDuTDezT2aH/DRD4MZpzFFd7hcR5EIM2SrsGDcuVowDjr
0G+SQOvKbIzS4uhKgwoc/FiZThRKu8gFR2w6e2esqXXvcvkdbdg2pDhZx20Jf9HQ4WOjqJpDRLpy
w9hVeSge2lkoeXHOFrQtKCe2ZSbALlHM5HR8aor03WaQchFbRaWP0E9BMxD8XqimTfu5e2wj+sjY
aVYDs7pzGaSvWs8Zr0g1MAoTTA2Y7HEmkKdM2yGIPAgQT/Bvo2PjmLuHXZoSqhgHYqqt03qcaIBS
ArqwqB5DHNSyC/OfasPBchrIG8BlHQjgv0r9bOp1emsBSqc3RkKNo3tgIBAIhDAKUw8l4gJwpmAj
ijI1WSfeizwaJCR/Nw8vCv71HJInWXnMk24nkQkOliMnaqHpBKCinVH/x89yNM5a3muLG0xk3WRw
b/R1D9layWIKynYd/owY/bd9xkXqKem9Du7RYeumUake71W0lDid0yZZBUcSz45xUuMA6ol7q+yj
FAP5kS3IJrr3oYvVB7U+kMdShZVhwT+7MeCIOofV3JlTtnanRLGUPwSLkblCPbfiC6ckDjZzHZNs
zYwJ5A3AnKqBsy0OYaX2BqxXBBz4yhisXNzvZGOSKDPZ8HSSYBWdWXOM1PAZWK6SvDAYaGlqJD/D
D7BiqiJa3yDXjApUNy72H3ELY0LxeYkCsehAe1MS8EvjvcO4sqMxFykaYETVQbXSidZVvl3WRGRz
p2maIK4DZqjwNgtT3kmDIuJ7sFtMExiQemay7f0hJNV/4TJLHR7FE13ix59tCJHvl0jVgHuSRySa
wafbjDt6yN5jADwGiEXeRD32sourzj8u3vVFDktwlSG1PHunpYxrWQZxXg96q9agHnYiZyLAER1U
stwsXlCJFudBmSKwveisZZ4n+E352pOKqg9SWYbnO0RFc76uYmouS/1Zrjdqq9Dd8lH6TlE+O/kk
FvnMwVIKyBa3zc0ErQ11TSQa2+HQiYF8ujtv7Ew+dFpnsZ9wJeeEt2dkyq+d5p4W2haTLoCRrZhi
epPSYwkI0r4rwAYjOO1bk2RmzjN1FPGqA7YvGq3r9/sKuggl58uAD54ICUAeUPnKmiqRSuxXe6Fv
YbpcRhDFZgcmy/hQHnouXJ5SE05zjS4DhKkH9G1yeJ7trs37lmBcfBLdSOzaYdexOYilQ41k066X
RrWg5Kwrn2AZzpM7jlJ89tXUNa57ehEcQnItVlRWYnmaq5SlAdS3FXyaf+XN+Mul5fe1dDvxtObq
xQZe7ZGWJW5tie5J02XWnYeuKmFdHPqp0S4XWexirGn7l93uTIF+qTtbHKbAvEhEp7jVI9Qs9Xzo
XfyYA7CzlNflhEkiEW3lZRg8bQniYXmzpfLnZWAihCjTPF2k9ksXhP2dKzDkdWGEx9/kby1f1XcU
IAvIxU9NykIPXHG1YRPecBLyix7SDVWc8B4+jutmnjOvJKo/yJ+KvwuG8VAm251GM65QkRmuCTA9
gqdF3uBJOXq3bJylhXq9zRolyzfW1OvgNazfJ8vfdUK6vHeoTBqN0oQhyxmSdhwYQePH5lwcM20o
X8twAOP+vhGFJOvz5fM7So/s4O9hZwAwlwI6j1XFF8NJuzRUS2pfu8jL/mtcMiNpd/jgfHu7qJ/g
ESrAqiK1MQxbPns3efkT/dzhDPyvZmmGNBFUILTqVofOTKIh6Q2dHNyTr40d5ObvqUnR1feedKWG
6hSrE9JxjYXtUtkMWNKHJjzH+KWRCXQRIP3pXcaEak4afCpg1hbI7adlvk+Dc8hf+m1Ym2TBRbc8
YEHNjVTEIVxJg3WCbt1m4VZx471u2x67gJCb52NUg39qoA5DvLw2mevJoHYLpDEu9L3xtYBuxtFE
8MLpDObdDAqTDl2arCR27UzxkkBjv7mjZ2vhg0JOFb5kfiUJ4L+YHnPWPlPw4qWVXfUoO+2Kl7Va
ABnuz2UA+Vh+tQlhFN+aljgelV2V9SZSx1teIGU42YQUKw2no+OT9ZqPxvGu7oRg7vO/K+HIn7pE
8KJhX/JCp2T5qdaWnm/zrKEqqa18FI4GupXuuDw1Cn9ZWV6WHZa8+5BWdIq44kJlsmQ7CHdDKxSm
BzT7N65C9c1UWx/BWwvJoXge59vUFtbtnFFHPZ5n8tiOiE9w9S+rYfUtjChILCVpnQQLO/gPlgsO
odJDy456/bk7pQDBACBs70XCIhsJyrDzvd0uV4ZlR5UewczemnnceAnlbvjvgDSz/EXfjwZaFdbS
JZ3mrvSR1mwCj7L4cAMXt/2PJoufstmeuefxAy/Xb0tJBVXvtogQOGRVmLwrq5G5ktFqlBSLHMA7
53zAKDH0bKq/ekIaTsruYaDgAcsCvIpHsdkes14WI3+RcJnSHflIFulRg+gBbhW/coX3GJMeS3Av
pHhc87TXniyZ8KKkMoIW8dDA9lQtqJiGZpSdxCEsDEFwzRkRv6JpRNhxXotbhMhVShcXJEPiRW3W
RlerKtaxoiurd313iOWj9hXOUeSV/guHuZ9ivv44Mo4NlI+3DM2TnPgMmgj1o/4D6nhhWrSSsf+5
hLgVYr3y99/ak0cezsDhvx0XULzkQtrAamo7Zx6OLswOFcSnO8TKTPHqFWT/jPTPIiKQCnpHWJtK
EsD7vqubF2ugF0ylQzddoAHYoXRT4QMcFoRwFPFbjE9MK1RrwzB4RaULcW92nUqUAmN3RaVJzdQw
1OYsWV1hdtVlPRThWi4te8Vu7lX9qkcrlX1ufXRYr4xfh6OZdaWZzpWgrNn1h2MyWkD1Z0UQUEOl
0+6K6kbeYIK4hZI943WcoBJE701GQZECQvudVbi7xdT0Yt8LSnPnbX5XN2HKDuwUFw4iW5alh8G3
zIN3b9AoACeydy+vvyE/IwM0vmRzh7r6VanHAA5pNs7Bdy9dyjNuYNqP7v7CGKO8m2lGdLgKcBI1
8afdyRlv4dT+/v5InCpWhSQ6bRGAZi8RTemn3uL8roTRMrgWV3Ub+eNDOUkQlZCks7F86+0kLa1j
F80vOxVCAfySd8ocLJr6keL4FKqp+YgTtDdJzJSnjoAKiVVcGIDvWpzUcLChMSpifKAL3zfTsUKl
rKeusYb2Z88GWoOtwFHuFB5C5vcz8nGF+LeK8yJFY0Gp2/quG4VWjBQ5Canz4ceV57eBQM86Syr6
Ptn0PvNT5UATHGLJz4DkeaGEPIzvSb4luWuFfBy0XKmw+i+XpW/oz2PvGXO7Jn7vhtdojDOBlMfl
hilcVJqglDJAHbx6k02RQ0I5S/2KX9aIYEkhJekh3x4imnaVWFkYdRGksoELoT6G77w/HrhoDrKo
QVkWuOyuJd6qbvudxDGaatmenA8jmgd3tThrmsqjkuaE/wLDIs6kLXatHjMzPcxWs35OvOOX/D6U
3dClYP+gbYFNNtRfh8Afepx3mrLL+cvFfKD5zfArWt4QNZUb9uSyBnGHyprh7Htd7ubzxbwG/N3r
M2EVD7SrWu4VcYQv3HxyGsgHTDK8gkHaunfyFfOBpXy8K7l8/JKO01s72ctK5vBfDlb56qjsntzs
SJKWvh7wz/z0aJU7Mw2wyiNFR2doR4/drLLNQWi+JMMYCVoeZXId0H0V+Ym96GzzWnXMEfbHb6Tf
wpLsC4CXpDCKPfrRZUguj+pt+TxpXEKsWTjfdTeFTsNm7BuYB21WbuzwrnjtVHBGYS2nrFQ6e6g1
cVujh7n7ho1r4BqKQJHPkbPiYvp5g0dP0SAgKO767Chi8qEkggoXPfhLiJAyBagO6y42ftFxThlq
WHSLDvIWz2OsC43n9eY40ye9S9LWArmjnGxZNqgHUZf26SzCJ6EpyEIj8euh5/57/ksVWoDPMgZR
gHOfqbJQy7sjXnfekDodwkYmk0YTqt8FKlZjFr4Y/Dw2Luknxmzob0GYRIrUWCwjVFWfdtQzERcD
mP9W3GtByPPTdN0eSDjjibJ1kSAZYEU4NKFwZNQbKhher+nYtKlJSA4hoow2/XmP/OAqZGDVIHYz
1vqLqVu9CGAo2pBuYb7343WlVUYS/X+/2q9RyAhOwLmWX+iOuDmPF6gsxxWsERKi/Vo80gwlUPKv
BKyBTfo9hoqa0yi+TEsr4AtonpGx1W16KqpNdCS4k1u+/vYc9ryJavri1/Nc8XVnW506MoG5tuYe
DqcY1kgo2Bpnh/PifZkoPqArSXiXrQBahXkZcIRwYtT4MnFMtEHkT/6IddohERFDshv+nFnyNFMu
RrDnudtTyNxQe7JAlFORdL5FAeu33Ghfc4nwBR3LFdQCqNW/Mbqwgv6hEsioBTaw/2SYJ+vQ+gnP
gfbT82FWsbKEkGOrlUcTITtEhf32OF4YnXReXmTy5O+o082tbYcLpdY8sjmZfZPSPqQ35dfjCS8+
LrzB5WVFOAuEITD6gg2qB0XDvt4b89IuAfiiRcG+HhZVGO4Pvv1ajJ9OrY+cG0E8Ob4NQ/hfDdru
JpWAL+y+kX4zaMpe7PoCah3DC8X+Q5JWi0Hq5ICOpZOZK5pbtzLwbbCl1sPhzXsoUiiXdQuWp+Bj
a/8kwLPSO5HYSEyKS4vWjlHphZS4pLqWySXHaHtQwxb0ymZnJU4wvJSTOEoWLQx1trKRYoNPSH65
VXxaev+Jupbwk4wUqUuxTPsBoFeaYzvcYOn08CKaRCXhgeAMxQ+azoxgucqQMzXUjnHPzuCcErop
Dmy1aksy2ehLuJwXKAhjOWJvJDNvOeX31h4mXPnQmnswoHRni3Azsqt8ugzz05NgIgbtMoI4tBxm
rGLm4DE0Hgbrd4L4rSN97c20OG7fDVFf3zEuRxNVdlmUgNfVfXE2TILn4w0HqCo1S0OcMftCxQQ1
nNlMex1mlkU2ccJdwC+eqU95BaC4o7Pz6X9ignpWjRC+CmRIMoqDwJsccC5Jm6RavIRNcHhhTOTq
eGKfeJG7C2pQSZcnGjWDVmSd33S5R3++lJbZU4414w2Pgn6J2mddInYmSGBNprm3IXnDYCimSgXq
oUG1P3kqNghmzwVVBdDKILxauYYSuneyovZjI5UhQ3AQ4DTYKcMTJosDKOFmmHDFc/lYKWdcKp9D
i87i8z9srBjmUmHinhwI5T4LZ8Yi4aQ4ErGFZu5RLQuSebBproeHGZ/Ki7nbfaCwTZf4t7SLsf00
TnJRCAAt9Hpydz8P0tykhgEvCd+YeBQI3+rjFHTWuLdT76Q8KQf8oiaGQc4XCzwbYIKDeUyjPhUx
iwWnJWwHEMR51zpmO4japlOy2eC8bD0y4s66wwyxF3NSBxsse+CKb3oEMbFpSr4srI0ggV01kYFM
pXcDZdiLE3TVeGpFykZB23BnfcHwn4KmBJcfJkrYZF4x6Yd10R9IM+ui+bQ4C631tIoJfjljU/mT
sNNcFyI0PU7RySs6gLfS4FVzYZy7weBmb91Vh9wq/xzThIrwpqAztxXXJ6FD48aDmGeV1My7CiJW
GqLt/7gKpNERE/wtC2v6+UWrP+ZtrnbXsGZhEqK7XRzI6h4wSW8VJ9hIYGAIGVViherJhUK2SE7u
6f5jiGowDcog1YnnGKCdJlsvnm3HQQK1so3qfTVzkC6GXGLukwMEGk3+GPoFwz/jNDBFYteYMdUU
sMxajUQWMdOTC/1k9INxMvKqH7ctIHmzq+NR3FLyIW3WLOmFgXp3i+d6qMr04RtfkcLzzhMPmXr7
N/wJTyMTmtyssBMI/R46bC5E0x0oJNz29+GZZH/bcR3UgQHrL3huT0raPvMQ31W9wzGrEeHBvb3i
fjy5obETolggCwInDYdAe6A4mfDGdMNFzFaDjJ2mYvXoeg4CyEzQmNehW00jyiL61t+W4IeMywcp
Ssy4WYs1EVDj90RaqzkMuhZ5En/oqFu70DREWU/p5N/VkUaFdswfgNa+luUTVBvU+EUni+TYdn5/
K4Y+CBKT/eEqKGZy/VK9YyHmZAOwPyJHz1+prVEgmYk1vHTzNR7S5xaX7KUujBZ9NzJPRyoV/zQO
wF3ofYAQsmDyah4EbqSkVrrSZEiUhpSfEQIG9G4c3jtwSom5VNax6Bb8kt1kh0RVqj7PxtQlWzMi
G0Cq97ffRxSU+1qRF9jEX9byhY2UFO3bVRbl/DNJkoezpl74cZKKEdYEpDrPq8sIS9qCEY39nM4V
EySg4S6+eLlNXpzw7TF0VahSC2lvXHq961HeFMIzk/T/4SZuAmII5vt5G8un++z84jLWKqaDNCVA
V/XlIOCKiIYd1gHj+rVB30A3OgGRsXUPU4UkNS9gvzFG5TKGSPFGODEvrtmZyH+WjcODEyl/MaTa
LAIOUE0gKsftEcSQm+ybMfk/7z5KNP/cOW5RCN6nFzf+3LU+WBWrvTROTD9znDutokZOkeg3nzG7
NN1BmqWUAnpI/FguXD8vX6GfMRTojBggDwz7y13NTB5wkMiWA4cWmwGnHSwGdEj3BMKkDUvtSemh
wRklyhGAHh/9XmIQeDyTcyh8NiqufFfCASZPIJfF96hFLwE12fxtttaONrlHAIeDVVvxWADa2TyQ
iO5BXNZau8Hhv7KC4JJ/85ELePmLLC+yPwBIizThPhaZi/PO7PrVOM0dt7djTe54GfoB5l3orWO3
s15MU14MhuhB8U0oMRYU5gXbLRbYkysFaX+z3iv+Uk2TWX4Zj04HkWzxRCkQLNe7vbDj1/cdi1jr
v1CrZrZFWr+80nQJexuz/OJYfuA/zGqPGkSOutS8wU5FHcMH9vJ8lLKAadlWkWCH73pNtmO1SUPP
wtxssDXg8SiyihsdsyWxiHioBcJA7rN72EgZIiwUaU4PQhaghmCu9/KfM6klqDxnVsDcgOW3+Cyv
e0VM7LSlMGrhIYwAo1KRea78Xxfkog0sL5tKulZ7I4FO8IwkZEfx1700e7DrrwgXB7VQH3TI+GO2
vDmaIJRWUR8nUWc/ciAuldSQOTxi/uyY6VuOQ9MbejpFRgtyACMGLxQiieut5lL6Mae9DyUkw/NA
zuwpNzYHZxpRUcCd+yMKbHytKRgQBZpDmzojArOAq2iwnfc0YGmEiRLL+BdoXn24V7EH7WQHQD+H
EVPPSRMEV+XogWNbUfd3AXiOU/BZcrRz4TSE8gz3H6hnh5WfKc2vg8VpcQk0HTdQm5xfMkdAzGrw
EjDaBPgV9srk+524Rtyf05+Bi+N4itEy0uUav2DpJkI8iv4eAiEzXHN2A6E9ItxeWtiYA+sn8svX
QOaXyXyiseww5nkhyHJKMt9wB4SBGSCIoIs3AVdb5opRtdXiydUzcsP+y8bBxPpjjANWuEakfYCt
cD9NsdEYbYuBs67ddHSMPKS+w0kSltAfwA0J4DYq1Z6KtofL1J3iIipaOZjSEVWlJRSNsOBX7ewv
fKUvlw5pWKklhI68EmsJrqrniwfjVN74/GrFXHiBbVPGktLHoFuqUANycD3KVyWwmhYKpTOFs2T/
lC762YJTA7FuqtBybcn6lvTX/5fhmPCtvrjh/s41QY9kDeujaOdnYbEDjxgPtTAOhcQ+ZUubnZQR
vpmlgzTpBHhtakdBDCYW0yGEpn/QbndcMoQ+EGQ4XQcU02HsUH0G8FJs6B84bZa5SjKuuBo4d3oy
Lt7WqyapuPxoWZh+GvzRDmQhyRhYWXg0SyTyh7Aup4a+HIQgYJ4dhltozYLWj36uOhOOxxiXMTcT
PT5WhDNgzkCAYGScYvxWwCpmKuUBInDbaaPJThh3e5GUCcds9A7HDejPy3hFBPsWsaIXefLdMywg
Q3QnfCjm2BLtDnuPwiwlSweOglHcYVKVI5nLPlFL4XqVknD1sqQKVA2hmEdZuD6SDVWagb+1JptT
EodqEnJ+J9liCRYZ/m1wg932T3G29mXUcK7ocBOardP8YRh4KhmXmQlf+/YS2HBepodPk5BYBGe7
GWN6C2dlD7N8IPRR+/ZyrdFX5cRwuea0o4sQ83rva2WnYRWCIYEpr8vsi3WNwcWiIcdc4YozJIXs
KJpo+DyiG3HLVd73mTvp0nN5/m96tkWyrSI3luDAf91DhBx4sGqAN9rS/OaX6XoKnBvqqWUELgG0
7i7IkflAUyK3p0OCqgmlaOdtDD0VTLz/Iv/wz0MG9vCS5zWCh4/jA5fcJB49LBnpRwFxs1TOtL/0
rCZUyA9FnvesZkx4pncxFpETT7RRNpzQkgZscmObxOlmV6lJS/J5R7idYFLFm6HLQt9Mf+QoGEtH
Na20dlvK8Jv0grYe0a8aj95OZuMSmCCoNuytZ3pWWP4pe5JGyq2DuqxY/lARoZr6Xm1Pn5LDedZx
d7ds68iKRnj6fnt3GS3FAeAyZjpCuoiOFjQ6JYVGvswG2JJJ5x/Wq/j3b2Xs1VhvGVYF67CUYz1y
M5AAx2MaOEVrJJswl+lFpiSocnzYA/yWkkykkRpR9u83qhmEyhDxOkNRAzqr5WmIiAKXlNa4eOmV
57T7F1PG5lG72Q4L7IgkgTtH+IzbaMglRVpg5k9PomZ6KASelxZ7COlrZ/O3Txo+2kpRJLGck1Lb
TdhesnYEzHBX1ajm1yBqYk6l9nE/g2hIueZ860H6pxWxhIJwNrXOILdNq/TelZvu4TeU74NIHlxV
5sU/NXkdDEYRo5Eid0Jw5gJC32bQPvz5WtkmFGszMoMQUDlBAwgVhWuz8dr5zoYEgzMAxpv5wSwa
2Bf1MAiBCi1htVtbVIqefeA5WTm1Lo+tiCdPhTIL8aGLNM7DGJ2brizqAdIHx1nry11ViWjPcHCj
qkEI6/WaR1TPghh/7vGcjO1caHHEE6gunUFBcCkkOTo5F/2v6J54fTBWbVHEqypnA6bXSTnSd2BR
SqQ1R3ABuhBQgErccdizsAR/kTPHHJ3bX1triC5Y7xIRPv0s0acYJXciynqVBNxJTywd44b47/Sr
nJwAqjK4ek6ErGWI+hRAiwugCXQzJWNEc/GKYZD5Y3waNHrOJSLNOz3kFzXDq0M/VhbaA9a/HUSP
MI/bEIyMF9uYNRvcCp75xkDDjqqqywg1KhIIAAtvvR9PAJvWkdTG7oks+wcdeBG59CYqM3xgBgrU
CqIWA9/pCpFMBfFfvP6IsB1U8Kgz8jY6F4N3+jIFY3MlvSuGlP0alEILvXKoYnb+oskPbxo7ZICX
sjmZDEAQVwFlBeV9vY22HiNRrfPmKyxKXzLq/UexLpk6kgfHPnPv//CGlu5AG1+2tAWeQj2riYca
aAf8mkfaDnTO+w7b18++EFWKuRiLRwcDf+Swd+exxOurEWeAd6ehvD0VKSqja2CjqQV9M4HC6NmN
E1RYnlUI73chGkl07Y9KnRyv72YyRfFe2gRUYCW+Fm/Csg4WPbi9r7iUXOmZ+ip290wGlnYY/MFz
BdXUIGzzB2nD4qqFgPs/Zc0RKD0OmRTr75ONS/ncNT7eSbVveZXvnfkQ7G4497RQ4mwT45ZsR9rt
d1GsSWHOKxYFFv60wR4tVzgoh7AOP3dkCGeFpUqaaDpCuFhzUUMe1eBSPrBDHqOb7NvzUwvF6KjV
RzxKkYBr/pAiGllUg2d43ncfNRFjdO9QX7o1/TRL0fSvoTgNsK/Cg6At6X/YBEBfzu476smLgYY7
hnFmcnN99lktXuWre2jiK2ZTXUaeVA5biKuqSKR2s7UkE2OuevjzQDsrKPyLFc2YYlJ/SsgGa4Km
MiqL8w5Vmw6iIGh5pwm2vzAQyTfoSFk38U12VgzYJH8AevOLOdXO11Ldd7fmtJYvTs1UlZo968tF
ZCXShttb57ZZyMlui+tV5ZW7VUqX71TY4TWi0YGyqD2llcahZXeXDmtWrqziwE9M37SJE2mSTadP
X+NmRxJsCRLfkhVIXs1+Ce2HxM0E6Zu2IZrYcQRO+kV5p7H9G7mzWkjtKFJwHSj/J29ssT26YpKf
ijkvRDJon05fpGi9ysDsa55hXqLflX5/6e98lbx+empvrV6nucRZjn3c+8Bif/qB1AzZU6c9iyDG
NuA+Q5bR/ykqbY6aeq3eLOtpKpkiuky4B5gb4zFINRKujrx46YG+KFZ8ZbT5BvdXnCS4Y4HsMn9e
0iVUEI39ucs2MhMn/LQ47RquGtwz3fZlVStaABjDStKCYLO0SFCC7eQpDE463QIueKlKCCyfC2cz
WJ/jgbwRa9WN2fk6Rz0f6lO4wpHl4FYJHCo/QrgijiNp11RgGcY8BJ32N6iZyxY4xoR4Hh3Xkkzd
lsFT4LxkGMKF6G+F6/ybExbD+5DlaStMT/+/Blww7L3OfNbnqaAQiGuIsYptcwTjujC7Esw1RC7T
3fIhs8IteMOZGy+s6wpWJes6ALj+Xr3xFBHvi6WlSseQgyDIZ6v7aXl/dPxXZSgkRaSEkzl6vHCk
kUXFD0OCIw863VRtpB+0F0I3chCxskw975diduHuJarqT5/+edRBXkqjqiRowHCtg6imIkzPXUTa
9peB5zPnYhQKzZ1zmpk420Tzpu3rNB9X091irJV6vZfRwkIqtnfRi6jNEjrg6dEmtF+HEacpSvns
2EfFgS65AD1lQY+xO8f5m6bkCEXpkxnayskZZlbtG2rtaTa10LSfjhhR50/FYRLBwbDMhzhay6vA
wZ1JwQMh9+OL5UGziGSyDm1c4gBs1Kd87or8EisvX7jZny1i9/525N4SYIZVQyebzy57/FthrPqf
wFvvXNDCPQtJeMkkGdzHFLiy/am1JotKwBHS5OcOXDxpm56bjxWk6EgtGZo0txNaD5PXunfOtq5G
oJlTIAlAEbATiBqOgabzIavuqfJvw5DYBQrEPgSUQtP/DJsuRfef2oRc84xsr1CLgwcEfdz0W/zN
P6exSnqo3eQcYtXEeogx9ejJhjDG2nfkNiGJBUEtoZwMxh07/lSPQhd5WuabYBfxXvGJaDv2hP3e
QUgNw1MhiFDMdZ1Rdn7CfhnSCqA5WQISq+glko1RW7OK/7vP+ZENkdeXcau+5K0y3kxEF61CCEo2
okOn5dVJH42dELsx5Q/zIWJ/PmvQwhF5gWjOyIoRabK7Z4IbK/QDBLmMDEnTpOoyhmTWh9ejOAgA
kvrXf6VOiNKqiHfDAm1SHgz5sa99WB1k9iGUftz4MlDrlUTbdWgblPuRNXKaFnh4fw+S8WDc4aqU
SMzyS2LylkgHfyJNpcD/RMg3Z9f2gG3pLMEjsioaxajCF9GWOKz8VIVbd+Qzv8ePxQO1cuwqH+VG
MWnZB2n97HP3V7i3bparkwgAulHH2rpgzZi7pHLBITT0aRHhVsUFQd9ylriB5BsgIn4wWVm0/9gj
7teUOURAx89/4o99QBsfnKGemdvmyFIpNlVHKFQYPVMMXNe+VEAqtLmP9Yd0pKwSSd4qmQIXUSNI
2x0IY+N8yKwpSVnlH+68Hyyi5CR1jBfLSq6JpByZ6cBPIyqeIqeaAgcNF5diRfpg8+JMbs40Wcq/
R1Js3tD6dhqhvfQuENNWp3Cq/3SzAQo2siIhg/zANlR6E7eukdLo9q50sGW2MlaHrCdHbrFGHwQt
sbE3HKKegv11N2wJmoRx1kKh2Z4XytlJlddc42hNNe9tUM2VzE4WCD6RcKxmKakUNGDQVttvB+oW
gxToEYpvEmaoNrFbEz64jWRN1dZ5daj45ecaX2pmqay4U4/c4Habd6rIYkJVDagLk5uQL6Y1eg2i
WqfUw307rxvQKrvVm0fNLHvrrq4RNjEaeyTdQ6BrWSKOw2A3tmC0PtJpWhOTQu2vPmopJoxU/YCo
nt/91m5PfRUegrZnRdMcfXs1k6uAK18CzTUS2/pgNBnyCXl4MlB353rGnJDWBOUiHQOlBpFmO8GH
xkwPQ/6k6+lVMNcnaAu/O4nwHU5zsgc9Q0LMtHIZV7ecV63cZMFkFKmwQvQx53SB23Bcf0XGV9nR
WO1QEqZibJpULA135v1wZ3Su9IDxgQfWF1iHDqFIZlPvg/TO9mGlpDvzkM2WyHxCKQJnrm1IgmVW
9bB2XMH0RDdCijhWi1t0W/+3MCRG2H9oqa3jcpPIFlQ5RQQ+MWEQwktf7v6L4/oewvnLFs4yRc1O
8dRirrEz9HEDlj0AVbhwiDTYKGYIsVOykKieYcUnIpLSaroXa3TPyWPFLgTdyWatoIyAkc9ab2Nz
c8DZ0DYmPm0VsBg0DfA3WrkV7L7UfIVE+uT8ypO5PIEBZdWQ5z2l+7pyRya+WfS7cqcdh8YqF+I6
y+uWvxX3eI8hHjz73npiMFXKoXGWDsURjAlHHNDfSMHuAz4V8Q45PgHILvPLNcTMMgfY6Lv3aetP
5bIewDawAwhDT4G8Bd+FJJThh4WOqxQtqJEacmGgp5eBrCkmxQn3YQBqvdsVR3NhMYgm39pIfsQV
6r0d0xHavo0fiVOU9mnFwhqEIejqXi3rxm0pEIFOX/rjCdAUChvTnc5RYho6oqvy6brYjPgi6y2r
J2SiFxnUZuQ9q/wIU77J8DmkJFbSyHREDVkDPQtYykKoyjPovvbq+FnKXdFCL8Rflr9+KziounJU
m1cvYMdMSUli2rJNbdvXKv6KC8u1ZJatxZkpJG/v09XIGH4fCCwmCPNt5TrDkU06K+U3peUP8qyX
/JSZqgU+HKEy1Y+wz0dJbuan8z+BR7V+yY25H4jkVyd3yJmj7kSq1G4IfEDG7RWymfhRzgzK7tTC
amxqOI/zPNOyGLV/acGiA6Bv+O0Vso0ce/wO6Yeb5pnw55bnncb94ARfP8lewgasVsAJMyAPaND5
PvcrsqEO6NS9TrMT6661qPPbQZWe/R4aFmvkQAgGUAIzHPn4pCDjZip65Ojy/x7GOrPEjiQIZCUr
30TBwg+zQUwZmgbmaO451eHRVqydtlE6Yvg3He4D4sCA0qWJHeB8ehyQDx0uSr9qQtEGmmO5ql+1
bqaXU3BwMgLTVSIfctlsGJnly6CmjaFXFJ8PNZmvAK3S9+LcIJ984C6UA+pD8Xx2uxv8Toon+/b+
Sl6qypQQDQmvV81zd18IdtwUd9Il4ClKZP7+ozJL2z1R5T8kQLG86mG+g9z8On2sOUS3hZo0uECB
wR3LI1R4ChKpHDIbaQc71e3s2solvC1nOQFVR3toxCVAVgjbRR++OHb7zyFqR8PzhLyMrA4iK1nO
7MuhkUdOvH6tKKzB6A/izY8Lr9n5oLbRx+JEgeEidfyiaufGFGN8wGRMia7tbKdhlN9V3kT3cL+G
ukQA1XDhOMdMngsSuCMgb6FflRa8TTOuro4pTWYw+sdQHH2F0qldQxyDYeWjQGzkahwOj7Ds4fdk
KA3Dnopxlqf72XGhhnpEbZiFcEGVOFTJGHbj6eAKqY8aJdZQAKsfFC44qCmkR1LpjMg9Qyt+kCvw
t2DQsCcmuHC9qofr/OEBD4tQPqrd7vkmz+V2fzkP7VxdbJN7nfe4qyCjx/a7rzLnJnCTLRuB5c8k
2XpmhYDVslyOvD0LtQGtiSKPYGvgpO3pvOzMwOYPNU+zavpbYvtYsUoC/R2H6UQvmmtUfv00YK1d
NAj1Y6HOp/a+Xm/i49zQ3YQGEnL0W/hj7cbf6LXTHlOqDHvYCC99HjiSBrZP2dDqpVIXkHJ1LACq
yB9ThP1pF0VZB8xQn9bq4wS2sZJavKMZ9+EAcuD5ikeMCaFbK6Krh0hGSmPXZV9IASJzen/L3ZG0
9MgwcLx/sYeSzHlP99AZIXYP9GcPVCmHltwiqzVFdZkJzBkO9qSwW+eq67lJCHEcdf2GPsmbtp9z
8nOvudDyFC5z7MQSop2GTRBoBrdxT0gH5p56+ufVQfhFsm3X0AWkxWumFEt2Cl89Db7w1aTvEb0a
uFsXDLnrYXjWl08U+Y9GHhlr++hEoMKlFXKEW70HbUySQwBy4VqVBiZcbd50k7s1eyPtaEVEBcDA
viAo3M9mg/jvH0M4Q2864k++Pdv/VWd8Bi2ESW3sVnFD3sL0SbEggA9tNhhlZQLk28Im5ClTda4G
4KVEEQ0oleq6U07J2dM0aL1xiG2viCdiBIT5vufMfCQBxaQNaotfS5lJEP4pr/+31Yh3ptIvt7Iy
228FhIEfJKx68vU1leaBu0kosVipeHL4rxr00dIt3IYjrJHBc6IYgADaG2RfVs1j7KqTTNS1TR3u
sxe2DUN+m7LjPcTNyXm33sLtlp4uoQ5f4rAcLnUNclk2VCE8z7Rgvc5kJVdPs/rxZ2yd+ciRNI3p
ZBDeY5TRr5TQLY9mLPNmSV0FN8JuPegHpSNJK80ZAgYavx0HPVUCbf0NzQe5d2YgCwdetoCroQKQ
bUxdItQUF2ZDxOZErM2KkBfjj8cDY66z7LI073dgprgoFo0R4qOVy4ET1G+iKeLKIsFweKyn4Dzc
ReMSUJt4QMPMU4v7Uh3Gug97/caS/3ki6CWWG5Q0kTZ/CkpCvTnEoC2hUBtf6R7bfR+wIBd/FC9m
Xe7JJnQ15KnqSJjbnMiTWuALyaV0rFByFNSBfhYeCcFb2qhPFhl28f3Na05NNn54P4yI1RYiu7py
FwSgr352MZJ7KePMjxk2cuPPofSRiPBUzkO7ROWAMVRHRJ0S1MTBJkZpz/3f53JQmj5lHt11ayni
b1//pcN9E49qOoP9+OwVGfs3hLeJDHYOr897tnJTONBJGnrr4hzZryReZS0aEhw61KuagiG0DNsT
6bJkm2l4afZBOHUVFhudV9zydM72x1BFVFSZ34UFSLVN59Lew8Goad6OFJiPFWPZ0tzIzWvegET5
19rBJpW4iqY1lHmzdgIsVD9sqIANr3yf9/6SpDzqzZ2X921yzhR3hZwypE0IAXS+vWdaXXFh9Tod
DHA1yeeeQzU7J40TeNMn8o4Xgr85ozUZ+j9r+NOk2E36pKe2KdWo3ab6zizxbiTAPaHU+RSs/vSR
msMhR+yxhJi99mMbRlHNamUbF7TaPMwyoTXh2vOmR6S3RjDR6vC0MnNEmQejYOBq9iI1+13yWwjQ
1jmf6MufThJdWPnUqORD/cxRTILhJPFjPTnAIAz1O40v9GDyoRdw2bFQLcHbGlkfIzQIx7lWA6Qh
JINavlsxa+LIlilMdts3RB1tyEOGqmW5G7MoILVUfqIXwCxY6AwzScimtixJ8twPoQ+WS0ru6cDQ
LL58NtXP5yk0ZiD9mxYJSLcz4Ty2opEMmvu2wWWYnT6d4aqg9/TTVVr24MBPKe+5S4AIEGtv7kyb
xkuIiOgaqykCYQxmt5avebaABvrhxKYmWqjS/nMKJHP/2RtH5rDdPAdId3JgiytfPvQj305+Buzr
JGBJVmUyoHlvLYkUuwkJkiK8FqIGNChUbFiOstVexO8ZrHBs/dcLwxzpZmXnzA1NBoYR3VJSXdkW
LVsXLjmmfrIQxKlyONerzqHwLPBcBZ45QNUj6JCigrPGmIDdDAz7oGT5ziCagfIybjZtuQvZDiEX
LIHvD1/gah8NZt1Rt+X4StxHFbCVdMtXgVdKLUF0Ha8sfZIL04KmRby6Ce+zGM3ydclm4okR+oLY
p9P7x12GP2Q51wZ4Vrym89uGnF3LqpVCbc/gm+EfW+wg/rhUPDktH7q850/dhvz76bgQSyXwsY/4
Gds+9gz61L5L8TmiUdSNpYfNT7mAHSiU5drXe9oCjBXbAk77TCzFN9qgx5Nhl06DxjrP1i8u3ZmY
T/N0LXgYpMniPh/n2iOCBjPF1LEKB9c+8PefwujJuVo9Cpk8c4zf5+s95PhBOHoIg/48i9GBppC/
hg29FZ5lMsEzUvsMhNoGIC+ubelhgHWN7nDuRmL3H/w4/nJ/ESHGu63Llr4NgWH2Ov9jMx8cXbS+
9UaOT8y2P3X3pEtF87HWokWVF+PULN+ta8Pme5VuTOPXfhPn2Op2Fh8cKxx6/nI5D9N/UYeA9wLR
9MCQyu0a47bgBjKVF0YbE5L2KvHgPSHufZTaZ1T3sHA9dDAXwhZMwctrb/nWYURXD1uDBPaqfbTG
N/nXfF1T/BwGppbOu/ABcKA36iJlGDPfNJJlzCKE9Vjnau5bLGxEqbiiQwenyifRJo1gWsmch2fi
UAO6Rdw7OUTmtxuUN2OsRZPEAkPmoMH2j1ciAPEQ3QEkYGx0wJBT/F84Rb5duiirVHQ2IxSL7cwf
cUMveY94SNu1m/iJItIrDqc+iKoLML32/qGapCLnbcZUTLqC8tURUXMwfHgWix+BhK26nhhkZPGi
KkNO8/gRTaZBmi/mkOhbNoeoFldWS6Y3xNDdJxgIod9dlS1hBjjdfg3vnbiQdFbUU5YFh4+2FH5V
AAhaVersqO7ppRZqjRAnj/aRza3yEezJu+hCU6R0f3tVWYLOnK7bB0TEZvd7m+305AB2la0XI6H+
cnm/2wVmkqbvr8cRa3KVnJcw+gDMCt34Ghb1wJUzOFekT/Y7+5bFL5UNKfIPf+oBTvTOKHRFruxQ
pzSvcfI0LXHZ70qiD/5CcXLjczu5oAvTql7lepPWLKI9p1a44/x0tyJZL4bzWR1IX57kDTWhF6JT
iBRAYcwLOpNaWwHa8NQsAjYfkuEK4/vRmHdZDE83LPnHgeLdV4Y3WHpXL08ih4oau27jH9ChwOCo
YQfCxsd2BSD4pzeY8amWzBS3Oq/54wrlN07AUyNuEs9df9m1lEA+inHJv6MHIAdbzsstqsMX8lI1
fud4uA00v+y/yuu9jQ3acAo3/EQRhXvNCzZtCp7EANRe5W1IvWOZy1vr4EnCrN7xauvhKKJz7x/r
RDzkOPJUsTLmkWjP+Fm5JtFaPJ2LxT3z0zYRdYDITAKod7cSCB6Se/+p+70EstZve0Zqn88vse7t
9Q38ErsOPSqqrbQOPgQnLr3z2iL/qhxuuislafU5330KCEt7y3KDV1zKIg2cJQKzWiKdHMyMLql+
Z0gUQS7MWXUuVZsG8DwAN+zkx0J+T5o0vFrqiVRfwu3wJvskwdOsw3aPkvvzWUbKyScTDVS4snxX
Qm7w90T8V26o4H6dUsP5lfTNcGD0g352wSIn1gjLwqQlIQXRp7v3+EHiy3MKRvDkhze3s8ZDaRq8
rVncgXbDQZrcGKyYy4u2qUMgld8ibFMt3NNsyt+QBFl8kvWISl0Gu4CxToHSih013ndLgHlHbczt
3lLWwQb7QoFJmSTjkbjALU/bIvZ4ZgmuFcW1DH4pbO9TCXOM2R6kmg++NZ4u6EM7wwvNdtc96aI7
0KKPHYBsiQNuUIHtcYnEHu6eRx0WnKJ5nzeToov3O+hPmsK9oOqL5cmcZqnRouzPLFeI8Z6IfVKE
bTVY8YdtYjHKirhDbaLX/6xOMTwinPj0Ov9uFPXpojEUnIrJvKIuC5aNst/Kbel9XBMeG7TvTqB2
+08/vRwcazpozoTKy+bgBZq/9DZjFAt9qWzriMK9lCTf0v1PkKFMdzI47xTX1DmAH+0wfEU+f2XP
MVTqFYMRsuP6roX5LhY1DpdNSMgC2v+e314kCMPhiLCIbBobNp6fVW9fWyvVjgjy3kXIqbaUfG3E
F8PmbMH1zmXNp0Uam+0Ur2T7Po16Duz0ZwYTrx0+tWxbM0MlEJfAL8y0aQzGZTGQyC8zX5TwTMWb
8y0L5ICMOM4sjhPrt9npNu/vlmr/NDAyNPMuaSfOA3+oOo7g5tvJWbS2muBAUIE/Cr9BLlrzGQjE
LjOctG1JvpwR8ZnaWNHoxQ4m7a1A+Gn5TiK5cbnG+jykWjxCpw5K8cUvw3U5GhbqWu210vofBRNd
l2Rd3hxPRccAula3TB1dTrcsx3JDRO+ERtyl99ji1nF9zr3N/x1Chfc/FpsacD/IAmMpr5nt4ayg
qorefemQtli7/RCnDUhdWVKc0mr52lXW5X+Zgwz++XYMc3Kl7oM9qqgQ9Zt3Yvx2YfEYNtf4LaKE
TFCOAU86EeDHTH3mTgibRgiQQcQ2xutSgrdWUX+Rt5FVX2rwxrbe8b4SyQ/OM1jS8gXV94ulFJZN
aXt3SRPn5YEnd96rXNtZPRmPyQn/Go1TqZfPYRObGehNAFH2MdTzU8jhgG7hiFnULSRBLO12VO9L
Fo/h/QAZz7G+2UsDuWxG4tsZIDkB8WNHQpNc8au+sL8HsBmRvow92YeQ1JQDKKwdKQjrOwcMR74/
TMF8YDcNWmpkB2NUpzWW6FNYzy6ZL/vLN7hdcwIDFQceoRP+6F0rhIeiS3HM/XpEJ4QjRyyvsWL1
0v3lgLFbY1AT8djFrB9W2tl14eHMzQ5YK2888wTG6DYQnzMmhZ7CwAuoQMuXRdyHaVM5Xt+o6IE6
CVbgjH32F8r9AHvBOwFw7oRwbxiKMEyywB2UA2Fqjl9zzZr9WTtoTrVmAEAD3TGTaXKPn3kPuK9z
hnf1oMGJ78zdSw5aCxkI1TCyZZQM5DlB8Q0byRBy6ASgpzvEKls/PQLzNl+NGa55q1a01QQQTSqw
AEQNQUfSthYoU+VAgkXLpJV86WOkzfEC8MbOmhA0qpA8zUxkBqMHi7eqVMuz31qBYtXEur5VxKr3
ZSAgZPlbgSSb2nZeZaYBO37uBvDeWQjIntngj+Lx+5RQV4S2sEzwBjn3ja3JDtoyCrHlaVJHBrsK
dZvdyCE9zvw6oY2yhoCKoG3ynXPB2FkpYTY1wF07X8iMy+Q2kFiYOOe/+m+0u2G2rD5Rgo0P8iEG
cu6Mvsmidt8szn1GaHavTq6izQbQGS0IfXoLz0xux6qV9aR86YVPu3wUtXMd+Yt0iRbzg8nswnKr
quUDk2jD+Ygz83Ly8q+k7pxXyHnHSNOr5ksVw7JCJAdAZlGiKlQW/3n+XozoUhrDKB00AInk4y7F
oc/hUjDCh4AGIQd5rEYOvdEk4TyWJHZd2wo4BLAgqOj/sY8hLpa9dPeUufd8t9MaYq+JLxPH+lpC
ViQUBGh1Ao8I2awf0jk7ttNjAlLqKCf588xsP2DRq24IfEI6sezp1fbNv7PUHdyovzdOhXoCh+h4
ZZBfN6YRzt0WMtRNOZ3HeUpw/hhMwNUNrZwh0NLbIf52G33padp2xOsk1rovfZR982idPZtV8m1P
LT+0mPAq36e5dJ/X+cg9G/xYyDoBaFpYxsN6/Kuwk5j9mM89+vUoM8MXOHFIFmiahUrJihck1yjZ
azzSW1QxwOODySyVo5rgGRsmeIcdB9319lGAh8fTpk0+9a+bUbhj/EcHuonrfHL3btNrC8eF8W1d
M5uqVcO7vqwymxOiW2A6Umt9/A7pL1VvTZOfsdGx21sWe+ATbBHdEpwVyh7Yf4YXWeWT2hN4WyWq
YbOE8E76GDuYafRhnX4ADnD7a9Ec6x3hgrdE/Km0RmJ6sl4yF73YaaqadH0U6B0p2amktfkBk/+G
HI9CCc7uXufyizbeVsuj3oSiDd0PjkM5Zn1YtHkneJksUJujBQGQ+jUNfN5XWCyRjWEUSFteNE5H
s7gMyFx6Y693olUJKVdAIS703h3S+WaFr9yLLaZlv714rSxtPGqfsCPhrNXoQQ5I4B3fyltwNhZJ
m52KRKkYouL1rfvqRWjN6bjNhhqb4ju9DRvkFSqegHuhw2pVvv+H04KHTRtygi4LjXxbAgMk68Aa
cBAvkUu47QVyQR/ZMYdcv9lTtZRGxisrTEWHbfvFziehiTeq6MYKqhaYvnVrCgWA2zdFAPlBBo4n
zywpO4SG/V7bcCA5RupmsmOSu19xYqpAtNt953ZyEmwsnSG9/15EjnGp4V3h3lsLLDlQCxPl71CZ
bbzwU3lc+rSDYIG0cd23Jjxbqf0h7VfnWgAiak+u6ux/ROnxlYoYpU7Tgb0StFwyP65vZb8i2FZ8
yAFvu+C1WR91OBz/6WaZZxZ3pXZ88YF/DK5h+2aFToWfRe/YKUWHCb/93jIH1hoNtrFTzKHrxmhg
oSvneY7qM7njUDzxSggB+Q2gbZM4mcsXfrqqKRpQwlRz7PWa0l9RjwNwQ/oEe/GjK0HweviUoxXF
6dOFwkZYNW+fTDWiP5PvyFnqJEgWlZySxv63Iqb67j3OS4vAeHUC4wWVLLKOjPGqMchQX6mrgY8V
cMaVIegnN7TbCXvSRu4eaG7yZ0nCGjNW/2Aq6jwRUGsKwdx7liBIj3ZAD+JZsmVB3nL7NLePf9JN
/6Si6JCrVcgKoso+wNH5mEFZzQ/FsG0Uw9tg0Y5YNmGn6qj+lha8ZgLYgy7kMReph0ebYv3T9oCa
nbW+MvSo5FhOa9NofWw3ctyplih4MLz81AWvUb/ClQ/qwTIQjRaOz7eOKGhZHv98e/lrL4LY/wor
TbcXppdI7zCZ0GwFp803J+iPbfGtkc1NUTPtEZDgPRSETHAQEFiJjsALqtj1IwYpXqnNh6r3TrM6
/zyRC9RK9TlLf+iSbBq9Cs05ojg0anbqO2Tz7lTqDEx9d8i3WWj54Six2gYH4Qak0fi1U9v1l17A
a/KeyIdrKnzHPydDse9IvDyP3LBTWVWTzfn6Iw/ZrYIVVF1UHaWyizPZGKiGQjDoPQXtaeSjvPsk
mCFs6885L/9doOGexIR2Dx0lhG+iHoNYq7zOYPu/ZoYXKjfzMzmSQaQ6wvHAXKl5P+IGTaai0liQ
vncuDKzeV7/6sfiWe2dqBdKdXhDyHWdUXYqRByW8ePREsut4syctSe03mtaZceZNYh3MY8TGmDnF
1fOg2iNk9yjkmnD077MmQf8aD5n7/cGZ86sKgN4xa5RpI8iEMTrIZVEvzfIs7mL66POI4pyQEvFA
g2NWujTYn+BTH7o3tYz+KnMDMVdR8qiXvBVgLHhTd8Z/2xiBVSPANZXp2zDLNTGOWe7xHXqNBHst
4i9y32szbN+4lRm2iCujTGv+Ub/qJfxN3F7k2FZb006E+qtoDWsb9wKi+nK5v08nVrInCmCJpl8O
VK79Wk5ANlDdFKBrTvCMZBLTianK8n336wGn4hoVxnqJon4o1hFq9SZJz/GgV5UI2kwZ/LLoIlPE
wr5GjjtmNggj8k8klnLJZ5KzSxYioUCubcVembF4ttA81R8a3EEN3RdtpuZjnfg73nIYsV0scw58
Y4e/BlgQxaiQ78wm9It1pODrTboT1OnqEbvSWg0uXDRHCmADn+eO5DPlo+OsKVZ1WxRIJkgtM/Nw
ZJ9+cDTlfDsLkgKrnOddT5hpoR9TwaBrySzMjsvnfuW4CU0AnDitjwdEl79LrJKCeckMUiNV13oL
kOU0Nhb7QgHlDE7cd6F5KJ6rlb/nhEn05Jg9qqt4lV7HpDxcMO4IPPB9KEJCtUf0li8e/lrFldEM
8uLDR65SvfYVasU16JUaBteXGoOSgv2G5nJRTidUNtBBZkZ2bTdsfO5kpKGmK/RvPhjM0SUjcrgP
4GuRp8AwL+wrNtKMyHgytvmJIl9v3qIJEJ43zSsZXOf5+BHoQhY5UC26O2el1zmNLY6FjtjNzeov
fxsb9LoVQHf2JhcK9YcnB/PXxf0XkRQ5YYPAqwyx0uH5coOwQqW22/vjC1skBQhbktmHkaT4OjQS
RrCLEJDMXwKLhciTQE0NXc53VvOdkjNNUkgf/JRhJcfZtIXemFNLEF+Rfo9mD9szhkxxECLgu+Iy
qv5q7Ybkmekw/fJNBSVAGvD2IXj2wQfO4qZWdCW960t0DTRW+m//LP/3QQ4SOQzJFDIvLQIgrB4w
PsdLyoHg9pEkYc4TMpykZnmDaypjbDjZWCbZASYryPumvZeAJhCOqSBG3M9pzTG8y0n1LlD4B0Kk
ZHeTOHzQ+D7NqTfK6CdXwLnbM7n5o0SiZ5Qgn/JlWdbXYueabc8AYYncx2HKx5dSFw6eSn2XG7J1
lGAbFCR/jm5JDqjrtZh/GCIGHMbij2eURcXkIBbYozTX1WU9Pb2nLSDHWS+2xF+WdYD2upEj9dnc
spihryN4Grn5xI7LGeQWvKcVUXRhSBsLzPkUwMB1Um99cUvxBgqROHdkfVSauvrmnFZneYhU1A0e
9W6klyHAVoZ9aW3aisIP+mQZVCO0FUYvizyGkpSTXUuFGPtBnNAMcmANfJ5nWmu0FdmM4IUzM41k
xlMZ03feWypGmejWd/9ho/Y2GQAh1wRJ+RWKohEu62rftBqen4U/O4gu92z9Cum453pi1jVr+ev5
Z2nhV556c8ZTr6LZtSGocm7e4zSkDVYqiFR3uTk3WWN6CTKjRrqnQZ2aU8ppsfghnnQr3C9l13Ea
8dd2S+/ePqipdqKUWbBLvJwLepJi8hEDDcdUuGvfSPI+7UniJ46nWW/J8sgQkghAkkcfJKQ07160
VHionWTJ3dnnwj9fjZ4ouWwDJf5FLr/hTcVDxw7gbEVLkoYKbWlHwczUcGWajpqxPGV6K0g553F6
3IWKOPGfKpfv0aV04lue37zjd3EsLzaB+iDkWPAtnevyllA1y+6xJRJ6Qm2cOSsGwopX1ka8+3MG
BK0n6ODep+GU5Rx4CPIWDvyKdEHhsVGHRgne3j6NIHTCESw01fXu8WbvdtU4cTGfyM8EIfCmSs7X
jaIaNn91U2T6XJ3IZ3WytboZZD4BPOM4utQKmv6w3U6fGuFGoWFX0KbfOQLmBHwBonYZO5XobThy
8x+NzdnzgQXVrS1tQ8v5C9d8wUbiyz4ki8Ry9uK2eTSwOgmDXXFlI9oXRE4MaoctjOTMSGqQiEMM
vlqw6hZndxYoB7yxKZywSFC5FKCIy/lB6TBnZAcUEpRyLrFFSD73CGdIvo9+EcgIEWyY+wNKhkke
7mwnxj4e4msujKzRhScGFQx91QaIRtMfGgmC5mXBRv8fthB6krkpyA1sbVPHf71Uw2JqTqu4lOxC
4QiVa/YTaFhTF9Svd3DAMp5ZUd26pYvgJsuEDj3VAaJQDg8KUGVdSdbGFvuOXkjMdRngpUCWDpOo
IAKScLmDV8/cav4noON7LOtVs/yLJ0b1v71c19XzOmZE2E8QPRTd6f1tSwm2xobo/NpTO9VUsZAw
QGBJYMHyahxgeq+awGH2Fy694vqA+s3zNiQ0LYKhU+w3GPm43TyluqCu3BMuvl6pRlWX8NN7+qqW
uzOM5dtOByANtrefQ6qBVahP3dkbdDEzfWyOqKz1nveMu9mt8MjOzI4PCUc+SsPbxP3dWvjS6R7+
1CuNlBjD7RIG4BBW64cJCecG7D4TvnEfxEIu1jNAfPaQ9qouSxA7FE6PzIOsfnBx0AXYzgxF08gB
1F+lNRVgI/KUEYDt5sIdh6847hCdPR1gc2EorTVPBUpVgwzDSxNRMnUa8aLbHqniHkMfcwJH7X4q
OM3bHNjeX2XTAaPfVtRUaBoKcp3yVQesK2nljnCFQ0Uwgz3zCzmbXejPVS/CRr1wr/AtTVZe4Z+U
B/lp6G83coE9vSVC22goE7nvVK+Rlk/NQLTNG72wSAPySZv6MxTydNyA8y9ZFxBHONu21Rv6vdHr
XrQ+9peL6on4Dn8fSQTRAxu39Uj2lRwACxzrYlDY1pl42+k9Xba7OoRczBTC3gTBbGlIAGg8uO6G
pSFUUETFB+ecdpKAtbbPeAM81wJdhTtrMqBoTJcaY4tObhSFZA2R7AYwE5j5z4HX/LKn38att6oh
s0If8PWcFXwYPkIM3OHDXxT1PFfMK8xOyhji2vpF4Ku3NQaPd/0xV6na7VQsmXJObyX3YjsA6/JU
eytHQY4CxVgMx5aDpMzvQE76PuermON1F+CQBItZoR/DA94MPSdV3D31LtlZlg03RRPGwQ6ViKww
AryrDgiNaRm431BSe+nDVL06M+dKR47Tfc5o7mLq4akotzh9Nc3ckhlRIgFLzukW0bIPBmPOL64y
22AJdP6U4EhlvTbMNarERJ2YyV4bfHMgL8dHbWEEraREp4bTpzGiaeObQdTTv9yz9WaQhLCJQgbF
nJsqiVTGKZhYfApq9Jmwk/nIXLw2jBZUrpBcYLRmQDc8b/s7Srv7GN7HKJsgL/uzX/u2u105O4wC
ETzf284j3vwVVv/0kPLqIQ+FNro/l9JYH1M3a2fp+Y+uwuK+/spe63STbj80UnKH2OhXhzYp+Ddz
M2HEFB7455JYrGkXtK8ZDEs/8rj/vSlT1TJymOjmlS10FBTYxYqtfBs/oVMLdyFtrIVWUiD41dIQ
TTvXrdSnPrGmnzKiTHqfgH9Ll8QRqwIUrBPOxN4QmPPf29zmI35QTHBnSe2FW3crjUZHE2oVwZWk
JbqVLB97Sf/juB0bQUrCpcZ0AXUewql5JLPe6gh7peucN9f3SZVDsRloHX6p0wm4RVF40MIVPuYt
Hz/nxmQqX2wkfTITKU8SZq65j1c1+Yb9pECZE4mqn6+looxb+6qzU62zE36ynfuTH9zev6OCiRRh
ySDLYa4izwlhYyXG4/Y9VoL7s4iJOsAoU9Pb6SFxRLHxPWi9KIBArvcLExwSuNd7onJ2H+YUIcDn
dPa/MfScRT1QzU9nZ8vfyF2rwZDVaqSklhvNn1JNwy291XYFOnWGS16qLesaUze65FZlDis/M7uy
EzJMHUsBGR6ncwgb9jrzhTuRSIv0QmPRz7m8EQLp+O8ZXt4vdh+EtGYkf5YnqDf9If4z7tgZGAOD
D82zTnBVYXEDMWQS/7f83NOMTn1/LcjLBLDfUpgf7QC2Q1D0I1d1Jp1XKQX+XAKNFbi+I+1+mc6J
NCboxUEPlLBCj4ZTQ3qYBMXqMnatgxbG193kWSu+DwXA0qpLUgNysyga8AND9tenGDoGXmUeFpoz
JjDI9nck9xvW9tnCEROsqsP19H3nem77sDBi2Imd5JT3ra5kbu4b78Fx9LbyNavXdC5c93Azzd9A
Y0ql4B1DQKeSkMlkPZ3nQnV3xXtvgFOdoPUMeC7tB5tDK93ZEXHD2ne4kjjyuc/I7XOC5PPD6w44
oHmcYrC98bjwTo48BYT8lZb3HFQ2GzltpKjy8SdrTX3W3gwcetV+1t8DYOpsWe6hU8L43TuSX3wu
U+6wUO78+spuX40RRg7dOauw5tDxnmwooIm31/xUkyNEnQf+RLhmDI8C8j4HEIx9Zsbp0RFqeBXk
HPHxT1yTKbqRJgzXXr/butyrYVu5TDgKRRojKuP72FzMDO7KI1DzYwQ5DO8jxwsEs543Npc9f5kq
696QvC8a0nPXjMemPeDfGisqJrAvo1HnchO4JYELWsRAJbKwWmm0dJi8/3ERdpK8pWQVn6POiyUB
EGJ05HsiMjHs5df3hRj/7Xyu+Wd8xohmFGD/6/cPu56ll1ZIdcBHTJHaQHTtQf5k3WNZbLaCybI4
XyvvThzswV0dyUp5ksInfUxsfhsFNF+be+ox1LAAkYT7cpwKf85UUky92z0xu1kBP1v7fXhjycl9
rSA0+7PDTsqp1jVu/GCqc0+TPOFpItt10bFzsJPBpVAs8MSar6LI17SmCtaA0AmL3NykR6xpN8oO
hkTCrh0JVf6LQfg5D7Ng05UrYgoNZxeNYNW+eaSvU3ndmzjCYoLx7Dg1FSAGbhGuV8xYXRVHHOk2
SkVRy5lllzylwcQPYBCxA094h08i2fShHPvETuru5Huwv2mWZALCs8a8jCSDCEXCwW3CmbxbeKEC
esXUpBGsBJhzOLOIDkfFUyg1DzIAWth+WV0OVw4r6QH1OnFib17cxGhb0bBJkTVZ81uUBaq834dC
wg3xlWas6ZrZlAAANhgN0f3yTtgCcDabHbSubxbPfeovz3aHa7K5rrD8dSISsgUfU2027WDuXuLk
ul4FIZQj8YDa9iSOB8e9H8oL6AzwWsJrQJCu0yNoBJfPsz73PLHuLxNHH1lgEfJ261QBVQ6iDoom
kdeVxEzL+iOcFycn/xPiHPTe2uPimLchuZi8qn9+QXvTDZKDv5ad6kG/xGf3BFHVKCrDvpp17GtM
Ec7oGcctM+gB6G82JUq98yDeYcobt2Fe+mgIAeuGf02ktCvCOg8ageNss6HzfGdSTYNjOBx567dt
a1WVClbhk4+BHNKQig3RLOzCJ+9YdBALdX+NChbXMcB+T10Q4mpKeqHw3SUYSKzmXALJp0LidRd+
hpkf2i4QPmNRBAECJT1W3BZ5tDg/8hQbeUzZQksMoNInN5V9ehzaVspgeUia+cBAreV8v6poO1Yj
iUMeaj+2IwFPqn+zMmYbJzZ5DKZJ0id6trd5SejPIUnCraubMixQxGEEyj6kC4ACwXgMDLlVWgAL
spHej6KQWlogO6Q0QD71G5eFMwBVClz6LBe6g0GhfkPvuxhQnOIveWX5+aFf9CT+HA4Qy2fryty0
/+raFY5BJZWKJ8eXiJRMfrgX2WIvmFPWfS3Y6gVpKlZL37JScucW33st3B9W5JxD1F4p51u/9ndl
9/n71AiTXG8AUfDbzFQYigrJveRD2abEnp/cLqWc3DcxPJhu9wGzfw9natUP+vUs7FQcvkKYlRWu
46srhTg7Zqq5C3ibW5yYzAzUKeHpHQeLU7xjShQYZLjO6UZQXgYyf0k8W8TnWlL3NAUmG/ipld2T
BqnhIleG3usl0YbWzDYh061BVvhE9kPWqg0bWkn7KT1JABny9izDI0CWRqOsOd0+MyNv2oDDUCKU
H1rvYDduaYQboN2qB7k4GusLTar4pf/c+/bAFgQ7r0V9GFizupGYYVxMoHkasBtzYlLKXXJBeZfk
rPByRCUkMMmhG2bwM3uAT+XNZrCl0RySxn5PFv1Ij7+qmrlJBiqHF/wvjsVzMbXa0BlwbQRxUDCF
6u/D5BnNSG52ydKTVKVbphafm4m3ZA/H9Dw1ZvSjjaYTeQNUbR48KBk0+2GLTukfap/GIstVMs3R
O8Fg45cEd6kdEGBQlbkPwWjSw8w3f7EvoxkRV5gmhUHZIrv1eWijIBx14iiIEFpUw4/0kXtJKb9W
q+2sg1K9dOCbYPXzxGou7QJFxo368wiI8/IaXaNqA1oXGi4v2i2BegyKjelJ54S4Yf8Mnw3jNuaC
+lDOl77qxeM5PJhjO+N1BltvfKow6Mm7xs4c/Lv57IluxmTXsAeTMDTqBJuqyWbQVYgEt7AuXl1v
lVwomSjKMEZL3pM/D6zIohTuDDavpBNZj7lV9O+WicE/oVdF7nz649hLWCGatPqR0+Z0iCHo6+E/
5kVwVBrwWtvji91hWUXWf5QP6pCpVRnZeg7ZgBX/MYwLIB4fRaLR74xwh7jJnAMLH9o+vJvh7Y8i
SRIiIfoJwc93yzv91WmqDxOG1C01wEF3WKiyfuqWF8sgjbOSuw2hj2Ess9MZIJrH0fBVgTqu+9yt
hkaXw2/iRyr5lFII7V7zC54QqYsbXi91qNl4UBPBIJv1RsdUPCT6KzcdXakayoT/NErl6/1zwmMv
MFx6YpqXiCyvOfzaipTyhlr9r2OxVeSQ8guiMH5V7xY/+uKOmjIEgx17FQKhYT/FsTwguG/QEHrv
m42D6n1vgifXnsQhEmMexc+fpeGBKkBFwJzNQb9glkq1wWSMHIFvChyYaDtWru7f4u+cPKDvgTqQ
XA1AxsqXCpeUwrffmxWJ8qTAOg0wI6xIrUTGpeeZIjz3+4BgjX0LfCuiwzUktolgK90uyJAjcLTF
ei6fkbImmzdFSmXF1PyWH79gtGY4t6pA2eWN44MvmiFNBpDwIH2doZmim+G3LQXloFI09yEnYITT
XG9ULPuTe6Fyb/jkCgnQSi8GbfUh84FfMzRintUcPieaUQZ0xWZiLp04JfmU99FqyWdJ+ZG++iN1
zUp5hZh79RjSxNVVinUYGLQd7DkK34ctACse5HvHyiX5xr90Wppy4txqz1gH42n8m5Cs9p3748t/
xo3hVHxlnD+dvdy9T3jv2cnYxo3Ey9NAZab+MxncDbptIPkZ/Q21OzYUIX7QIxNLuzfYtzrxSnD2
y+njyucbqMyvQt3xLUqseEe9Ntu7uq515i69LPZ2rMj8nGN8DHv19K5H/pqbvDumkoOgty9ozFKS
Nl6ULTmwNwnVlnGgqpDplhhyjbdM5lI9sBYgdtA+KPF2Az8UI2n7horr1RyWbFlZOAjk+qrKfeOh
17xURKNr0O6cIJ9QSFvi76+pL2d6D+rw704yeaKLS+GYIZjvpSkMGkk5JPbyPw3DV5t7u+RSPqI+
9Uv9cYHnuONt70v9zII49hLxdN+GG394rBjZGhZ8OjU/000GX22Eh9B69cR9L+RbcTQvGkvdqn9R
bzE+pRoSJGTwa2ys0ZpEVAPlManx0Pb8ImEIRoW2PbbFt9QrPaS/pPJtbkXQE4Ro805IPt4QaIFV
A8OdXhmfhWAC68vNnmPtRU0nPszSV8r7dzumS9nur1FQVEHjO+VQNvvL/OW82GAJoAodW54TrYZR
8SE9kAjv5JiXbYk75X8zvapZUhAD0e57tsHDTJ/Yztl2z5EuM9C0xlP43gOAa8jImnJLvo5LXNkL
FL15fSDIQz3kz0r/tU/Q+eg0rj1+DzlhTp1ZuhtXaAxh7IQPwMO+jzVaWSECDptIZxbyrBq5XSwZ
QRPaAwCryPoL0oiVuBa0k/nNucSi7PWHc/oUfyW5wQ7me19hb5gzCzUWIOnrqZZLQwbqHAeHfdK3
DzLB6hOFcxJhmGjcwEPZWp8xsPntEratVkbHI9zPNdtkwYw6lwcmXDIzv8SstU/HD0zO8SzUIe5R
q16aR/c5hqvb2MJd/LcBicUAuCUhy5RPKa/aUpZaS5RL0AlpRok7URHOrXaQfNTfrM/auje+Yp+F
/N9w0j3E6JsOKWCdPCXSoF636jrKXjLnUMgafSXZjae0TjewrRWAqW/4TcF82DuO1Htvq9JfpG5C
qdWlMfSjSKPzs4Z/8svN+6ticmEZ+GxipOxrMvzoyuF96EcBlfd+wqGgW+NxfrH6j1O7xhhvgRMQ
ZhqhuqP9VK8wqJCaD5PG8DXk1CfZsyPZ5wy9n2rqUo7leT9go8qWqjwzRCpS3gSDSvvJkZ8hqvuK
9Z7CXSOOdjE0iQ0ee4gwSJlabbMqcLN+83cdbxqszwtgazBXDBsFu0GvfzwHaAYfqyKXsdnFUu0k
RaoUFRFnhWG+brIQ21DuEBUJ3NF3GJ795vMjt4eLJeJidnQ/9EXxFwaPqFwAHTMdf3AhPDDJU8mR
JFN4FsCKVqIFTYYCa3+Gk/zW6fEhRj9ZKB4DCjXLl6DmKQX/rLS2C4TO/y1m266jB2H9TjN+bgmA
lxkFVhnqXvJfOlOi2HGaTBeTcFifU/BaevK+dVPzKtl/TmImkDjUbSw7c5TWNtQauefe/+5vm5xG
C7ktBExxfWmv0wF4gcSO5MzTsyfHcqS07VHteQ+ddITx6p610n8838wstGz3QEtQWenTSddZWerd
XhwvGkq+iuMsNMCdsgDFjrwKTnu8Ir378dTquCiN6FQTNbtHqA4VD1wqoygbDoMH2hEQXVF8+8ze
LsecQJRCEKCcgr0W4XHpu+MGBse+8djZq1KXUCt6iBlxAzkRJQczeVAsSv2hpre8cRFt1+gQVpkQ
Fs1gpZAPgHtJZD222F7bm2j7em2VPIXooevC16ZkrhTQALxKivxw9xDGiOIEqBXcuZW8byhEnmOO
/5+7V2n2AwtEkDYR/fRPv8KopvJpUhTsyeJRlTDkTdh02ndLs/9uHRftdagKoTAYCKWAfnURMU/g
O4G0qBZkIfR1FF43OHTLidUgKg3+fuDb7NQR6inRwZKzMjMK21o55wvIXovarVDayvD4LPWsOBAl
nxaxTQdBirEmVKZHwdNGeQcWCI/xdUjTB3yDj89sQCWOsP17QREkkC+uiwR/Yv+iKi3ysC0Xr09v
Kg9cjrpIXdiuHAFDpuBjEOAlJheh+E3XtlpIyfQLkW6NVtFOHtTNDoi/QeB8SRqEEy/hA3NBvLYH
KwICyHT6ihUOmbyy7iNK0jTfexwZQkYrWTHG9UKFmnotSmgTKgOA7NwbUi7/WEzXKOyA5KGT15xc
3h8YkgqILWWlQ5ql84hy1MFLliWRP341IfxuXw3fASTpE3lb/ysQ1CVhXYg5y8guhf961G1SsYUw
o5NZ5QKea695TaiLpEj3v8S7OsuY3i4RR9Gtp5VAl18K6bH11ag9HhJ6qXz3AvYEvkkDqXtY9ldz
Mgz2UbP72docRqBZm51fPkJaNo8tctWoUhTON5JWoC7Ku91W+e0HYUIxl6mILFmwalv94DiNtfb1
R5NJ4lXaRsrMMUqgpQCZQakkqeKHb5PMg+bOdgIwKR0ZOS5MNtq33KjlTRxf87m+IDqkxKabGS0v
VRGL6zBuuLxcI/qBjgutmAqw2pVTzCeWHCTioF7jJcSikOD6/Ou704KyJjWtWPkBIHr8Yy3JPJVz
S5J20JvbgwO76GaRCwGfTCgOzLFOFXllFrQ1ZcO/y8vVyZPPHlqRfamAeyADYFgI+3L8YDYuXsB0
JZSvbqTKYGmwfSHp4x9WwI6EWMkLteHfVp1YNJzbXgRC6gMcx8H9/3S+wEhzBM5FH9txdltpbZax
XnHCFyDiJ2mScHWT4oGbXs3xqjeY0sl6efnqef4hQYrteAcGpdmLSaO8a89ZqWNeAe7x49I5fdNq
WEO3mYfoTP9Sj3kkxjAuP87oe2ICVLPucSa4YcHi6CsulNWsQwTlf2LkTn3IECarRINRPCsKOkA6
uiDCTw7Ko4A+p1tvTIdfra8qQ3rG8J5XntOzVn8cD/vpsKzZq5XbfI0wZ+1ua8OFf26aOAWVCt4v
bqbKtmflv9t/HG+CYDJE4oR1cCt+Fk6YLIfWrhu/8JGUJJCe1lt/c1jGf5qMf9T8vWsASt4jV9FH
DRwfyX1Tuh11XW1DsLnY4ORqK8B58xAg87wXUIalGJeSJlW+9ZiR7X+3yBBDVB/A1sqwgGbxbOis
VgVkfow4vDapXZ00sg13EL78Pym4mNGxGDLen2QUpUAVH9042ixSoOZrww4Bqd87QPln7SW45hfn
MPRm67/obK+MPVoUDSB1i15rjGFL/O8FvjOtKwQKRxCxfEs0CNrMraAmscNACOnjbhVoAklKPnP8
G0lUXimc633+LJERQGpHyG7tiG4C3dpKSQzihVOq/AZvcZzzNxmwdStwjlMrhdN3z+aoRlsOa0Ay
pDweJCu7Frfczcm+nK4ouQOMKgNRPWdjO2F8d/v6LiOvJJSYNwthO7zg+SnwFQtGGaIDPyIRNBHP
u8odhcm6pBaqjyGzZGCzbQdtk6cn6CZR2UV2os9TPt1Za9hew6QuEL29WJHISss98vSrUw7FcsAf
XNGS6TNg0qnDjMMqzjvZ6JX7QOp5Eom8UkSKyNOx5s5jeUhvfFrNdEdSugyad+887rmY9jyCMQf7
5h7L8bX5DIUpsFHd7VZhTZ0N8MIZ2lLwWTb+uaTTmx96lDBb27mSl7iDehQ7dw7XTyG+SXTBpnre
4Y3PMSwOG7igly9+R0BNRynlxveDlv7R9CEMMgyHVqEctqIN/yz99h/922zi+3gc4VOe6jgpohSt
eyH/YotbuC7AE8z5AUrg4A8Dy1OADcnh3FaM/5Jb7zQqbyHZQimeNrbAOPyn3h7KuXYMsNPsiWQP
RqZerYgz0fkQ0iz4sPTQBGJ4vRnl4gkwzXyOZZBg5zS9gb2YDtaWPasljI3BGYsgBqHMdKt0nk4m
FvKl9sv5MTudztpGCwxB7Wabw4jHtQHpSEXmJbwayBUnTVY51jHPoFdPpEo2ybbAAxkXT14yik/R
05TzuBd6N0rnNLCXfIf4YN+9hBPr4adP76A4nQmeROFtOrXNAvJcsTzJHMULVHu697Z3wJ0YpO27
VEeFAoHcHPjvMMJz788iinrTr6OLAoCrOIUlFmyV0dp0LqJfY28OEkxDyGis2/LhADu/0BnyeYHK
3lWXiVs1I31Aw1PXH01QP4xkJBg57hqv+ud0p3xJ3arENk6gcfBinQ45LXA2mc4G9/kyscLUGWIV
56TtWdGpY2Cj5HssaF5UvcqcaQcFXPp/fKHqDFkzCYhi59WC3njVz3GIXD7L68+zRx5azgBiSuE0
xEfP5mHuPVTijq2I3PxYwqg2ybkgg/e3AO2AygrJaILXgPGvMHvnr4I5BGha0eiHE7B9jsGWvKyZ
AVSCnjSUkUXkPdfYiKiTSQ5ulgtsKNgGVSl+L+SUHwlecilxZZ9fqotVe4wTipk83NY+4NXlrr4r
2OOizuPz7swdyiGgyBGgrFYbi7qqbvJX0HypU83zI8EpNPEokWzVM8wCIA8cAqrN0xkSuRUGE8QW
pVun3bygMCbXioczXVWsB96MFozuugIYy+XsY29oR6R8mvkCMStLC9iNeEMB7m/emPL1C2SlkzML
ql7femJCHUGQYxTcDfgn+qap2HYVlXWrugik/oSbXek0EhCMdNyekEKnSwDtByA/imDR1KPkn7g7
15qXAiYQZn5VPol6Rux4j8zoLGVQihmhJnE/SQNAwbfnUNZA16JDpGQ0SWRRA7JD531B/XiKS2u4
UfO3onZ8i3BVh7+QKAMsfyBUuuXMcIW6CVJSvBy00EsPzuVHm5b1xTLxlEkmSpaqLNAGs0NiSSgn
CwQ6ff4N+jH8FO4xVGgWX8Sd6I94hvGX6B8Q2SLLJOqrd8c5SusarKcnCzQqpNn3jYSCDL4UUl2n
e1UBgeqoAhmtiHdWXmykyJZGyH++Wz5oBLoR2ieYS5pUNYhYcPaQXftpzfD8c+BgWRazQG2N4fnR
ETKrMHY1NoEWm2an22AOmLxxQ6qazzUPGA/dWKlNWysQU4xa219/jk5e0g49dWqtvrMDYOf5Wm/+
2TsJVtJd35EHjqxkS5Br8SoTFCc4xfwBJ25q3rk6bP9zKnTRqZZM1MgWDimsG/eeFYOuSmRwpJ5T
mU/1ioSNvdOrBW+xpxowgI73/+NrFTPeNZDbAP+irISBi7Pjrk3TJWhBwIjq5oMKaxjXfTB48leo
ihB8luXKfl296knCKq+DrPbh09B4hAhHVy45eNVHQptuNreJK8Czays1L5Jqg5zvJzr3X/scTCZK
Ouet/ed1Wp8VSjMYoOqFuF1nFf/ISki20W8g/HPY01eXtqTg1wmCSIswil+7iaDOvcKYD5slpdUW
vadesoEDOxxx3xydxvJLPYnAJppBD5/4/H/bH5QpPInP94GHo3SGoOF2UFFS6JZeZnBS2BViai+x
uVdsTcBKBXvQSanvlKWyIBnNR/amRxrtbmubxgmjDCv390DNY/zA9oayBfMGEVwUcZthCSWXw5le
Ki1X4ZaBvKvxSGlj/KeYL1duuD2qALgt0+TP1sx5MUaq+GMB3Wmx5fwtNdt9nst3bgwusSop53Td
QWrW59R9DgU7TTBt5vWW/sRtijuaM6XY+dJz3XCt11kibCEELetr3xWarIydTMF2CIwBTZGQUG61
1DOdCgONurkNLDA4s00KEPeqUB0xElWh13qF5Mw6DvBcoeflKnIpCVina88b/rHf56uB3rsx2I0x
y2YYlkr0VXtyBNpulhFxfZu9XEa7TSyHx9U0sA205lBuAd7sNhfplJAJP4nWabn7/oOrOgyE7StM
BSGCTE1z1YVk471wcFxv+5qLyf3gb+/Iw6UwlayU0y9FNDQzh+ayLbrQY7zTimvRXvmqu+ewdMsX
OeCzECr9eQrMUDrJ8jw8ON4ZgB4OdtLYM6F+8dMc+OA64320UoVBNrU4b400XoLiFJrW47qdRXSE
gZP7N8RWbt9I/AFWIKWnmpSexXxSe0fwOcJClfMLNVa7iWx3uKw3yD5S7K9G6TK4JRaiiyLvdBwo
y6aBzQ3vNRYQHN2rTLVxfQyyRb7yjtO7g9kc2qNWZDEaBnXpoWwSQp6DJ5VoqbzcQkjaVgFBYnPS
rh8e6lIdH13sJqNm77JKQUrzS9jyb6yNxK/CckXwiKnkR3m1CIDwqCH3IyEXytRPALHlFuU5ECYV
exNsomn2GbBskKsK7OOO0T17Q+z9lhNTIL7tu4Ni4rx/qK05TzUR2gSkxxF3uO2uTdsbOvnbDxMr
687HKoraGME+h3Vy1gLM5wpQijyZpiVlzddI9nNc7c+ncC/5xKM5oRCFhLk3Fvn2GgCDe5443NXv
V4vz+bew8RF2K/TsGtSP7XJycpyjTfh1hTg69jv7IT6AtN0NSpgRuD67hSc+ZJNL+IYw3nZvqi0r
A2Nx+7S9dTJHq4TFYi4vfos6T4LBVN2nP7TJyJtx0OKmB/Ki+ey+2leB/CNdHXj3z7lG8dGaKg4J
GcFOc7bcWhnEvKn0BDGD0dftFxdEDllOSfSHDV+rgtVS9XpQoobLAgaLfaXAOxaRnHS2Yy66CB/W
HX2QZgTv1R9ZLytpcgNw0byS0MXItT8bA0AudPXfFm/eYCQKjpWLubsf2H1ZDlrTyihVbrEVoekY
dsBJnigB4zMDtyp4WRHrXbd+fqbrduUMb1PO291dpbgtMTAt9d2q9IThpG6CQWg51tMmY5rJDr6A
71zLK5T+0OX09z4QEKXfWA4C99je67Xc1VUHlU1ff4Tgsqr1A9FaZomRp7kErifGXRatC5QeX1mt
bWpGyQ/v8wZlqXMaEIF1Yu7BiYN2azbnnmBPSUfOpGR6y1HCuzNFFhek+4aQPOGfB3xFMurCP6n9
KEug+CHrkY4FmS9g1Y4P6XCr3froeImyg5NujkMu9u99wnugx3YS6ABdXreZabd3xC8/vpysIY3K
LOcQvKNXZOeVJR4/8wcK24X/8OCl7lUNR46iEewEI3lriB3fJh44RXm3qxSDx8vrHdZ0X/udeGv3
1TfD53/6P3m1vJo+cKUMShSlYwV9XGpsi+dr+Y7bt7zYxuayC+6WgH3vRP65qEMGpbyU45ue0ba7
z6Nb4gSkDsM7G4hq4ow0AdOkmoU1/3MXdgz2dVRlRcf+Katu0VKinSR3zFKNd/V3xsa6nIlmh1oZ
4IE1pae1TX+TcAg4EgGCUtPk0rEChj1AU57dWDpmJ3dmslwAIwDXqNXI2pllFirlN4sQJMKvSgTu
mN8FPsiFbt8GqVcrVDkePWUFyEmqDNK7oBXAp+c1E3AyBqqYMTOBPKNfaO55uXoHvM5+c4UXr1py
bdzv9SVo8Xd0KZfsIGlpwLy84L5yVxc/UzTJ1FiRIUvEFXbhLG8/gEliXua3SPXm/dvVivCH+r/i
p5fpMVGuvbVC8Y/Bpsf4udug9Dn+Lk+BSbHjrpjmUui3OpMX9a5SfIh2x+ly1jv9gxsyTD537gxB
4GC7Wy2Yt0RrLCszqCoIUqOWktwYVWdtmQK96Dhgl/1xfIHMN6v8urk1AK4d7u1QWDniQv24VTg3
4s8oOudoXjU3NF17qX/14hQuXLVNcLhvK2VwmEFrLzUH4IZH0s2dTMWFJNv2xBwrCQJbUnUZPd01
T4Dv1MzTA2Y5mtc0vKfop1PsB/4tlNfXCcqReuzL76Kb0rbiNNvPYKkKNMCPjyY0Hj6prNhIV6qy
OWFT3zYkpPZypbVDiRaoiW5oFLkYtGFfBbON8YhYv9SUvx1PoLpkcm6XmfJmxbrbUFHZk2TOGsxu
1vQr1Ziv28ONM4VVZebtVQOOaz5C2win2vdsopw5YF1X1wzoHUb1nKnZD4UBi4F/0corHLnHJUhF
EQuQDGG0P3dXp7jp0Uz7QatHGTrgPZmC1+cElWP+S7zHYSVTc23IHHWzkNzaGKcjvmHlELW6pWKS
sHhoFmCYj19LJBaPAy7U9AzjfePwkRqw5J3pPsGxn0qYYuyWicbt9njsBoPxzjhG/+UmSL8d+7DL
y9mGq0xAZdHd40Scl7b9jCAd+BNZC3CbBWPPYrPL4UY6iFOjHSUkO8ytdEiKTYq00luoLA1gSOdj
ro+J1MTQMC+imMIurp0dL6umsndn3+/Qg99euTgqitXrcvEKAfG6yTCSr4GhzZrdzEGtY0lj3Jhh
dfnLfUwedGFsaOW9RibkIe0n3hNxCH564Zueh64j1UQqh1CCRF1TzHnX3V6udZ4L0VU7Kd0KrHPi
dnd08/TigI6w3DOwNO+puY3B3xNqnG0RWgVPf1PQs16iDQPDvPNRXNTKooJ+5qbJTJ5oNEGrF0aw
c6e0db3t8XMG3/9q+U7Fj/ckDvMBOHeEONez4At6FuuNL+IqcfIQRsSf9ultkV3AAUz3/4i24jXg
tWns/9m18E+zJBCh3EqXh3wUISCVdsOZTvfeDQry4m/oRnd2/hwev9oZZpGXenCjn+yO/oJFpydl
FrA2ya5mlAyTbgT3G8LOB83vE4xyUVTSk21eLjVtDb/WwrrwV7dHUt1QZRyA8IAI179GSsvJPvzh
nPDKDWVnqbB62WvUaH8Dy2z/HZj1BQ0LzXIn/8KDQknZgYf/c0dcuRatyB/bZsGvLxXIbqUlzuqc
AFJpJX0SfgsM69QNLzZqCzTmpgGibooTkyHI+UZ/+8pvoO2JLHw+lUE15xqqqrV8pKJkQKiDxh3G
+YWuJYEJll+Tjpz8/WPYJ/Fz5tKlfzA+uO4g+uSCYCi2DvxLbRRfllw7xJWfY1P5WCBidNs6Tyt1
6YoRiXAnQwQiKhsz5komgSbpNMI9TOrmQTDzL3u2veMp9wramzuNyLfj0ihFMnYAAjddnIAYhMPZ
EQtGyAzknZYjoUAw9pLqJyAasP6fPzNDvB15PPRFBPRFFZrI+U9afYWrW7SnuxXM1JBkneWMHyAF
zHhLUFighCKB39RE5LkFFdzHal+bA97MVMEJ1FMdGrFkO1o6Xxx+7/zzORUkfkuPzgfT1LZsQek8
kBFu2wAZ6PdCUcEifV6o0P8294JvRjYCLWgB89C27ZseZipA3R6/IAW7X1k4+JlKWKO+nZbVVz6E
E6C6nEvJ3eJZUaIA7r488lm9GZmSv1Q7RNOx+NJCeicu2wlZEM/HU5E9LSBsPmEPF3Y8dAZaHxxO
iJNNScXivGYC0gRVvEg/GM4HP7/L7wzWMGeqRUgYNN7oCrt0TuelPyC8e53O7Ijre6HcKWAdA+Iq
ULlMx0WE1cD3eFVPXtt//mYaAfFINYcMjrNAoGcG/sty5BIKMTLwWwVUl0s6MCJejWucMnzCut0q
JnInzNUymR/ZaJT0wvZMtO5b9iV1MUXmNZaK/W+dOhJRhEL8EpniW6S60x7gi/j05LdDuU161zfQ
FQ0T8jUUef3fH5aK4oGEc3XQkQdYE5NHKou1pXjKDikHZ/PajD557fs/dSQPEa5GNyEX+bs3QJyF
MHKn/f55eQ0X2UPvncozb7yNYP191vTXmJPuuwd7cr9Umbr8DP5MG//MftzBTDKOP7EUiWGGP2IZ
JjFOKlG76afuwlrsX5GhyHgTazaw0M9cY1plea+87CSQRgF5lqCNIBfar7PyFrRMtLzKWimFbjQd
j+b1Eb5xi1leTGNaI3oDz7IiMsYF39rsIrScj9HmHZ0dQO7TxMq/OVgrB6klBUWLnact6gvNW/n/
goST52giNp3tEfLyhxZiATysxG+G0LBE4XaIbGQT6EFefWYGYY3NMT8gU3+qklTS2HWbFrXSGF39
8olZeHIlatJdo1+Ar6iX3Pv3l259OKOnzxnX2fx3xeIrWtyqPMr0EzQo9kEmRGJ4xP5gxD8mXocC
wxk9lH65cQV8PWRlaKnjqKiryjQ6Yem8q4sUk8OSsJo6AlYhIrjB0qONoy7b5ON5CAleq8/ADXXG
p7uuJ5reRAPufpeTNM+lKk0/PSoxW/lxQadr2wOa2YNZSV8QJcIr3rnYPV/PwS/vlTkQ0oByWhgZ
soxyDqwD7heNNxOkgpVyr2AcGXN1BccD5w58qY0Zm1QYE+JndDJAOQx70Gav/g44k3P/k645LuXq
BZRm3jV9N9qkehPEaw9KObiZP6ExgaToGwVtfFhfEEqxJ/GdyL5zqPQZu8UeJ5YkASGjR99v2vm0
uYxVqNBpWwoFMp1VC4ibDQoIbrmFcRNL0v28eutO0qDWZKlVz4bRJAS+yzq4k8D3UQiLYClB2YRJ
Ou0X8zKgoEe+sx86cXGrLbmHgGUotE8wXNk6emT9FVURkbg//vdE8+cffhvaK+khH8o5hfDxRhPw
xo+GIo8VB3inHtF5i81TtXGik3F914BJEngyNdX3T2k/pCTrpjbhiezRyEOJGuyvLfCeDPtytzvb
Fscrg6TeaVwqog8C+MCLWPY3IBt5/f7B/xkqUDvJXNYSyyB6VS9YziXnvtt/udUxNQ6Chyl8EoeB
nGR55vNRbBBhLqX7z84aVbFfZ0/I02/PZl8eyxe+keD5enGOmCfqho0vMXgDnl0mq9O9PdQ4Ap8b
Y5AjJeLptOIdY8G5GwhaI0LItQcqW5nJIc9avbI2VV1LuQKGCQvO8VQQSlG9pPTjBdoceAsBM9Dh
VmNnoa2Dk40TSaXi5fsfV5lPcpeFMKF02or64OmwNg4HYAwQxbU5dk6r2dlnlAFhdZAH4KSg8tkz
2QM/p59stZ3WR4XjxQNlI45KP9y+g4VpPPy7AgtZvQWZZaCcGoBcubKNkuOEvTC2gnQbnkiRu0Jw
6iAHPeiKbBpdPCxFjxMXz8aqjvX9R1ZG3gHOCuJiTZApdzQ9sgDMe2gwgiqnBTz+wYE9CO7MlfuY
jb5YKJ8M9aRTH4X+opTniBv4DiLp31lulxU3OMXC9wrn+U4CfjkuZHlM5fM3MKbic775NWrORhdK
/rYBQ8qvAW0j2wOfVvklrR4iPKy8LNuS9soEh+A8vdRwUoiXVfDcT728TLm6au3+SV39aYpMKcy3
fh9kazZvRiRxa67bensjCAHpa/qbfHV6SlYWomTQSq73XuEDW0UPXZN6hBkkc0T9is6QmlHSxQjl
irEYTDhzENWZH/42Er4hcw5Ckb1dPFPm+2QSTFWMSW4t0g8HdspW9emD7A/6xLOKsHnOK/jvewBG
XzkbPYiNIq+NLT9LPzMkBXkt6e+w+EN07R1no8HFipsFRpEwN8D00Qn5EzJpazUUdQ4A4V3BpOI9
2e3b6jaWYWz5kw000l72ZaD/Lqso7GkmwAc7nWZ45Yb4SBOef4Eo6yPCjfFX8oc2nnqywgyvLN6f
MXvahrptQNpunWGnD+Q928W7WVF+tlzvS3avO8+chK3pLlkGo1fizZKVL/UPlj2cxVjO6pLOLOK0
xGcZZ2Rm5RfbOtR/QVmk88ityMAR/g2tvsTFbbd/HA8r+A7oER2Drwi8nVLBOdNbqf/N1I3EGE9M
6LuFzHIEIay9I2chxQMXWLC5L3jVzYRIOa70LpI7bXM2bvILXSO3VlxUmj+CuyGPDm5SCrCtwnbC
7SMmv9rqOFo6OWOuKudvIWn+DsDMjCRLGY8TDtIstl4q0s/OFEwmUe/zONrHO4IRvys9WiQEiax7
/jSyDbbq5JeEx0aM+3N0Aa7WPjr+N3qp9Ag41CQQDkyn5yZDlqTpuQGeoQ9ktO61ap+Uw9m0tA7R
K1Snv0xQD2WO8i1LERMS9c8IhVXgNNdjYl88f/l6D/Zn7q5lUj/DNja7E5rAI67SGltcHLDpCa+p
darz5Z+Ll9mLssWy7x5nVwJtnYcr+MX2ygYEOhAhMLRdKADrZahJG9iF/bYReIiTb2XkQAVxnGIw
GQ5mAwLV8Ckwo6WmfDs6euhDV4uugj6gbkzXeSuA+J1AdREF/tfxcJwPfBdN/jxMAd0KEYWg9+pV
Ii0GYS9ZuiriubcZKHizbVfrxKnfz9emsPykEzdSA5/Q/FiABB2FpszU24HJadOGmOMVkLxKzuJY
IY0t0/sj0ZlOH7SF2MHwwxYDd6XCdnS90GeKzShRAAmBpsbGsKmDfdsfs3vwvU5Q6qpDB2tByPYN
qcokLZBCimAnHuLQO75sDow8MX7twndd6GoYXv8f8HpK4a56q02Rg29pQCQAcLU5U9tHmv6FKCZ+
7gtpqK0nljbb9XJDQzXOS4x+jYLxyuLXtCda5YApztuWe980QjENoRz9dUEfClSc36YhMDYwBMCv
dA0sTLp97ToIEVRSI6SFK+gs7H/lpKA6LG+CKVU51pJRd5d2tnBK5g89iJezIFdDSIm4a9K0ATI4
C8FzTR3Pp1t3M10lgbRayGYyeN5f78Y1VlIImofHcOwN4coJ2BYN+WdNiW17WtE4vapmBws2UgnY
YFbp+m2haeAiuzeD9b67ac++Jsd6XkKf4RcBoR9HW9nyz3CsGmwf1akjNgsqsEqcJ/M0Faf/eheJ
SKSxz4WXy2bVmV6rZawoPpTduaj/NQrh3khd7XA7tyadfnXpJec/7BLbUbxwAgqSlNezt+sVgOcP
alB8ugI/RM+1h51xQMIcJWdWXAyUQ0/juRp5XAo3g7FipkKy09Q4knAH6F5+ZrJFoRTWe4gg9Qic
vtaFFSe3h0B7txS8j8B0ksi7IvXU7hjWjDIgm6r3+O+a2sHuCNQ3u5FREaRF62E4xsV74jPsHq9g
eq02GeTOVRjcvIUhJG6KxWut1NBXmrMvQ9IaaxpXiaGf7QeXxvN6b40960vcBNXW9RLnl+oTEC1c
QNXj6bijUpvUhDMhp7BrcawiHq8CeiVyJvG5FiOSyqvJzcF7Dy3RSUwxpTJRLaIkcUa5DrR+djDL
5nq/vK9+t+4pUUj8s3W6uUbf++N+Cw9RqCdXlZmiH6Nmj6JzfXRSjMB86obDnL0EoxHwwpd9Txka
IY4GXPPAmPu2Yrem/oxMXFTCr6Uq3JxlV+lEH141rZaMC4N8zcmjYjHPGhFvHq5cjEOL+Ma+G2B/
XZyvulXf0t/zQlrQdRUwiG9PAfQZjLWbltqNKyuMZKQ4GHZYp3H9B0l+0w/96Y8n8+Mc+BurPos5
JrjlukTRkF3xDSzQFWkPdOUsU2/rNtavEvH+ybOBcKKCWeT3WE5FVTe3TA2eq7i9Z67q3exMUb0Y
x8Xvt2dVxVJngXT6EeA/FDyhcAPJChfumzFOTLA3A1JZGbz3s09eT/KnXenFR60IxBz/C3mBh3vx
I1Equjm4Q2ZSd4kds7FfNXP+OtOYi0XLbIm+J5eSUtIrN9KYtHTMCvR/1u1+QoWEVnvegf7ActBl
uCOlW8wf0LwAV+O6I+dSIF5m12hsiX4vEeLKriux9I3quDPnjVa4JZZ2mjfxN+32LfgTFaeimT1D
xWSFT4lz8DPzOwLOVTxuT6YVnSlyoDbjHy0X0EMR3zfDISYq29v/zuqilgnETbVuYKDhrmc8ulUW
gApyIUR86ButXFSDgNnAr5aqRoZ5zh1w35WOv7Xf9P7akC/MiXRXhjatOrM/PImvGSLJ/s+7kcyp
w1QLezDYmWcaDsXbzN1aK5hXg17PF+VIUM8E+Gj315NsNpJ0NE7gcEtTr9zZ4foWJbIpRO8YsVyG
UKXE+EyLQkLaymogkAmDdZK0Ghen4r2Da3G7qYXc6e6YHkxgp0zHL2KU4mkHIFnbvvtI7sa0bZCL
wCjWvKMdzpo/N3YgANSp7IYiddN/irbzC4OnUbTFxgRDY1EXfM3F7g4FjNGQDmfgvyzjsbVCKAjO
OkrCDXrq7KMGlnckIb7FQVcyb9fEHMU06pd6rBDOKO9uSSje1GxVG48Yass9eBic2ADkplFA/RDw
653jnXs2ftC3phTF/UkItwOo2LAAU7COMHgipncIrRAVjH1InxZckitZJ+gs0CydAh66V/jinQyZ
Qol3rDtk1Hun+k9n/1u17rk9JMGZBIL8QLzC6BozbU2rsWBas1YC3tsqz3bjIfP6AfKInL7dr/Da
GofH1kvOEdpB775FI5MBlKAB73Z6wDbgu9fJ4B5wfr2OKCGfdqQFuMI9uc1s30Js1n75+pVEs1Zv
TCPtu+4eW6OlU7UZ8KSU01c5ntIy+WZygXcTpEOMip6up4RgmoV1oKm26AN4+5Plo7fXneizgHNC
YUjDtsk/xCFJyQrOTeQAnH2KiCF3npCH5et7zyvjrT0XjGZp+7kY/+hWbqyxI0bEpWmud2lFwHir
1xPuZ811n1hGyb9wxVx54ERQFeiC9/PWo5O1diYBUdKehltqb5nuZsro3cBDwyOBt8eCruSTuEec
8OgC7hqXMJedelHC6XU2uu6rB4u0z1RMtd2pAbwWwsudDvbfH6o8QG0jKqoPKikW105QzUJ+evQM
TyZx2q8qBoIRsipmOJum851jm7IAaVVDnOwqnFwsJzcE8YwxSSqZxP+riyspwyTSWuhLB03OTYeU
QJgHERfPlO7ghNYy6EBwseUJX71qyz4EfQj+SfNuYDLHebjCZpt0HCnVyoZRPNrT0ZyKQS1cf4HY
erbccYsogsBJ/PaleuB3Q5niuJRjab0sSpOK0EqHnEwhp+gPuGBxlJlMXU/1uwpvpSWrWoQNXSAs
eB8Y9BZgHJfl2se0pudTb/isoZTe8KM/YYSs9OoO2qILqXK/K7D+iOTnpcjjNOcYy7NrN8DCmG5O
Roy/eQXzQp5oFEifVZbHhQNRZdu5LFZefwHlEM32OA+09X5pfi5pAy/48kpHZGSmAmD5AK6+jNGD
Dmvx1QFm7nZP5qz1vClyZHERACdmCl+aIloHFzXa82orjlPjPK2fiA/Wf0N/dpw9JooY3PWy/jHN
wS2ZmmA0eHDwrtzqGtTmFZgBrz8CnmSwPGYTTsvgzJA+Rhq5vBXfTp1oFsHZtWNzg9vRj0waOuNb
6lOGcqMhgwciKeQiyNhCvO3hpbOdt+45ipzB6gjgxe4kEBWThXz31ozdrJ6yKZiyrjg/jOLD5ja6
iGTs2awpofsDuQy46amnguEpWje4rYnhrcatQsw7kzRmQAZO28sQHOZHfSbRqY5sJOD/nO/djjHu
xZmNoSPemwBFayEYU8f+r/JOstWfB9VUjZc/BVi/AuOIKVt7HBoLcxTLuoJg4eBkwE0JdgnPpd85
CdJOGijLoIEJrULB7SKrOTjCJfaufItE3c/dwfTIS0HTnVo+lOlTJAAiL7sej1LWyq3q8I8gqNEp
IbxWGjk3VOIu3WYyMjbW4zSfLoqihoQrua5e3ffHxtOplvWlwuKugxuUbs/1b9vrMwkR45goXX0T
NNcp/v3a06aDqUNO8DlHYyAjUSpip72MTdW5jtydjrYWHzfcAvGunA3QiTDG2dAEoIefATBV4mkZ
cCWBqZxVxc7gL96kxPoRBePYtr9oHLzKMxD6GVAzDMgI8apiGwYxu+H6HNhhpAVD/C/Zms8PSZSf
FD1cvZPy8OS+e8d0jamC46IUmWl+acHblXTub+pog8JjS9NdVb34++WGpOfFvdhYvSfTk53Sj8wg
airzJDka2il3M3NsfEb0gLRKIgRk3aq8XZsa86A1gq9XHGFna4BcL8bYMApCYhAy62YM9K7MmtWg
di+MswaVAijwqUghIHyXg8rTs8LKpNygAI4suqLw5zZs6rSFpufhDPWVNFRHCR0ZPMY2upiTwD3U
CsQs2vyQVS6Y8yga4keJ2xtWPaw9BMQCqvafIKumWcFJ4Rm4cv5ROJt/EzomukqJu/JQaNZG3k/S
nWkBxb3wme8bZXm8ZZyD3JWe9tRPZQaY+HiI2duvGRh/Ei+zVIqcuatpsout9hJtP2rruvbxn5sS
PTZL7oudoDSvVaJfbjVehaFDcd8qpabt52mYAfp3s6a3+J2X1is2rAM8cr+2VG5eG+IMbYMb4yYu
41L10iXv2zULIcyKKLfFGFzCj0bOxB9QACBUxR6loJLFzjK49b6emEfISGfJuQvlFJmCmuWrY7pF
mr2XTJbbzeSjXuxqp/pdZysl2VRGMTTOkvw7IhE9sniI/xQuWhN69A3O7/RgGi79e3SIZciQONYo
fIIC3O6DdP2dBDhtnOJECupFY2SzJBm9BhAKvtWjjCAWW1EAHsd44oi+3lL9BdLQRGS89OtLTMin
oe7r/OsRa17mS//aKyeW5XvCLrguUGihc0yGb4KMV0jWRSWyezDSoW+2RzUznHcib3VmVRPWTgLP
7acILsRhehYlxRVmRiNdoiWSOojzq+qD6Ukv45v9udp+xejiATY6CHk0iIcsJ80STmiRWbwkrBNM
dGpvGhh9ItOTd+yh+oSMY0ayYkkRFJwHe/6sU738GqX8iVr1J+9sshhDl8Bdp8xN4ulU6WxOrHBT
RlpHD9j97XfhIF8QvIoSCTEvjsk6zoB+ilK5yVOTM6Qq5V/Rs/0+cLh8rPoQ4M4WtfJOhSYcUtVC
yDI6R9k95wI+9ehcaOp0aYu8cmlO8cZ8pj/MgdREBH9hqAMn2OcJ1KtnoN5n5gyCfJwWMbUKh6v0
0kK016Tbv66Fh3V0Z2Sf38MonyTwgiqp499EaGJq4MtkS1vMo943xsymhtn+MVsw8weAyugH8+bv
JUcA/g2BNdXy82pO/2p3IncqByrtPrvvvYey99fyPbssXuAToC0ZS5VxnUZhjzmOv68wlkp3CnRJ
PXRlvpNWdAum9eNzK0GNrOMWt0+EyUGmcdYyJmIWjhOE7LIJgKvkJtsuyUtAUIdfz6PCcmtKaBCb
dWyk6iRQMhhUsK0uiiYKYt3/5FQ1uSdMpVblCmb5ZcxRYsWkbR9z0EW97SPxOU2kxrqhaZJltLr5
Xr47ke6vykz2jVGxWnOAND8/1rzdRKuW5ko8D8UDBAurJjx1irD+4Wx2itoJiJgBq6B4OTNk6jVb
Jbs92hnTxJi7HR3nKkuVJvruqCxUqRpUv1/Odeo+Aqr+bM4a+Y7MvcwcUZgaj/YNxux8j62rbTen
PntX67QE6Qv00R0KwHEqyqF5k9fx6iM8GXwz2on9gQxiUmI7g60e7hBCGyoKKdIAtVx2NueD3vDO
QVKMDLWLB0aKwO4LyaP5tiu0mldQtITZkt//Mrxkc5SAEiHIf1gGJ7lrhpqyW1fPsrch1mD7cC4f
BtVBbHawj8PTItjxZ3Cq74oQaoM5gQjL7QJOWZNHz3Et3fONtQajliMt0C/+IYUQ4Ad/Q92/cLd1
pdVaR9lcgUpJGza1xzRhVJhiAxWxLyD7lyGQ0obKhnlGYN/ZIF2IiQnj5kmOGCoiAbwVmHQYq99Y
vteIoJv1GRqEw3ZhgN2nrV6RVh8OxOJxR56CGKYMQrtNiN6mUH6PgR61XT31fO+yJRzhVBOjTztk
t04WVhwxjjaZ4zvHegw4j9dfjWrlTYpi87NLinvYPSF8Gic53Dk/jfadmpxI+kXHEFmQ0UdR3ySG
NNU2wXA56xy7qydbYR/FpJtJhSP/3eUmA8eNK6x6jQN8hcGOmVmTkBeHnql7leWHFQNeMgUIJJh9
V+HmBLubkjv8Mq5rNN4Nl1AQdqEEL8cX0nC/m0Un62Q5GUeoEPjN3hdFA0rRiiI/Kfq5jG/wTIQR
EqOutKzSEHzw2HSVGvdaKMMpSWsXF9/LD1LV1MkNVQZ8T77OITsXDvpPv94/tz21pO7VlnRJ7sDf
CwNdTAKrZ9q7Wg/YqHxYh6lBnDZVSEDddq4WL0fskX42DB7AKwpYMzixKcy9IRLCZgRtoQw5fk7W
iS/cTKYproffctkjsQdP+35FeCAy4kVGAjAwdZHMsUvq4iCyspJGqW3nqII2w+UAuz5/0QoyALqx
iIZbdizCabtcgWSE/sl+3WQ8UK5KR2OBvpImMarNkRkZUu/nYlozb1ghuPFYOikvhEvvzuP+/M03
FnJe6I5QKZAJOiYz3Q9sxJENdzk5DFH/2ia1ifUn0N+VdSN8CqH0EJuN32ZjCYPz4Tkly6vowpkB
khBXDYQqn8KDKWDpGveHaNIUh+nAc12942A/31ulFopZnST8blriplEV6EU9vrOUG88k072Jaswk
AsIbnhFVdPBXAzrna7UFxm17zCBwIoyEug4DkE7K+DdV3K06OqMaW9+KKlH0T6vc4YuaX+c/o5ju
n+IQPYvl+jX/dpg6yskR5B5XFjJTyFYQBdsNWWRusKTz57UNaNcHXZVVDSces5E25zOg5oXMYsBw
nw0jUgJsH8JOgIL4UOGmpfowhcNLJxMj6/Ce9/Hw27VzLD9SEeVSB0yl16a5wCXuhlTFPcXvwtnC
0sa7aOBoBRJRF+JNFcGw8uf1ySVPfzyueoSqhiQX1tY/vjTQn/Lfv3R8wT97jRJzlNgLDs+lTDX6
EkUe3QemdrBm15VUCTIizcEnfgSwoX10DmOPnsYU9TxunUzpvU7/fGhoSRLzwIiLtD+UollG0+RG
BpKuqAPwejVKmAh89VWWldkCbFEPyEbMjgY3Nv5EOXyIcxx89HP8puKVWjHVmqsaLCMyC6sxGHcw
DXw7cSRBha8lDHHdGCYOEmbrhqIXHW0EUvTpZ+fSoF7Rr0OBO3/tipG6pHwGZ7rE6Bq6PA6GhyJ9
OwrMQ9ab2cKebNbfHakF9QqxVl7WHRb7QWb5PtRdFKYpatO/1Z28EY1RW2VjQf5m+dBXly5FUiFt
yqZLsqI9j2j/6lTq4zU4O3GdG3Wpu13c8XTWuSgAcKB9w50Jf2tUaUoTYOvZswt/0jhlIy90NU9M
dWddzbEufi61UuQgRWWX5xlW52nO1eabO8yN/zrt9v1brtouMmFuwfOC+EFJo9NBntzRl4G2OoDu
Xo500KTbd6ckoLTbXN9fFv7Azo/8j/uh3MM4bP60Gf7/GWKkt97TlS7Jr1jtKtoa6iaOlPYgxCnM
hgj9s7JIg0B87HOaItBxp+Pf3JR1gKobjGQlMGhAZvxhD3kyroc2LNT5HtOc0NfL9AQmz8KCynFn
gB7MQ4L+t03Ype3ercZtJL5TjqcmpC+5BIFc9rbG2Hm100hk/DgUPpn6taPKkD+6NRYMlciDOkSJ
8mBbVQyncWl/7rp5uwZBCFAhdXjABT5GeB6xfX6+uhiIi4/WaE3YGdKfGPUMrgZNFzh/8bSyWJFa
Qbr9HkHr918Cp6KZBbGmmyhAuErb/hX+GyudQWUxf5dmmL/+0ghPo2aTVr40CC++3wxv9OF6qSfx
7KtIaP99JhWpz/1en4mRag4u1D9xdDOvxThE7UY5FKJn9z0akeuZ8Vhn6ykOpeE38vPApR9/1uuX
JY2ssdXW97gcfWmjm0x5e7m1ny6IwPVx6uBviswbZuz3XHIk0dfb+S0nMsWHONnQBDUELn8gocjD
w2lVAhp4h+NYZcLMOmaM7X31/t7S8t/htqU0lbWErKP3Pvtobd21/jezlYjntyGNMArc55dBSgqr
DD1FfKTghI5LUIcikVjo+9m2hO4WWquS+huECHfRuxpC9wUQ+0WcMRjcloe09KIcqCoi/vjNpb+T
w5WWkptMxnqOjHOlGZzhU2JwbaFhCAORQ0pBdrUeEBqaHutJcyBwIVUIETwcKiFt5IibtLPzWbmc
4liGTG8bOA0UlJDcOAAGHtsIlXfX+PWrx7kTDeOXi5RItz5RiVev0vjkuVrWPNYG7mmhdglLHYvZ
VyKALKm4ChYkM5uXvh/QrgQewUM7pLsGjiu1zz+IYRKOa727UXKCBW+EHqyMwRyKVKUmmtV5Jb04
jBTygp6PbDwPzvmtbW7Z9t8KrhJZaiIZqUjfqoN8cokE3UfRTD/40YWhxC9Ul8TQoTH4Y+5WQuYc
f6LTEnjMQUJuLZVkSYUPZVAwmH9Gvs19LUhSJA4WJyFCZpzw7PIPTyroQjZR7fqbDyB2D7ZKwwaD
LT2b1KVdOwQYCRBRNbjkOx61Z2HaN5J02s+8pUQ4mLechr8VfH3UN1ZItevfRSMyDO5YfuD4kSyY
1GNieY6pckEwv8WZB1ATGSmQj6elIG85VaiUURwaBjN5D387jjs6aouVhJd6vqPOO5xl/WLMAXKm
VE5hOblGG77kcn1RSyUn1kNvhby9oUcJ7IAFbNcMI09otlO4TiMVY31sLp71fJO6gzO4w9La74Vy
LkGXSEpCXZbIAz0bsFyBAYEYq4NastfWpIXQjGNup7g9glvHoDBiSGioWHKKuFAnks3lT2gPIFLx
dLngGm9/NnHQZjChumFbqXl6Qg9qURVYxb7m+NNKlvkpUaej3ll9TSwCN0Kw+HXn3tUvB7MOyyZP
G6Z5aGlU/HgX04Biucmlj9RXzm7ENhG1dnVIznk9fRqRY7dldmKwQWH84bajAdTB9eLGInyopkfS
kjiZNgHI+g8VNJpyaezO0pKrpds+LGgj9GRZtSB2uxJVxUxp8e/k7pDwIsyF6SAmPF97Sca6oKeS
gIi005HC/5nLelUUPJ4Q8iUzivaAbFEvJbx7JrMosTmJ6mtwV1Q6NQj7/YWOHffunAwXPp6ONcyS
Tpeasimo1OkOHqB0e2c1B/oAjGXFKK9doy2pviMc736l1HcHH8QffR/cvglumB/bxnplJMPZUexV
jgTepFFc1Idjnj6jnJ5cDWYxxUYMgY5P7d+egdgyevS3S3I4bNONy3Q4cB5zQA03+XvP1LtVsesG
Uxr0XaZhYCRs0TxjhEUNxg6QB2Fm5XYY7VUAEzQEy5abNPxTAeAitOoUQnglMAHRLVXi5rKBPsAZ
tlSxfH2hE5c56I+nffTqXZmvnEHCuF2Idt1jaxvW45hLnCtePhU2swfH0mZJvDd5woI64BGI9hYO
44pTZhqDndE7yXLM7x/8IKCFsKCh+IRcNoFI6FO+QF581hrcHq5Gar9xJhRTmjsm1MI4o/fZORk/
FNQQJhzbTnVPKJ88DAuxl5baZWQ0WYlbkFsPMkBMGZD73LFoBTwOZ5PRge1IPHCg+Df4XEnJsu/Y
ibu6FUm8JJSYEDpC78AVipsNvU4EUGsgS79MwgHZJyxUL1FikuojkjmrzSvZxJ2ZrThIwUme2MOP
0dBZJT3X5EP3hFbGBN/7U6f1hnccF08hH1hppZFYJOPi3uM16TnZhpAFk64x/wKkXXq22fyNERIY
4egN2Ci7oBbJuyaEm+Qc08OoQAyCeP8ifmHnaHo+StABROQcWZ3JglWN7+43tWuKIsiAVfVGun3f
T7os4hbLbRAHrisGv3dB0E8uZf0aF9SiNL6xSJIdGCig+8/nD8wPJwgKb0qtlv6658iai509nyjT
5RFnRxvpQm8U54S2olde+M4/qE84xoCvyMEv48/SHjvL3JBpsi3iDQOxBN7R3tgXirQG+WIMWbBd
Xwd8ux7Ty/zybAJg2WP3De1pCYEFkFUQWQUckUNEIiXvu3jvdlfOnykqMe7kH+qFfNJc6baBidfP
Gl/hbT0BJk8fWhYYt1oO+bGhsO5zwnWmdPc7zCYhQW9tSwYu/xYnnEHACM2qjPVsitt/F6K5KlFO
aff2tLg0lC514txCPiDceXnn/hbswmld3yfEW1YRYlnP84up1oUZCsHc38cyJUIZA/vf10as1i1H
oQVdJCLyH0EIM3GSyX6bAKWqh19sCv7l0MSKH74NcZxqiBUpu0xW9i5P7521giz+gQkUhYHe43J+
Yr4pu/GrYXZZeO+kmLSRlDAZIuDDmvJv6tAwQs/X9OkJP7bn47T8iXNAlz+YKFwVzmBapHKHV0M3
3jv6/U2oQAZgnyLobv9TaKogtL+lSfTPF1fU0FK+18AGVJO73/aqYtt35Q3VUXdX51CsI6Ks5tc2
9N5YpakmI+G+vmu9BmMFqg5EDs/43axio2PC6ZOvkfnNAeYffE1kT0+GYgBz2JuzhQbDaMrduXkn
abMX94HNW6He6TtS5yMV5q2k/uHpUwZcB7wTuzK71u2mlFrtD0g9vlrxOogWpmFjCsnOcgzVY7bu
r9/iEcje0fGdH+mzX5bV0UM32bSGmMaOgV2YqlNNdQwhqF/ppxlgIzMHtCdKeW/RWl0e5LUoD8Wq
wmEQodhGE+cr/lL8r9PkOOXhVUJAGv2tej3mkBPtmHQHOUD7q1sfwJLhnRaJdsVNZUJRlA0CIM7z
k+UYVrOBOKt82YycPChwtHOKTjGzB27MzWChq8zeBOoliwi9jxRpjFYp3P4h5a8b6vGlip9IVLM8
9KmwJT0ISw1DfDnnO5cXLzD/+dOp04osQRDkFkIY6QS9Ca90IjPVGuRgJRjF499sGGjfxlO+HF2p
Sta/5XKWjgKK0g6vIHg2I5RaWB3sY9fGrdXnpNEfGOqcNx+a+pwhuq15oHc9MsEy30syaR9InMqj
Jb3r8C0Jzi8XB42tOJ+IUyUZNlwXNnT4laoSloZ97qEDzOjKp676Br4ok5520lUqTnPPyVtvll2u
IIV0fiZn6GNvHPIpTZ13a40kYrwyqA8FJvbBLHVB3C4rKWCqLFPxeuCzSNUYZs46yOC3iaZ9DMxg
KQwkMWTc5RgzNDHE9QqJu4IOHCEbOoxk51d+1rOg6Y1N4WikiMOuUBjtrRWEdQIYQqruz68h/5e+
R0qWOCXlV3Rs0c04UvmA0zvZJHHi4iVhoTSH/Q0NyW1wLBpLPIcuqo5YAjntNrBarFJJp7oGsRDn
mwPizhXuwkOtk58uQajggnbbJLXTIAvv10oIVoHOC78zjfgnzEkZAkEmymr1/XEVMPETGFxDEXDF
/7F+/pIMQq6R9tMcPhSTvJZkooia5KhujTfBGgGqytuUacDSQ0XBT/M4dyE7YVt8S3o1ER3k5CMa
dwQHZ1b0SkRbCxj/UIiMqiXuTE35hdAnU9a2Vm/yBnqxsD1y7uHF8y/JrbDt+31gbNjQB40KeyBb
hQx8Dtrj3Akf16Obqv0wdyHbgrom/68QE0phNystHpkbDIuMDLGr2OUZ69QstmWIyUc32QIAbIPu
D+Kee3r0R0XZNCnwkRcs5IBUNH9ht+2dYhG4UtkR4NvHIqBB37MXdzOwNszbLeYIzUbHNTXdGPP3
NO5x8kZxTCJfAW1EGP6SZMQyYn0BRSIycCroTiAGnNTNp9++M2Bh6cf5yYJg8TLl0pdnNT8HH4Di
3kibMJLFCQTbCbzG5k+c8oE1Kz/JxCw7qJevp/81xcpQnA8bAWzG6v/u1BpOd6TLKx7zxgu6gMXW
4g8aUp3InwT6s9QQ092O7srNe9cgG0uV7BgcZX29dnv5OBKEUbhZYRi4XW4IHpRSlm2AE3yDcQX0
DO05Jj99CYrptqioAmuP5r6njKR0E/MveUZhM7OSufxY+pEcI21q10L6WBGZY9FiQUyYZbYNtTln
tJAu15Eizgnvs/Bscx/rcOM9X1hHy/YQWFNKjn52ne9x/jL1RonYLrG/MYvRougm+wvV5GxkCx5w
AtAmRXJdfJKbLuWAtMLOi3PiegvCWI9weUgb2LMadRye2B/A964ekBWiFdEK4AOBPDSNhSFuZSyB
g7N5F6ejuPHrz036IcsVzKLHJzGxL/6HJjVHYB/cQPUX7P6IUNeeC6buK+EC1xVrYaYgBXUcdBm+
rJNuhYaT18UjvfPZvcmTmdCbt/tKqRhzc3xapPN98y7NLpdhdNTo7mgPmqGll1ZP5S2ZCqLWnZKC
JcY8Sc290+L1TGjDxsWCNbyLbltKGb+pbAMAc2CnBxV9zfS6fokzxxRaHMKYU3jALpIYh5lwIYij
dYVnx0HIS9WF8zp/n54GxxKpxKGJAfPstdZkX9VK3xDF2JqQOCwxu82xOS20HsYT/Bmnkc+KjQV1
bnaaViLv8FIqHSJdZs31+H5gsRlJqgvSetxZ5YOQFGdb+GHJVm2rm7D1gpr0YlbzulsoC6ihicQ+
NpOEz5JrTediIAEb4BRSVTBL7fXrU2GULy1EDqBc1Wn3jco+8RFKNuwG7JHg7cok5fqCcdb1q9UU
dbTRrVy7V6YOLiRKNBbU21A7MNSXctpoZ3eHqzYARt1Tv9KylvUb4qHkb6B2xwswsLo0TGQKRzk1
WpPk3Saahe6apyffrfY8GiNl2UB5I9xbekPDMdK8RsT3kqUjr+4W5Qc+UIC0ZgHR0EKNaZU/vvpO
IfhuvxOZU2CQolwnlr/wIIXCLjTE/N8wx/Psgib0iv+YW+xEtRiBNokT/YIznBxeBYMbAksuT589
uXe+RdDQ5BeDpTD8h55GppXZR5m2PpcC1S208kNl0vinvFRlvF4IkC3BoLzwCqmapXlmkqZaRwk7
GXJgo/4PIVXSUMT7RiFgAryuyuVdseeCZZtOGxbyzjrV2Zap1p7I5i9WdyOrqEy+fMROyZREu9xu
1mWhY4HbRpykHrpAKjGyfiIIbn0NB+COXRanHcc/tPJz5kXYvbdBNxW9m+NY2tkW9MFnfrIanV5P
DIvAzGxrhQNWQxKbiW17AyvJfwrpYUN5THi7Hkb1cUr6sZM0BsExjMIaaeLy6zbWUqIh/iJdm8hP
OhZSCeFtWL3P7DXWXgpc051zwxQjlI/vN50zy3jk7GfP/qsov4qpw+uGvByTaiDsw3vJqEryKAeD
cHYqGBJSdrvpiGlDh2fKY5tvcO5h6kuP4iJbW/XlppqYqxhTApAexVWcYx2rthSWjFBR7YV0zWks
2XDKrIWK2uBQrR9YIdV+GDjYKyj33MHa/YLXzmk2e6LLEu0ZRmhiXpowiu6268JPSi7SN1QTpKrL
Z5aPprb2A5GAXrSzAj6dx7tuUeUbzo8sYWvHeRXDhNZoprk/pQPdPq3ZCGqXk5e7FSezyHwJ+SYZ
eHeWEX/wOonlYCXs97k9g3YSa1Jhb5PFH0yaZcXRb++bvEs8IXtkdZnp2gzhtwm969MNO7P7I58D
2NJypC64mY6inT5sg/gDQXBLE2B7Ckk3crCPVvWqq5keuNZvJapYpLM0SFrTrOFkNYitcDnTtVGE
PfngYXYFR3VnAAukM4kneTLl8k8O5BybobOlB9bb8CunVg2XdNGiv+uA0DBxE/ysTBmorEzOUGiz
tB41Ca+om/k4JSCOIUSYZuge+JzB4v/MmkeQFoZfIU1WbdNXW2GBzDO4+mEuxKEq78vN4L2Q3Bw6
42zFujWnaQzSQAntC9hNQUQBdNS/A1L3VNQmaMQXpxIa3uAz6ckorPN9EwKdAdSBAS3ehWC5fjHE
IgmnYj06PrmTK4MAGLsCVV8H6QNnon9pQf3IGWjePQpnc80CS5o9W/4gIX1OYZm7EYZdPjXpPw2a
4IjDDk7v3gdZlX2ktx3B57eMU3fMWsQ9HB1JFNmoQ/36qoVlq2a9TR+6k31nHVKTn3ymUuCjJxyE
/ACfnb4mjgVwuFBBegqsmBqqSLdUWy2piSuhWh5wSB4Semp3xahIQGZJNmdFAfy73HzXqw4gyuU/
iEq2Th3P2/mSFphAtErUnVH0Ldv+zSOs+cVp9jN0OhxgbIydnp8eiDTROHhOUq7liwNfF5+AA7ch
iRZBEh+JTeoHmH3cr4pDdM5KScMnQWlgf4J/TSq0I5TDtITz/7dJBeDTqbpZ88P5XO/CRgwjHtfb
qKnjb93o1LA261x9M15mCNpw2SfeoL6rBSIwTkW2CdeYLwsLxFyT9hzhSZwJvogtjTfdG2dGVMNS
6XuKRwV8FNOCsuc0ceyXOrtHIRdtzYu6k4hID/5e5kakxJdq0howZMwlT5yGZ9GuD7b+pY791Kp/
VX5/W7mQnm4tGTZ+9qcnbAFyWMDVzdo2m9OD7/XD3u5CI26mzTIFBk51rQMjgN48yv6vQFa9DMGj
o4vu3KgT00qO/XfVAPBCRlB8291Yo0g8lOoHYfd+6MH/lFgvgF+JtW06gwj9y251o2ISKh9B+UmC
kD3hEJgoUWMji7R5yX9D4czGd9uZTVf/LhyFWzXhVVcO6iQQYuHFLZAtUmeyABjUmgLDTlOPu8EI
nD4fSettCBM6+cJ0h1kVN1f8A5jSksk4CztTxadIIbJkcAOsGkP6xy7oYOK07qc+GDx+DA/Upc2A
IPgJ8qDvo+eFTRCKlfQ6Mpm/im+7NxDaZH1Yhfd8HHnP6IL4+71HGHwOSmCQOQVSht2Yx0nOPukS
kQ//eUC7DKldec5yr+H8iDPIpUqXE37L3UVWoBqwPy9s+ejaIkTyl8UMXy32zSiOjS9FL/+4wUMk
12KEVtAYj+CnUH3VdoYEk3Eot0UgfUwjC8CabDNNobC6LZWST0cZ2vQ7OuVIFpEYv8RgfBF5VTZs
QDUUx0H/jYYQNjTcteUX8xSPhZ4Urhi8Bq5KAwqi02JYra0V/WPbgARfIZ3D1ysVm9RQjf9tS5mc
UbQpd37T3zAmocgbXUry9BDo0TSp28ECH6Zs6XMdLcHgP6XuXmya7TfBzZbSH7QogP1ljJGA1uB8
sNoc34U84t86btNDSXlNJZv+BCkD7CwIuBkr0fqw/83rrxuHYbzHqT4VWUusz8JfgoY/OAh4MTcy
nqY+i1y81hxSMr0F9xt0CziRJPCSNLjwB2/Uuz6mWNGwOJ1ZnapgUq9K52IOYvSyLlolxRMd/S4S
gHBtBcfXHaUMgYJal5p/s4xOtviAIMpvCjMJQnkNJL02brj2LMI16HCjL95TJjhNy0sl/Udu9t9o
ziIWOmj79A8CWAxWnLKu42MPK0ez0NMPjpse/znmnNJWhZ3ehmuxizjJATw+2xgogVHue4bozgix
rH5XjXfkLsJzcc/dVD0zsMhjyeDAZscL1/0e3pqztX18cETWI23slp/4hQBOzZOewIDU1qTI4Yqp
QAhVxdduV3/bv/NxzDoLIPiVVbcSszpc8PTgcuH/T25/FTiaz7/IK0zdUxW04IeO6DiXfyMwFZSC
luUJrB57ZXIdAhTAfjEm+dpktOMrbq2OubRgNfHhwQ1GuwLop3QSii9EmTl3366wfdFBDk/1Xsq0
ICz3DfnE6sqcn11yY8RkuylMrtIvUiytDyHtNDsJCupjoTmr/TULlkGe8GJeCk7g8JO3MiEMsmMw
vu1qhM1E69MglHuIeU3d+uAJ9jF949qilQbgNRHmqRBeo3NKtkJRgYZSVODYwHdXozUspIo4iTF6
NkVUqVdQvOehiwMxYIjn7OZVDSPulAj5L4p42wSJ5VVeBK7r+dR0xk60B5DjJaR9EAb2NC9bciJR
4SHfCLeGqeBxhsqb400HHOJZhpcViFAHY17p4OJJ8Op7iMHUZjOApPPvCxAjd9f3YcKrfjNVkMu8
2MsITvvKuJAp0LOYL3rXrgmUsN73spb+lflZo93r5pqxNWfJe02Km35OC+sZV4cyTgwmxHTxKezA
hTrM839HS8O0oAh9Ul4Q9n9JROv4ZFHHPL0UQsgwJaa34OwBTsep7FTYk1hxNtCmoh8Tiq50Zoii
pnvoPtDFh64L+cMLHNpknDGA4Ya1w1uNf+iBCAtALTwCtY8uvzCySZOF5shk9zzCiq15BfKYtpzV
ppM8Y/V7aqF7SXEQvnUrWJDLn/4EdfQS5xCIOkhjfchrwZagmgcbcKVmNv3DpxCeK2I/BZ09cfLt
0JcVda2Goi9Gn4/V1gLOzPo+JaxU3XvFeo677/dvYY8D8HlDlvOKAW3XKKYq7xDQEEnOX+y4MyTg
QCPdF5mnrEodSnktpcLDeyUfXYkSgZcvcIEQpfcOME0ZjzcEFBwDvhcMT/SqgI98bpauJW270L3Q
IwBBu7ySyy/yE35YXIwT+NXXkFrdrZwEfWLGGQXFa5GWziKDgxf9wgp5TzamX8qm6/V+/VuZfNZ4
9i2zBSLGH5l//HiKradi8WyY0V6IV+dqY1wml8kzrVQQunBDhI9p5F7fOZhaikwir4oO5S1wnChj
BRDTy5dq3/dCOZR5Gm2TrEXMF3sYEpD8kDZKbFEBqEaIP+fqIcTRVhS8l+R3TaNs6fZwi+PdqCux
dxwd5uJYNVvaLJsn/JYfv3J7QAz8froFPtHM4Y6ZAeKXHBoRBE0JaEyTDE2x7cUWwJDsvwahsTo4
mbhZwZP4Ggb7QMk5vJ5sxBlJ70mX4ERp59V8xp0qIS2TOda37l6U7mgTbrn/vOxXsa+bggXqfmdR
OFyrmRm/55YIfjyQN7SOMpdPd1nMnxXD7wT+l1oJDhNdzKzgb2zDafkwfudYyZQGbfbM3KwCi78T
XDjAwr84vmxiaQUbo/gptMYdzOXuYe7Owowh4ohZfMEuwGFwSpUN3LB8t6LIHKWXWSlPUVIrK/iu
sBis5UReybHG9DF3jmT2c5VLfL6piODash/mZDXp/ov5j6rxmf6JdZcMPEsp5WpmkAEihrvWxgQZ
erotcn+NupyZXuwD8ddDmLFHUWmRJNYta01Qzd8R68lHGkd1xMsPXN6qjzhvqKTFRRb3p/AcRb5Y
XkL537I1t2vhzT8LvriNWLruOeZ6NmheMg1mo5Kv8ciIAQBvVAVAVE8iArTWmcOitsjmoDR0PnGk
Kb+5L9yKK8AlkFP3Tpk/EC0HdbrVfgn8ihA7XVaJk4d3vhHVFBW0V/8dxR46KhNHkzi3kyBA555i
qEix1Mlc0Qc5/HbvwhRCHvf+Y8vLhr3TYKgokjBYU709wKhHQiwcoq6FmzstijPV5A0UfGQCaOx1
CQ+K1kVz6rKYEssxC3GNqzYOGTd+rZeF0PSPF5PjZh0OEa1cNtmAjxO96CHCg/nxkKvW8/B1kYUX
S+eB3bq6RU4nV9Q5DdyDPPvY9xeUmegxPIILm4ZVGrEzKY+kqjS5HMSn/i16Z7p3ZQLeUplp3SjH
n5cZ0HtH1cLrBgqAG7NqDYYFM8kQ3IxIAbuTyfDxSxG8ptG6mm19vWpFhRG/2Km3BLZgD8hAzdcw
wOIIrHQe5wowGsdke1xFZ0D3efCfAFFj4APmATc+IS0XpPOdJi0aS6dF0VLlLx2uZe5wu92snE+l
CXfAMIH99+mYPo2M+h4ZcCiODTPIrHLQvp9fOBp425WgtTr3RKLmFdqkWmSJzWwMLcKmjWpjMBwS
1oawss2FYK8efbUsdocifzhKKjexr+FdUsgOSHNKiyIs+viD/J8pmM0RkdG4EomFVaZ0QD8y0oK2
elbx3gbafSXDmabNpm9ksy0mUewNXrlJMqFhNPPqLI+uTHqX9FIYnRgj4uwiCYm1peT+G5U708Kr
Srs6PGnbi8EcPYwRvS9CKwXkjOS+N1WJX0hgGzJ2xex+KhztrRwwf8odiaLvdmKBdZHQGb8kd4U+
QcZ565jsaQjd4+/4a5knRRySS+rhvPJBh26z+DsQ6ygkwCkmvjeLzsCW422wfIDmJ7y2T9npThCz
Fy1F2uCBKs2rGxRXq0lYZ2sn09XbI/MHxfyTJK4HTONQJa13P1hXKO4NwP8esORWQ1x/FtgnMy0V
TPNkMCCagg3zcfWRxaZ75uwj3U6W7hHUj+5sjlAM2q2W1kXZJrEQxQeaiT6DjMNwuWZhj+kVYR+x
6SHvVq35RcElsp+Kj4iysbsFb/t60lgRqJoyVpzAG5IgLa3PItErveL2rJbf1b1efSZmdduCt+D2
fteIKxE9j5cpm/tzprHCp7DdIlKi/G+k36DiEFex72hRHPnkNITW0m/nqMN6Hla8UGfYQNu3auCc
Us4jhDDgINBp45JgmLK+Iip+p9ivUG+35HJaTScZqmexYaWUZV+yq0XDJJy8dmkSdXkC9fYqA72l
nCDXhaOW3tedBlCld/dVEmoHoh4958naFiYrWk6hIquTGBinioyjA8Ex3SS1UZxVi8QdW4Jvty01
CWKCPv98DSFSyGbV6o8Kkd/foxcJ9UnwAh2bUbSjWM/j6GF6vzq3sEm78Q4sHv3/uPoHf0DYoqB8
EOl97KH7kdYXlnulCiAjg1XLB0o7ChYLMIT4I4aRuIt5IXv2iqXy1i5K4Py4K4BrmdfjVtxwFg/c
LPWZx0TDRqi//VJT93zd7oDznG6x8r0Jtycy851lkVBc/GdQUTTrG5bzklL2eh7mw/rGaHvYOhSF
HZl4IWzEIF02axIxXvMgZIx4IyWnkuEQJDOhqFC8p/hMYA8xtouydsnOaAr6MVNvGVNkGbbAT164
wktKI2waKKwt0WVCCgyD544X1eIW7GhgFxOdjPKVfxSDIfx2KoDbxf3DaizPXc6dWVdSF9oiYp99
Kfa9TP1RavYvdrISO9JIBzN66beQIcHYih4x3GfHsOWtPetTPIY0QNu+G+x+qxYx3w3W98n6buwz
OaDmxb4+UWRr1jQ2RItauO6fc8QACN8G7g8bkiKLk4UebCFsl88az6DcJOC5Prsj562TKaC5LTWw
rH1mq6h9NhK5rEMdesNHmaACGKQQuvPG52VfQJL+Dz9fivwpIjC4TUlNSfpT+JGTthd5P3Phfaxw
PEjLTOj2EvWxmFLh58T8FdsCQYPurw4aMlv+350bbi97GYhf+E40aPcvW3INh9r46o+Gh5VlaICb
5b66xd2VcAzER7LvHAQbo2arhTMQg50lvGBK9o0y9jAzJfNxzZXL4WLwyVLSVJRCYJyVRPYZEVVY
+YYmkc9nvEXL0c1Qc1pF0THryDojpWho9m/6UaBPcTuVoyx1mANuzj3ZWI7lDyI4TLV9e1aj/4Sd
j7QJUPXUYUHZTKe/NPMrOo9XK6pC3olpYpgz9pGlf3H5zeVlPXpqkiHbEytrR/VNuAIzaRZEe14O
xw4VDVJrw16B7iMpCiUqs/mXambixzWKWZWqZnDUoofgtBsMlvc0UTr8qFiKYLNVcx3MYSeIs/a5
Lziscz+kOv3+nkvXdzh1+Sm096knxPYUH21sPu7C/VuJ/227uvPD8FfPrll6Ainks23QcmVf5DZy
V4IlXeYQjHq14PYwh4rv7gv6fz4tR9fOELIeTbvqi/+JtewrKqleg/F2nNwfbG/Ep1IennIwUlcR
v/eI3GcMKmP/x4LE0ZchbesGO37pjiTENA9XxHhmKiLcUhuzEOz2OvU40h4v/v7552oKlvF0uome
coRl2I0ub7rJXkjjxkm0xY+TXzKck5708L+qZ0YVr8TTfUh4t34AzM/S9nlr189FnGAa9xKGKqg0
ix3gvcl6Bge4vj7Kj3iFFvGxOdZ20IVfCGj6PYwDBLjl1LHdMufbxG7I3d2bKLd9pDQzuL7BN5aV
MUu/IigGJNDFvP9ZF9y4zdUv2FckEDoBy4JC8KpNFDi1Mh47KLNlgi92ulmc7n9NPhO/tyTpgghL
9Q5FAS3sp7at14Pc4omjG1wvlizF7TG/ojGe7c9WEXMBRmB2zWFt+ruf9Y7Wo/Kl8rPPi/6+Pezi
XCwDr39zG8eabpDQrwv9/T8XJQs6bsAkjoqnodmtH8Fs/frvG9BgKo3HRtEANb8TFTZOplukpYey
0Cw5Wd0PCmaGR22DYrjt5upz6ouW7W/EThY658rnIKuQVTf//yg3Q/HMEncmWomV2DG5xIbTITnP
pKeEdJZzrLZIElnO3uLtin5DekfgFXPfMR1O9OsjRwb0/URu4pPQ450eQi7hT70Yd/zHNM+cQ7YN
lG0I82FbGTmREsFJcxJm+3I4pGe/lisfr0uv3QH6gOLIWc16fBdzkiSFWFjwA715ru4jLG0MNA1i
LcGcw/E+f+PsAa96+UQJpJttyZLdy4COjzs/ze2riiIlRffXm5xbTOTxPrxhAGFUOhooM3qvzfEf
2dmeQ6IXsFyBXNBvNrXZzO/z9c/+oVQqDk12275OhjglA6Rbrwvu65eElHh+uCLZWOTqC/qdGSGe
LU2j1rUwPhrMZIasjCUkcgj2aZLRNej9vdojNU6UwCFxQ1GXzqlUpfXmBBKvuougr6/I42sGzTsC
8mTrNPt+GOkOWuIww78z+BIg8Nk1dy7vc6TmT9suRojNkzdDs4TvMT4LLloNd8ahwLaA/kO7ZnPD
fAr5j49/ukI2zyph6iDMSMtW8zNoXNmyKuxI74xm4gKQDR7EBWoW+eFf+TX5LyRZOAVkEKDnJP2p
bWnIRJjXKCiZ0QhYlK38Kxg8r6XhKybINhmXZYtFRlBF3Toxuwm3qnsLK3h2nSrdpwKrQX7In/dM
3lQ4PT6JVmVALadqfki1R8LfyPYoCWm4Ir0jx4IvpOCoL82yKjX5NfbrmOQ5aA49Flol5+OhnXsu
1leSATGlYTAW4pad1qXirh7FGllUQYkSbe9R1H/JYCWcyOs2YfGLJe3uH3aGXLM0aznDqoZCV2td
xftLirZ0HsckO3zOLEFXbbzmrUcMZFmmbVf1dgnzW7jubgCRrOy5PjZntindxfa/capxypR/w0fu
wwcxLTpb7ZzB+WvemQgz3SmaWQnQ2q+f+YvocuBk/bpWQ9tgJZG8lAz15HzSOksVBrurIkKuY+bb
hAsk00W9qp/MrYfLkUj2q2TNi+p0GHW/sF42pwCsUWeWZsBcpockYpXw2CHP1WT+VAUz9RkQ1w9n
wpn1XcV8E5N1Aw/p1cuoY0XEjAOXSmk7/XruBaPCp7tSvl5s4yoXaJU7342LOK/5RLJo2xX2MSI1
lW6JZ5SwsFcVznxLl1iphlvRhOZmHn2YvrFJuI49Fy401kyPyl1NAMcOdJFkl9tbxs2kgNDOCxvL
6XrHBuafqhxjAkBIubLVvgSB9bQDbwOKF+LMijGe8e3hbzgn8QKG9F0lXKxJz686cSN53WSA0DV6
n0bEee11dlYuuimJUwzib6giyRFUnJKBtlBqi9RJkysSC1WAKBpGDNKzcME0dzJ0i5BfhSQd5z+j
y2+hpWGe4YKJqBIsPO5K2/kc+l41xYwiYZf6xdohIsXZRekMVZ/1SOuIZ7QmmYQdyqKn3Dz9GRB1
hUW5ed39QjZj1eQQlgTyOGlnmZbXv9GUTYAO9FdODfJDTO+89MrDYZms3P2fi74u77DNScB1kajX
qc2mO/Z4j+UhDVlpO4ihAWXkNSzYENTsHMTcb7JBfgyBMT6uHBQm+hbcVATD94lF7lCB+s/mM/W+
Ol9gRTRDDgQs8JEP3iTRvmDnst8ADvk8K+e4EU4cCRj3f2uba6e3mXNbrROnXGTFLmnnmz3Da4DG
I3MMcmVKZagfd+zy32lXBaiysEClPE7JFQlS54r4qQG2H80HSnRbqxxZsnhs45e6e0mKF5+T2gLn
lfm26vm2uxfqUZa3Na6wqm6l4soWiTeSSkzePj3gpjjnBKgtoWeld/MIAMhIBhiVO2PS3rWkFdvM
trG6MifdZ+B4OzAMLqwoqU8w6ItkDP2E0X3sSsN/VkR9v6pckMRyou5Co47i/L4FEOHkT2fWPxLh
7DE2rRSnbJf+NDcV9Y0+Z0g3PS8FVjrxO05DZ/KjvQ3Uhr9n/ePclfxQptHWo7ZXfpOL+xSnsrBg
NRIubqnX9Xxbpcbl2DFgUd35IGZq0uQ1jb8KMPHDUZmpywfqCb+1uZ242OWcXnbHKrpcs3VcW1k0
0M3y8dRNjXa/CImbf33/I+nGXDXqVQGBHhuE0Ugrjb7ySA5TEZqABSt/b5EAjJku+iADDFtGoUnp
g+gN6hNYN38gtY+fJPgT4xpaBl8e4LaYHlJ8UiAk/ublGLDHEpX4Vs934d3ty/I/SAWOeuG8xs4W
9Bi5qOAQQM/4JsJc/Jy89ppbBxZ6X4dziak7qq6Gne7tUgo42BHrr2SK7ZjqK8+rFalD1QaXDgSd
s/lPzmSB8juTSnfBNxG7e/B5cHYbn/0lWqg2glSHM2svhL6R2+nt2vh4Bw/fySFfW2km+PVWI+E+
ch1EXiW+Q7z8uJaZmNIDGcslK5XIB9vGn9AHVcyhtBxAoZTAMk4WZ61k3izWrBlZLrBPwAM4WmpO
YCemsRysiOaIU+PFPT+FZ4xEb9o4J8ywq5uSIVbH6qB7nMCrPzL1L7EtkUM8Vq3WBfeeD1g6OVtH
19wrV7fB+aQ4hHnGA6cHbylX93zlxe0PJgx5Nq2E2IXBoUUHRwMsOCfLLKThn9Ogmw045HUTbtZY
1xleVYKZjvsACWFh2I81iYYcwpNAAWr3/tI8EsmCEMiUJBMgGJaLqr+UKTZfU7Z94xHPu2Tyh6oK
T/xTLwdFRpgoBqzeRlVvBlmMEj6HLa+vArdDs3JK8L85NrmdUg/0R8uES4h4sJoNMOMORVTtR8BN
+hW85Z4PtGAbus7wNVYgdCQFnpnw8inauM3GP901PDjAjr2o3am2gf509DbyT2amD0ySWkeATKnd
z+VXeMP8HZosj7YKhfnBhcE5ZROMib3tWW7raGQ+1dsQhSCN/pyHPk0twiZXpVYzFY4NnwO6+sZb
JcpyeMShwuyyMBnj0LOcrrw4H40sZoXaafA28V9d3OfnzZnrYx4VPoZzXVrE00ui1um/RI329ypM
S+7+W5gwtDw84CXEG9cCNJoClm3i8o9q/o9tPPftfZBo7wd4+nywri8KJyep5m/ukKVAaZe2KbEn
qp0nK0eHu2z9/hal/AomitRp0YF7z1TW5YPmpasCPU1Z80kUvV70NEYItk582BR06A1Emw8lNNmQ
KIP5AnUtZ4BDiNzo3QMX3REdGaiJjgM4S35L5XoF4QGZ8ZQ4MhLrOZ9SaVwoZck0lt3Y9ApkPTS7
NnwxDyLy4eDKvhkZsiOAqbVHqRAqWxV9ZVXklWI6/F4RFr9W6wGppVi4Fc/fimtW9YK84XLjNzG2
sLVpc8SFbn7CeB0ClcjPHyo6R578iDvC4EkN06HrQxicBXK71COQ267U3As4YxzhwUA/GpGynDtQ
/5hh1zbs30kflfLFiHJ4Z3DtegrUQs/xm2DdnnkXhnBEgVzoPKgGNehPsAH4Ozpbpe9YT99PyNwQ
yNs/vtMn+C5pfei4WIKpNnLpITefF2JvUz/UcwPMukJLh2TFP4WgS++pPmJDXbR7vV1lmnWZTAfY
olphShv+pwHvKe9hcnecior9PyWAhTHLY9XaOy50Oc2ILe9flNEWLU2N4rotav6LQMmUOoxV1/GJ
OFlST+3ZthNeP/dvbsHtEOOm44Z4qWlaeH0lLBIEyCVSU6Cdw5XK3kuZrdS6mrVVFI7kUd3lRPsS
FWHsQugaK1VNdcuypH+hnMjysPCsp545c3NyjoVee3S4Ur3HimmH1O80Mh0AsOTsQYeo1uWOgNqy
MqJuSx19OHJLeV4e91m36craCYxHzmQa+DWN7W+Gi6AXLwHlFJ096khVBAd2+qu+VFUp7Rt5cB9f
YW46p2WzagucrEUJF7u+dAKwbL+DbRje8oFnhdjqmhBOSW2f9ntNU17BGkiMw7Awku3+nzQf1xo/
VjsQdobg26aCVgrkp9KdP91PM6ApLRWQR2S2j4uaz8iSd0+JCBqOChpt0wX7hsgn1Lqoydnk1iKW
isc7nbDOurWNu2I9+FsZ9t+LyBOvOTNuWQy6q9WWtT0mD0T+vvGY90udQsP4j+UGf207vy6ck+Dr
KIrAmuocsXnY7CXfEmOAAZu29vQYFpbrjExaTz5w30AK1Q/XN38L+REtbfIeDAQTQTTA5yM/bt1L
9o5uHnk7958DJaR05CfyagZv0Q0JKWXeR93XD7DTgKyoa6XYX9H9MYHYdrUVmjaGIqP306v2vZcY
X1xKKkUjRHkJlfN2Y8pdkWmMkMiEhiMDM3aversdiNUyyi52HBRKQILBlzlAvkXbMQzaIMboO9Fv
CJIInxzpUlTfGKrXDbs2AAJS3WlU+A4WGacveEAGGmoJvweR8AO1XqQam1bxxlTszcwdgsLPhE3v
EWfNQ8CQo9oLwEmJVEQY8/IgrRStgHS0RyJn/tRUiDu+jyMBsozT8WQgjllgilrmGPaqAQ+F3vti
1samREjGjK9KvBUt/7FYDVZ49K+Yvqj6NaAzlqU8hYxOIGpQhi2gzLth2YzzTEaTei/9jltGEg/N
K0TLTdDJiZK+o1tIB1j6wnZf+m+ZCTIK0rTNk+/lCmXVKniSHg0/sVHURW7VOc/ZxdI2SAsMtcrw
Wigfv2A9G6b8T+Z+De4sMVZjRXlWtmJ1BJPxHCYYJB4JPX8MjcrLx911SZyvB1je+zYlUyFrdAj0
65Cog5Ipehi5FuKc8IMO06XkycZqUHdb/DFG4ipZvu0zul49TxjarI9tW13Z9u2KVi7meN0V52AA
z+1N/Od0Ju45LlmC80gDVlim8tP7/Y8xN6MPl06/aJDj2DL7zIjKCd89695ewDEWe/K5Nt/trpR7
6YmjQjWR1msb9FJJQUDmH43YJZM05Hb6TLxN+oMf+0ol3u6L6huYK1mcGCQv9kjYpjP2NPRkgi3U
GFmpRqxHHI0AhMAadxFQaQSlrFhcE2cKoakMu8aywCH+lDAtjIDf3Uv0jmiWfQl1OwGzlsXJF2nI
FahHOcEz+SVi+A0WP8nH2I23qPTHeP+2F9cAdHlI5GP9lWyCZZGjkrPrTBrYjDMpP50nuvSDJaf8
W+VS1e+H/LoAQYYvWe8QU3PGoVs5XPiDoShNQl82O4nUXKoFC98RhWGAanjf/IqvssONb4Y09cAH
8gUiPYlaHWnSS1B9mRJKEmdeG8dYnUOA8h5GwQGcB6p9iH3xObdvQkZZzzhtMzzm9VhEWB7pvI47
Qi6W2/9zgNMiAXJj32zIcNjlfDZTeQIFUDGGqUbxhDcBqerelymjAlaen4Kij4/ub+pINP9ltiRv
8io3c+y7cwmuz9Qr6jGZViYw0f4JAsr+d98LrcL2tQ8Xe7XZSn73g4V/61gP2tclUeCZrs6jWs+l
FPCFvB0XM1DOzGtgQeaQHrIn/1qIUdbKOYtLvBavFPckCWQ/dm4BwYDmgPmyJDUOgnHM0EC4YSMU
H5UIw/5iyV9K6/DqnkZT9GzNgsBpGOXEwXsI21ayXsU6mHxjSGdY8xdV+M04ni5WAVGW+Vk/J95+
05eXOIRQfbwnHK4KxJ2I816i7ShnNWvGr/c2PYOw9F2Hy83nj+7qnesiFjk4gqLo8hFkrM2UlCsH
Z9EucQnH1TJvEDVjIjN4XcV4Db0ntT676RNYOI1FasEp+QV/v+BFT3jlr9AfJdciO9yYUHMT0DqL
fGKUCz10NDBx6kI52ac4QLu7/H06ZYaUmQMf/zLA3bcgcWkW9hdepi757oK8N2TIIXU9ocyYr3P4
9xCLT/2R9fSFl3W2z4tF8VLsCJAkQuhak1pQeIlvaONBqJpHbgzEexb47s5CmSph0dmLwWymlZJ9
ws1iqvcyfGIrI/KDest+lauWj10ZX3pxP7qBmThp0zBAu5aR7c/Kwt6C5QqolHVRObX/Ih5+Bn6n
X231GJCnYLm3m2aFo6A+WYPQ0KCCxBwt6WeS43G48ZzwUSqnza23DDbscpMkkCBrR22LzhKVqdpL
C1EOD3J4xQIOkuE8nDTwjv2mfkEI+/BaaqLIIrUqoA/SRDEWawwhe1Shy/guXC7iFSRM9OJVxR6H
rTFrIY51tH6dNOQ4H3aBEuM4/z6HCgscCK0cNTjdNSiSwA6UfD8awQD16m8K+bVgMLMqgGH4yqEm
kyPEtpGubtt2HgNrYAbCJyZxxO4Zx3oKVMMM9H3ifdpnfsOrlbCbaQ2/d39u+MI98GJ3doNFqte/
euM84lSgt+EUAoFZ8NtoqBmFm1ZJADmnlEdbexaQ3jFVhdT8rRbmaoIbH2qb/kBd3u0ea6Gsz112
MFXKx5xxHZ6+Q7yUmxCcUZv8mgBl5Zj9mPtdi1ndeXFQHXnbJIJAwBzMedjQ+9Q1iSMHq4CySlNu
xBZfr2W8WmdY+RK+EKldv5tWmM1aUp0dTiCf5LZauD2HK6E6tB+D7MOD4IAvC01PxY8NAnv+3thA
VCij9TQNDyJuWrdRaL7Tho9+scO51tMBK+seqdWO4DPUneYnE7MU4XMrG9FScSpBuU3SDNVheFmy
o/lwz1WY792vHlXmnV1C99Vas8NyYwe3TZOSN2c1OOkfavHpgE5lx1/D+d6AMxOsdg2AKDxVf60R
7dIgxDlgnUftKoKrXKvMvNagoGmLQ5grIZ/l3nK6TCoHZzB9Ce5PplAHR9bcDkM+HbJueSY/eKCB
jJr1K4oZvWeES172mCUhjT/42GDcU+291v7GXnIqjuqKf5a9zlVKQUOCrClwOlU6LvS1AYRquug4
l0o0YCqo6RSBPg3A6H59D1XBWgpvL75GVCAMzpJevq3bx6sUCzwv8/5pWiYaUgLXbq02gWCVEZTk
atZUsFMSHXpMqq3dwgqOg+FFniBXK+HpRx0VaVL+x516hb5A+A72UFipKPft6c6GMMHXLH1iSl+G
ThmGoGRCpO+ANK98V34gNtGSoogNjyaTnYP5RRyVx+QZ3jxqITlzWfyinGys+yuLJZHAc7n/k7f7
enUtRDMi463Amw275DRXC28Qdyi8KJExy2zX+w2+863Km+9Gp7exi+07Ys4hWNsh111258uLK0E0
siHNtB/jD8PCLREe46lHmKnjb1Q6mc1U22s8aU3wB+m3PXvbuIxvUiYqLXT+tROiKa+5zfPsPGBA
Tc9xIJgm7XSu3NaRWkblBbzMAQstZ+LUstGBPLVxd/Q+3aZ4/2M3FQ3OzjGkW7KXRZwgN8DRpBAW
R2LYtDOZ/vLkDbKNLH6jwwgVIjj0oblrwlo06c1m5U06dApql7g9GkqbjAfgCKFUWKvuP3cOXgUm
zXZwvNerxU6v/1m5Y0vPtusJfh0Kvu0IoFfAuJt1zJQS3ik0yUiKWuoEgysmovmXnZRz/ILjVAdU
dOVoTpn6gK2iXfJJ2GFztwFPKFtPenn4mVFFHMHKyort5lZpbYCP/yr29OIKUs1XXDelYEHLblAo
Axc595YyX9J+bxPCY8Y58AZ7QedKy599JGZt1g4zXk1L7Ljv1Ly/IHWK4JNmbztrjorFsPh+znpb
a7prTDedr+kD4XBDAexMtdX0QL7fGlFdJ8K7VOctaXU5jqbbnYq6s1bXyLHtS1E03mTxbeRwaq1y
XiW6e6ii198dyLhOAIvDqiTdjI9L0Y2gCeu4sgTTEdzxYyf+3t3hKg2RnpvoLiFvdmA61kjn3C8K
sbbKkIesBhjqtX78gRkFsppxzZlnXrj48cA+Zxs6WfjameE9UhzrQx5IKG3/dEMr7ocLdJWjy/pk
E0+4Uv19PpJH9c2W9cOoMMsJryORhfkW+QLtZc0BNUdKn4+AY3F/92zETpRSeYKnDCOuf02qijJo
u1F7PArs78+m2Kwe3hWVjwWqLU+YHL4VrkyjzpvFDlmY4ULHX/V7lVhHcmc6uWGSPvpn4sPmAhIC
yBfwDCFyhCOMW+1zexN82r7LhMvNKa+8iRDchkbZh/KfkGhqUtgkdQl7lpg/9m//EEU0Pc6qrcrP
f6Qv2eMvCwmqSLV+NUQqomScdW5ivqIV4eKyXhPkhNoWlLL5SgThM0my1tykpbMJhwnNC0xWpa6p
3nyzxeEkUvS6fPsi388t3yNSs82Q7kRBXbSQQAL/9fzBfC9Y8x6KFK4//W8iNaur6v6eGC7M4CvP
EYTh3yPtgJJPGLw6gbPDn8Bk6ww+rnKoPTzL54FoeqlNT1bE8VwE3Ss/lBiGGd0AYw9zYC8Jd66y
eky3d1PuQclDsezQWCzuoFD+qDnvOK19DjRMueT3iMX8I230GpLnF/9P6ugnMp7/VC8E1G0L0AoQ
flVrKqIsy0no5OFtePCljRx6WHX7onjCGVYAv8npygVImJQhbaywIqYHq5lGc+LV7o6zpAvSJ4H+
l2zMHHKaiB+VVPFTnHvirVqn0WqrPheAAB5yDhM1oeVjuR1JjoNrTsF3S0u5FEiyZEdboK5QD+7x
x1EOkVUNfJS/Y6MXqc9sNfOJXKN9b6P9Yf2c1RkKnkWevxrK9ABf/V9c87mMUI3A3wxoca+v+YK3
GRwN//XsXvn4qWUVUSfz1x5BCcXAnxkgBdHRXUzTZJQyF5wB+48wcu8wE2vZhkp0gtMCjcmExuoX
z5NksELJf/MLP5nNRt0MomAjHB6qrgqWMTWOX8cAk1OIUm1XUJucqe1LCyLJnJu3D2AabWECIqOV
HMgk2XtXthLCYeKJ5jy/rvFaAjhNRFAgsfAqtitqSPOPXI0SJe26Tx9x+bMwfoIAEU492aE9ckLV
zOhX5DU/QAR5RkglNgrefcn5ROE2dM1uf3WObItEvUaNq1mXGFCY3aP2E6oki+1UBmmnPxGPl6xK
Qh+oEc5vrcQ5kTjVgCYHMnRKKKTrbFLhB0TF3i9Rsa2DBZHeffCiG/5FTPcC3rfJQBX0/mKjSgPC
5b/8z3y4iZAMYi4eVb1Cgn1R5yyC25IYQQ1VDnXHnXt5xILsVbzkc5fV9HLGT7sDXcBuosI7EgXX
C1Xd+pAD35qYFjFKpLA9CoDrZRLUZa7e8YOaPkLr8jbNdCElx6TDLmw5vtCQiF0vjLHNhuw1NWC5
DRHXdGup6mFSCyvzrm+TzOripo8cEAhW9w3HCNe8okuwQKXH1hhceq6DwTdYPyKjjUviNBuT18gw
YcOrup8/l/1wzC0SDX2YRS/1LTvnJ/18ZRiKGC88+XwLDxxYFuAzQkWb731VC6r2q2gYkftUBiyR
BE6fh1rVYIrxtV2V72ELaxjpe0bIyu7LvSLrKgtZSyP879H0e+Su+oUIWWLRMV893Zct6ZnQfu/b
rhJvIl0PmI0nlscBW3AHMc5I2Q7piuEQuJSopA1NEQ4GuT6JbI2gfSS5ULDkcre5ZEEMmpSRHsGm
5xOPoCibP/DCNEG0Zv/Av6qQLeJUTOdrvGoivQgWHMphVHqjwsyUO7ZSafLp+4/2Dotm7PyvC18o
0aM7Br/y4HDrvBnupKXuI8myG3mq0D/CvEua7G1UjW999cUi87U8R5L9AESaZE4ty3s44gOcmdU2
onE/59RoqHfCr/R0rEJj41TPJciAv9JHlB2LttchKcFkawjisePGFhIxeWvW2BxggXw3JmyZMNtV
ZY8nKfcoUJAkWg7hB47jHKfdbJb+Tx6Djn5oyd/Dbzd7I6BRRTvtLnZHQOmqTkXKCc9OwDpYFSXn
A543AhV9QWyCn93r62ewgMvpHIwm0lvI9But8mQV74Aw4dJUAf4V0AHgKyAhPr5ScH0ATx/gk7Tx
96wsK6cIE/93HY0KLu6ldP+kjIfzllh4UxwXp5EGoBMqQJc8lsQsH9JwKR+ojXnaXl+eKtFYJmCi
5ofAc7hhLdAWSwGW6jJdNTrGUYu2IzvhTDdsElzb8umnfA1MagXR22QPwkgQelnhEAUGv6OvtQZy
dtJYsj3DfsaGGnQvMIgumRuz0y+xCRBfno8jk5gAK04Tog3QkGTNRHb0Wm41ZEr4BU3M2Bjo/WQR
DVOiDi4tbvphKOTRv/TLg7i0jDVEkpysKU9WmmECHuf3G96uYOXJ1y+qfjPdNZ+7iR3hmnZSmWK/
UQpbLTUPuGAAFk0Z3VrGAw1N6kZHeQrMyLb2502Lpw9Ou5/+uObhe5ksnzZPGx+ZoZMcfuKIPlxZ
APgNqnPm5pMDmFawBCp5kYRs02lGMVN0nHAhzf51miDa7lTD0eCBE5hGhNXeBbu0a4OoE5qENXUP
s9nohWMmlCs6phKlnxfXhvN5QMDB0Cp2x1W6ZVvqsc0jO+gIkTozxoBNuI4QX/0tUPxeq/tdjhAx
9z4yv/Mi1eF7vsBbj6FbyagCSwF9FmQhS93pcEqlSor1i1DGPJD1LZIkEX5Cnz8fJ4/Vq6+XoJ+V
h0DerGZWI1iqGEilHoAEfefIIIpszkNBMO9P7s0CMR+GUIZEYumGuPU0K+FYMuMZHVtlJRj71YQL
nO5k9NXZLIde8MooJprzG5l2u1gDNYRjTqBIlVC1ZREOZpAO9SUKvphaeqYGX6MO5pgTPRsWZza6
W/7e4ndRqDhC20YcZ+bl6Tpnlr7GxvSxCgqsK0MM9mvBC3cxzWxntCy4sAfszrxmJwd+vDGJiqaG
thqHezmwcZ6U9vH6FMHjfYCQqxOIMn3D0A4cBZe8YBRdDNu+hVybfu+iVL/1OL5ojA/djGiAl+eF
joDPm/+vnnt0UhQBwRrw60K7ef4BlVBnhnjRlf1p+FIPOVuCdgbCJ5X0LertuApDFbiAosnAgoid
vS+YjJ4EWLjc/SUcPpEEfa7N9HkLcmzNtQVu3f58f3fNKvmevjkwO9NWEpZCNxQNBB5ztPHdram7
8FmGSbpi5Fqbb5GPgRONaJrNKm6ZgWz3pprZCqM4o3tgUZzyFLq5Tgk/mS1BSlvCFFSe4ss3neCH
/y+qf+XeIAFb6RMg+TdaYGStUZN0+1aJ33LTqtuvjBjnIuklKi5chjyn2r/ovClEYilLUiTnc90P
RMapLdacPn0LyMuyJj6SiMByXyWnWO67VDfUZ9Gmr+8yokmzC5xWb0qkEmNey/UzDJCXNtX7GFJp
uX0j7Q3mI9xmrtcVeLbXDmm/d8Z87IX9/BSmyfzpU0MicDn9nehtIeaoiEugbhqVC1rUq0hhGyd+
nLZMi0qSuYXc1PdYU8QwsLBmeFR9V7jFqERbbQrrKvJFdpuV6lw++uEcIb4tfQqk8/DKSjGfCThU
GD2OcbB0n+abHHrlC1nxTsRhv5EisfzfCpjQEtbMqZynST8/ZH9VDyRPdNPwSK3EQoXJ05QnuObT
/nC26bbnw8Fq/lIU5v79bXItj7e9H+RWUJw2BC2P0elL9V9PLepZhvgHSIfW7eUVDRFoqpRsIW64
vDTx1+b8L82lg9rfZjOePHDiJ93YfKunmQ947fg6ilx1Sz/68p/DM5NyCz/PJs9YPBBiuN1HBpti
DpVXoCoEIkR6i9hArD/CSqAEuaJtuRPhAno6YQGjSTWQza44GLaV693YruV7HSoQKJC2KWjIFqbP
j8C2qVjKiXsaPmYpb3xiyUPABVve6nik1/cTLkwugxv9PgJvW5LldRtpeJEXUwc23Zi84+ktqAtO
K8aFfLZp3AzX53fbCH/nGSuFyPRnFp+UqVUGcCpfn3ihqoo+3KRw5Z9ovrXIZAVxbCfKSOPAXajC
CGaAGNnraz4aqa/q155gP6q3FdP409fIiUaVrtQ7H7bOvGeZaRVbrpeh7sTUu2aqbAVTir2aO5R9
WyAw1sX3VHpVE8KJodVaOhd8aefZmoOIIMt9jTRMzJVwRHiVArKZhxSiXh1Hh2P1x3E70g5NAEuj
syhCga42ZP4NxTn1+Utp0NbvdkID8EVIjnciAOamE0dQtfsnl0oDX8kmXyVv4Py1z18Oxw48KEp8
RFOasZNoz3M6HsqRaOJ7/0c31ZTNrGAjGbolEvP+GLkneMlzAAHJfZlB9CrwyPF21m9W+7/86uN9
A6JCuuySKyOIOU2iZy/7B+ZJPTJkqWJIZJdqjVJytKftm0kr2hKZQ38t7AOCixzTLQAwOKeNvCVf
/c7ErxWT8UxQA2E/+l7kvBDOZEuKUSFRot/uTmCGymb+ioFDFhOAgFX7aVUTaPH5dJASPoNzDphC
hJsNznx6wo0NlT0jfh79CM6wO6Vaq0yKXmcSDtQL963k+H7FMZKz0ikrJAsMtf5JdE0jdpWzJdCG
cQCUUfK8yfRU1tUl8NaAAeF5MizOuP8RZLuWIS9shXvf4SXz9mjllpYG1RUjeYI0d+2TA5u5CvLM
Z/VB9D2kVF6TtK1bxtxJUVxCUE6+N8k0nTRycYB4FL4NyitK/3mkH1rilj/NdXIFhWKGqicIScY4
Zb1p3h73UZqONH40xJMgsuNI+8GkH3pFx6mggaRqJ6q1ZNYXLGACVpZ2TyTgzFQXEr6ElpBlPwpL
Nc9EdZ6xl2Z8kEh5BLJQCBjZ3XFPHXZpdZA4Q5zXhjCYbTv+nxj8/zz0YYFv//yo4oDTxK7RkqVO
sgNcjJemXAkR6w0MBUE5FQAoCNIj2veqTcpcecAaRseDM4q40g4/S3zxxPQTlOTEnfrKeKlYy+hK
Vm07Q+VeKOEKROObMD/n5HLYYP1Q0nBsEsjbo9qonsBbYBWNsxVUL6FrdsnIBDAYHUeG8zNuV3z3
XhvIwUQA+9RC4c045JUNTlaMGVyvs2nWOYJIJ+6iPJ9nwX0xLd9CtA2Qg3JIioJr/PPZR2wDBBLk
0XL5Ov5CLkxLfh4lkr2X5cDeCponm9FHHijHYFCm1nbUb7vYjHa2NF/rpDYQh2xmVKGR5McQT+V+
n0F0wcjq642nLHc/CgLiGgLefW4If5H/JQt8/BBZM265B4VQ/Qx4rI03VxsqoKXGuwhku55Qe0Fl
f/F18TuiFIisfs0tpCn7hk6yXMFWsDwvxrekbumcOiFIjsIVu1t5PfOFOkBDg2WbmV89kz2RztSI
nkLYMANxd79Rhs5kgqY4n45z2ZhsRJmOMVsmZpAHUDTDrlj/ELaIjXb+7GIKnt4DY5h1xKjuFBiV
3MRtbe3aVDkVa18lq3BMajrjekUkfkQRXCJlx2IpnEJCm5V4PXhVfKymMz4tEex6lOUKO6JYlrgX
ZPUBS9ZxNjY1V3tHdseeDgPfeL/vsOF8hD/K5Cr7jFdq98XA80Y9mkH0c1Uqy/bp/0qWlhIqJmro
wcyz9hrYy8W+CJ90k8ZnBNbuYWJ96PuxreroO2q+NiVI02v77HC+xwQJVZ+7MLL2n2CeYKOxDX57
YEjirCESZXLK0eq1KV0itJXF63hbCuUgVvNK6AsGoiFeRBlIrgC7iAoZww3FOOA4LL5Eq3031oXA
GoOZcDGpcGEtNErdowm7vFyiGe6zkUJK6zcg2BYZEb8FqDBy329O97tUk4jF4jwFEQ0lL18Auoc0
AJlsqD0407FdH53TkfvncDku6e9KlbSIytokR+ImKg8tse39nbGimztBNnK7fcehKLntyndfq0dq
5a237WAbCnj93BpooH2XhcfX3b89UeyDX71T6JsM4+VoY4cLAu49e8HicPKQcuCKLdYzRG6UBB6B
k5QsUaGn/ePQT2xIJ0B67O6qfIWa5gzS3MiRTBVfNawo0xsNKskLh1EuLAhikS/Hj4fmaiFf1xkW
sApe+Vg62j+XXrwxYNnjB9R6/XZsYtMlfXB7KMNED3P35ZP1PZot/IOY3D4Uc6sglzbfs6RfUKJr
ClOfPtoJ+GmtQhrrjo4cJxJMnCYQQq7LfqDUnLQg7yFUVQ3Z1c5Vm3USu1oqX7OwY+ZGetCsjlI+
E9O1TVfIZubTB00Jal8mhZM71S/mem1e9UFvad2UovIrDroDBtbMoVXQNGVMgiSK0HyDZgpt+cr9
6EHrIauiNiI1w32asDCkZH7jpJmzj+9ATvxOkwt1K+kfMOe0fHvt2OU45evkly5ScU5j8QvJboIg
HLniJ7PNXhzdzB5CBiexxtWpaKn3u0WBt/0TrycVGixbv8hgv3pYd5Aqn9Omzu1zp/GFeo6MGsrb
ZKMYJHiyeFgwk43uALanpg4RJmthHK7KBF1+HygjpPDJDLpud3b5zgkAW1ctfNlvbRIAcCyGsEju
39H0PUpC8U9mdG2sGHn91Tsbxstr/4CbTBrIWkcYomWBRTTk9ePPY3lWd6USEueOgp9nKjnoVKhD
3uG6pgL6NFS6mUgLAVko5DfJYQwpV2sw2BUcd11moh6ERL3kZoCZ+WbDppOTbHOgoaBTih4T6weh
xB+UvtrF2sLEysjVg5kZTtZgKNm7gVaxErGyncyPycztCI1CX+X0EvYf/uWhzCw47u7EX3oxy4PD
1+I1mlaMYhliLHh6AX3B6BwbwkjSc7y7T76MbfV/CPMLXIjedHYFBb3f+nFzpRvGBc0zQfJfznf2
RZkOo6dBy6vDxYBkyMEnyHL1jLwuC0OuuXRTLx9gs9JVjyzF7rQe1XT4v8zk2wLTgQIMZWz2NxZV
AipozWLYz145nnKUOLTehckJxab8YkW6SUAIyc6VxlbjgAUEZRbRHc3ra0SvNy6YNIgPzDV9KgsO
ISzHOoylxo6Ydjkkp3Y/ndlWZSU8LkvZMp/1czp6HVEALYx8pQFExFzoNBjy2cITOBSRWucvQxmk
sKEmhxr9QYN3SQx4t8bA7Xx25u24969uNYi0RD/EMcj4h0tekUHf5N3aHsoIrVkmTrur3mxw1bZj
nZatwyF174VYzM3v8s+tbr7GJm+v0ydmMHJdjGivNR5GPi89/ycFpvKJq1xA0uzDYG+aLhw6bGxz
IEmPzMaP/WA3TRzBhSSoOP8ByIfpbLpeqd0eNKjNagnX8Xzey+iZ4qfkzv2Nb5BQpahO95D5D2oQ
UNSesYlqw5fsNfEVCtWP3uUEab9+7yWh9dNeqQ2k+txUykb+kK1WjwnDclzRMJG27nthd/NN2QWf
EWt3iYNdhH84OqRKHNbxilCo6gRg0zD5+KSxCzOnwnEp6tsFlXOXzrsqMUMiLsyqcXGFKIDDn7BU
WjHXIYzoEac456EEij5mmUmFiuBf7oai6xN/JWdDJPqxGkHWp6WFlqMuDzfof0guiA3b2xGDJkwh
lPtQvdYTjPhPsD72jpjPvmK4jF2Y7lreUoZaaAPNPXvUmSmX+aJkcdtlbDY5BMs1Nz2NFQ/69iom
/6VIN9xLuEICAr0UVUG/YHcrRM3foI4AKYC9r1P2ZnZ7ULFiBX6GCf57cL0Ju0xaTrVYhsPv4mA1
7kURKY4Z3PtrucId8aScZ8vxE7m8hzZ2IFxRKlEbi06DpTxKQJcEktOcUnu4cGC683pkUML7KawT
MVGt13+nwy6hGTFqW3LPCMf05fJAXKmH2g54Ca4+M1C7kgKMSy7N5hyYbjWjNy7920PjmI0A4C6t
NLsnlKDwYVql18L7vp7d5HJHWpDDoM1VPsXKqcM746yOx5g4389cD36XTBAy/Tenz2UBDUWyJnRG
oWj540it0IiJC2G0kr58BOgmYp2OZZd1DNMIpcs1z7aYnb4AVz1kOIYK2q+IZPTyh+73ltDoctJe
QBq+RaXJIF5V5rbo8q2cckaIYwLHR+id/fBBp7qQQmoT3fHjW2gWH5YZ3kgLthgCW5okJ9jLCOj0
K+XdjuAuPkayET7N1cPlLuNHwVRgy/GSY6pk1F5Opke/91r9CTBrLWSz+ugKkw52WW11SskaSD9Q
EjCivWm6DX7q3tqtl3zeM9Wy9ZzHqRcukiom1WYqj+FDP9/Miy9n4nktkTuE2KzF9AhO6O3UhMq7
s9lT6gBSQIYUh5TBmb3gqe35ZItNNyqkrQ43+XhdKhjwv2OCtSwgWCH6a1WIpSiZjbKULtIUzxGj
LUuyZ2vD+18fk3+mEjqOEDcjSNfeuJM1vcDjYycBU13f0Nd2W+GuCJ3YYmQx/6nQ8FDiguk92C/T
4QvXhAGlxtrocWsKkTOUyVm1hRTiCim6bUVnyUFqA4nr/6osmVt+Qfz95KmJVN5nIhPuul6gm7G1
m1aDhuW4pOeVcP7OGkoI+AVWIsvzZ6Eqd4DA0ZHN9X81qEZq5kRVqQKFHyajEr3TsangQNAHdWM/
6rwlHqUXe+qsihgVjc/e5pU7uNfAnb7VThVkXsyS3Zj+ypmIF1CpWqCKtPs0LJkHb7bK7X1j/6jk
9pDXgvuFMaKKKZgVZlACAODB+KsSRBzEcdbkja/gUzOVoH2VqOWP3SpgfzHWHyetI8kuHyBedIFz
ltLmElimQIOP3Fuq0TNQaaKjgrnAzdqMG/oXTzZMeo9BcAY3wtyEqMRb8Tl2fndy3gebSFj8aQu0
Wcu9nXgt4fLGNK+HEyF7Am0utyN7Imd5BAUhUYdh/FP9pIJeSjdLw64VElqHOxrhaH2cRF/U6Jz5
RKlrdFKr9nOXzzvVgCVpsXWfnwosFPmmVqfY971xPC+NK1g4ohm+byulmDp6Wab1BKUCLArF3Kxu
Qtc9krh2RxEJWVnrn8KZabPwU3kpH6xEQQ8sqt6u3YPffJB4CTlpSFwOVujpzZP4NnXUqsXu6UxB
l57FBihJiyRLw4r0d55fyy4KmaKlwFG1r4kepAmpzpOjZLLaZm2hjmqAMEBOp2SVI58lbENnw3d8
HqT9BmOXJk8sx5bR/b3qbD0ifk6KO0UcHWLOius/OQx/fuVhJ6Rq6Ms2t4qNVJfDEFqh1oinLECx
e9e70/rqdoyEDRIoNJfvS6El+pl1E4vlrxtKd+1ae9qo4F6iesqBBPZ09yo/A+FyRY/N9eQlrvjA
zLYXew6D9zQiHZ+ecgB6dyE3vRMT3wQYaQKqgb1+xg/8pfpIM7F4Umbc1IH+xsmmVLE1PfOg0gX0
GT9uRSIbZOPNEQZPMdlB91Pl/A9E/tLssWMEXn/i9TnHsEahLN4uG6cZNRdViPgzi9a0swdBb6hX
IzijipxFu2cvHYwdQf6P1oIxrDasFKLS0ruNRA8B67p2cIQkd6pxLvKlVylLzIxuYFcu9mbW1lbM
t54I0PjfTDYkRHehw62hto4Cy8p1h5OTKq6ffdF0iR3+Ues78Z8BXR0u2toa+u7JfRhuejf4gTkF
SdovWSNnjMcr42VYe+1KxBsQU3yQeRZkoCq8uGnQ7DTAL4BRHUJTdRjtVd37oJOway7MuE4pJZr4
XUdFnja16jBfiFeb4qOKns/B8pvXcFk/3ZRg3rymMVOc7LRVuTyj/cppc391o3pBB2h7lxv/ZEsJ
1cvbywFfQsKVgdOyfKx8S4+GBW4D8tSDvR+AerrHQGcJ8VB0W+IbiX2zCIuVOiXeqTUtztSXjBJB
p00xl5QHEmQLAISSuEmqCrCQ7sCj8xjC/KiOPsESrve/XlGQR0F5jWYa5oIUX1GMWUayWyyQ6JfE
lTuDjCfd2jcnnhymdC5yu/B7SQmJXAYXTPn1gAXs6ph+QVTwo3gWgYOVtzsJQZHmMsn+/yM20RsE
zBvPW+cZp8KByEFyF064xul/EZfJhurCCRTWHrB6upLgX33JDdk6Dnf4GEKvll7zcIw+pdfqsoxy
q4lsprznJ6dDyqZu/khIEJjm40DWaVK3ZNl9cGckW+GFbl5WcpwXJ8ZMWzgnMg60yf2iPi2JqiMP
jJ0SjRvxzYs16EFhFh48QO4GCt+JZKtPJoiUsg8lLxwWYh+2KMAPb3ktT/Ll4T433S9XOzjg10GF
G3W0BSj1BHyF4cNvQz/nm2fPuXeKe5JdyZcKo2RWDasuViuz8IlJ/encumxnGn8ijyJmyLItPOG+
pyaLlElwRsbe/SmJ9ONPhPc/lpeddrpWpDUI4DZxhFTWv3mb9TIHrSuYpWU5ZSiakLjkLJKrsZsP
Ie/SqUesheosKum+R1YUfNPCzFg2rv5AcLpyxYA13F0g0+I1kfbQ6OKC7/DNu1z/dVFpBudDmB4C
WyrkfXC9Bj4X4lPh3j5khs0HjLqx6w+TUGfeVFW/qITvACig7TzFeDamkcLsHA/jxNN1Am3bO5jm
g9lKJS+RJ63QAZ2UnyP43JyhKrlnSAJJRtp6JTEsFBWLrU/7NArXgMHqc7Jf+Ljo8QGRaUHHaL46
1xm4eHCU0hN1ixcyb2dOQDRXJy+HGLynjyhk4b8QxUDF0+R+sudZNkP2tnfWiBxuWtXhvMG3zSRx
196qctQ2eZCaVXXaqW42sAkhtpsx54lveNn/HrAYtu3I4fSonBLEiOCCjk87r3sCApPJSA40abd4
B/XDDQUqeoZSCWmh/7ylklYdgDbqi11L2IETj02eXitAjNOnHz1Hnqcd9HBXrj1sdkJqsWYUb8j8
1ejoOxDDAfD4F7FX6rwH9HpHjE7tqaDo8cXNmIeYzNXDiE2cWrnuN97BZpM5/Qjp8+SToASUHo0R
lionLAurhlPE7yssq6aFUVOf6+oIXEHLg5GADJ0T4YUFdNZzzMpIV4p9/WHVWzli4dwuLVF6ljfX
k04e71YT2/uoqtSxXOLIr6U1J7NeTM3RIpmn7Q+9FT0guFKfv1KkPufzcUoBzNuBgzKe5tnRJpyd
GqYsD8if91GSFNqsiLBP6HuT84bXtNER+bIeGGgDVLlkR874BbcXihpF0s/vaW5ZXg1BRDrVruDy
n4/zT5GHA7nU3+vukO+jZFrgEs/DewKLwY+h47JOvp6ee+Ym8A9z3GQfFA3uKDmQcGE+J+v3MgEj
+9S2sXBtt+wmwQXCg2PUmOYw/AmXl0n5DOxMdB9FEZuYlt9vaLE1Z5eyd4XovgrgdBv45626yTpm
hwkxRwWDP1jbp+NuEB+CpGJgU2o5mxdRHZCcjefic9FPV3FTQfERNj20zEfT+bXdolhtPH+Jhd9Q
wev7QbZ3SGv8D63UU63rRMfOgEvFD4IbLeN5a7UWEEJdaZ8zFPrElZdUNvs5DK/r9ohgJI9kQoX8
q6G4JB7dSORF44BvV0rAvf+0CfTcS24GmpaevD9XlIInmEIG7fmWSGvrYiSNS4zcAD/A+cYaUTt8
i0kDLEIS+p+nG8VVINB+q2tn+Mrx1hI7y2iLMKOEn17aaVZe72WWFIjXOiTg5WGUrCgxlcPrWD/I
nZvr4Mu88hDcE25JdQsjv/0gb/LE+kRUNoJoMhIEVXN8lQLvLajdcTZ884cWhpFgCRYYXPwN6+eC
jsMlQuflrdJFI54EdLwZ79i1/oFQ5h45bpf5abDj+FuLK/t5cXgkbRChxgEm0Kws88UN+WcpRwxw
qPfzrZo/CZbZD5TJJlyu9gMWJls0rvEONvJrK2yb03xsn+0IvDQIIgNfNtaA/lG9deZjo3qOFUG5
iIzGbHzE/aDM5pc8/T12aVs4IlI8wp6WrGP40OWEoEJFAjJ02l50gD8++G74sY8TgvG7JnsD+vyu
IHOf4uU7KIlWs/1xPcn2anWasUyAqGW8O94iqPmZvpv+iK4EwcEsFwJErVuImpRYDl0uhgfhot8C
gAYfRHTN7auK4ZaaTergC+RwJq8r1XEB91ORne0kLrJutikPCo/Cgy/Jf7Tw5C/n2w5drYAjqBn7
2FxhkKIPO2g4Dd4RNWy67wSajg6lsdkG5Mzm5q30Fvo+Y/iEoCpaCn3jq7FBeN6wy5HL6BSy8Mmu
QaonGo85px5y0Nj9eYFJcgqrGstkCN8a4ezABGABT78gWYEPRb26RE/NZI2bSYfJeMk4CzH6Jn60
VoUL0zeyEW85/IOllG1rDJJjZgq1aJyQ5LIA7fxHYNECjWTDJVr9g4uFf6AoOFtRTB5GvcDjmrTF
wU2pBnC2+L4gA3HEuRrvm4KlIUPH5osbwEyA2hbinWiw+aNuLG3bRj+csz7PvkBa8hn+mnVAIh9t
czNCXvmdKz4/X7DQsHVT58O04rREggbsQa2pwZfA+R21P7KHuJBhD5c0HeF6bUMWeBfk0MANp0tM
woqrT6kaOvi/ohsQba6WpmX9zIaL3r0paNENcuauv1Bsd/zG/8FNISoED1WhqgKiX0BgCmB5pJry
/wWo+Wcwr+fKlZFvRGdhjeE+53qdRMv2E8Ted3pYTf8SnB4Gm7UGottPgrtYcri+Zqum4twjiRIB
i41UFZfCjlF5bTkhlSmZRvp+qndBIS21aIsqEhXdMsmS/UHwDoW3dfmtS9hEp/U1nh8LtthC6nfT
sw/YQe12oPYvDlICbKPmJxYUdQAzGDUCMJB72vEdDZ9VH0Isq/oXGb3NmJXfvU62waZ4beCJkWdf
a/aTIGLAb7bze41ZjN5ilc9QGBwnVsdzeuiUY3iY+gc7NLldYK+/REDvEEgubFEW2GCzf5C8lovP
+JU89tBguI75gLdUU5UDQe4lGPqeRISdOUQ2YQoxDKsbn39NmuPJhwIvFYLN71OTuL1SQT9o/0NA
mous8WEjkdhHGwhze01WPnZhzaJRCGx5lFTh1Fy0LT/fWG+EHGh2IDKDmekH2WOmiS+a0xSdelXD
KWfiqBljnPoZEQ9SXellN9XLcVYMhdv4tbOCwbIP7KwNF1X1xmXmWbw4B3KWpH7v29hGz3+R4M0T
KXMQUzEX3h2DaioxDF4njO4+0FXHlZRc5igTE3+BGKJfNVNYWvp31NjnTl0Jj9jMKDO52IdurCex
uHdGHSHAmx2ru2ZVa+HO0zbpIOV+nHYHFSKG9Zt266fp0MFBbU919DfYFWjjl5FCiAyrGNlePft0
rfaOU0PKnNOKxSRj6ficd7AWHgd6710n5xx197uVGiblQSIOrSods53ieX4gJDG8aqgL02Ti72Cu
ffBbs75wM50r+RsJBykGf0bj11erQr6VYtV516Vr3zs23tfS6RGXm9fLEHeY26A2AfAagNDuNfC6
Ag3W1RqXNu2rAG4YrTbq9uPt5g+FJuSSNnH/gsk2cQJooRZzIUfmh7yhQRbHuiqUmBee0ErMhdd4
0eQqfmXmXJTzDiTEgqb7U50fneF9z2YwgiUcSY+BBmNuAw9aiHbXchfnp+gru+qmWLiUCXq+MpGL
d+iiwZylv+9jKyPjGtgDJA7dixmhDALO1r9k1lpZMKJMQFVuPrE4n2fzLvusMqScwY+uoIQrT10N
7sHl/ZWUt0nQ6L3zHNwYMLWDO0Q87gMm4MWagrVE/UhrSZmHKVOmS0U8m8OY3O+7ucNttYSi/uk7
0ben4GBoyxuGaiA1nes9skbM4TMiTyTaytL5LUwD3L0BBXXsDFzUq+USnoQqVP5fTWZ7p+u0Ify3
N3Bcb4jnlRuGeD+3id0UuOOmvOdCJA03CBQ8OOPqzheW03Tf1gluneY52DxW95dCAgXfXbsNH7kW
719kBd+A78xGMgX7rVx8WuJKieAb7qxFDfTja8cO3Hr6ZYR01ZvwqU9wxVRjrmiQ5J1tR73d3dL5
x4tY+vrnBzFSI5nqDi5QU5IEk/+eA4WQGMcdS3fFSncVUnTTYqkKM5hpaU5ZmraYQGzmvMLJhaIS
NTJf5istSJkQKvTA4BnUBm68HCumP9umcn/8KSyBMr0YQd/TtGpIOoi4J/LvUReNtsz2k14F3VkX
SPruT56jsKyckieCUWn2JMjA7FmndkrbvWE6gH3lXr1hgYmU3jmUXhgICuwrS4JR8rW/2RUxbhvn
xuXPlOyRevLYVtAysao9bLOILMm6VUyuJwpPEIC6gW2QzQl1vHgPglfA9mgluNmD9fGRgZ0eK3Zm
Wv5mj6z+mZbcz0/dW4aFgPpbuv8VPCqScW+P/La7eZebkyGD5EUTFO1fdsP9pDb975U4h0eG5/2t
OlEXm4F25ya+zPVMGf0+DDPrIE5LFyHwoKNpktFs5ka3IpQKM5ndS3MWc2QCGh7HFCTyTb6QXaOy
U8C2UloMrL+KDYDRaIjbob7f0GsZy373wgqdu1kE8gWimTy47yZ09RKKWlnDvo7fDnAHudc69shl
jTL2G0ndtE7JAHTDM5nHB53MmETOkSZaMVxGGxmsSZq3f45mjtlhG4x5b8KGR1ctZ8PU+UHIwIEL
Oydc7oMA3E5nglkTF8jHFDBeDyW7O1N7gnV9FQin/iNnkkF77yMAIYDMpNtmCDTA3+Qxs/COFbc4
oQ4Roby1jBd5WZkF82YCXYulf15Qw+3ZBsbZKMLEt6+q1cEv52ayHHG4paQtC9NqT9KJPay2jstu
yyUmOUbE92bf3GYbNlDXWv3qPewg5Oj6efHKuEknrwR9aYhgDiWfmhixMKh7HCKRAzZ4j1ul0ONv
kR99keV/vm+7mQDA6EeYXKQSet0J48EXL0tko94+uqajnwLuTjgJ/lggMFrNUBLVGlVTjRFpFv20
xeFOKo5HDAOi4Sxqcx1mA7L20xgYMAlgAJTNHU6ZZbcaYHsX/VGKUmZcar/wxVZm5Dx6zS92e/P5
A4Twc6yj1rNsPnfnUIU82ZpPmPCywfi39GYvMgey69n6alzC+2ZFvrBcutmJDz6MxakPREolPln3
/LFe007umFgptsk88f8xgqgz8pkggmsBMWtqjW4684EhcbiExS0laG13ecy/cKuhKXiTgpdWXpVo
5eUMnn90uGoiGKUE4EWE+o+oqfZ4OO3c8uNGcagG0zSj9Wd3IQS6jmUiSWbpWooKXBpkrmn/lJwK
mmAqLOEXTn8U5Dp8yWkInki+P9tM0nmDBX8rPhySNsHlok2EGfqjqxEvSDuFN19YGZ9Ame61hsuU
9ncN+xezCxRWAJRBacHlYkDR9xT08ktOoLBG9pRxg8Uh6X4WSSzHc5/utAsPwJfaYnOBPnf/X3hh
840KipUAQH4SZHWA6PGAABayAgIAbK6jtFjjcx47iWdQae2EExkWdunsiGTRCHoxxuQQkx9ClFoQ
4+n5SRxUqopQ5CpptjGgPWcBpFkkf4Pwg+ftx0MpHn83Lrrn6wCGdn2GyWFu1p9QyP2m3TL5ITzb
kMY1WQTjmLHKBonOuPAQTQPTbU+Tl+BWrqIHFK4+1q5BFdt5NdU2KiuImGUTQx2httIYy6ouj7cq
5oM4XQZxTxQ3IkgSxYbKuegjL5pSBR+hsoO+49CrIRwc8gLcXwXhdSSlprTCKfES/pzE5apBm2Rg
D+mXczezXoOfWmPk4Z7N6NIP806fCxRhSl+0TlxdN85dgomR4SZ3EU2N+9ELbrlYkOP1KRQJKTeC
ygk7yu57pZU+Rjz9sTrCavDtlmWVrN/3Uj7j0EXIYodunMM4ntiBRRW8OAAQjxMt7sJxIag1Zu7B
othxaPgVA8Nueow7nUQstG8As2w71b8W4us4/1/N1Boai4V7KtjKcmfIMay6JKCDjKI6UdRuYw1I
++4htVbVYxhoBw9vh8WhK+Nau2PpN2wcsvWKR6sKVe3w5VzMjOS0E3lgtxAshd/fN/n1uuVoPxZK
P2l3SMs0+xgg5uBnTumSuBxmOT2W8fsXEPt6IvXA4rHeHgJMqFXPGAx0MGoY6UVQ3njmzTvvYppE
e1YUtjr/ukHZd5Q/wnCG1xToysBUIOm+STc+An/q6RRVNKcrBMGLBqmOFZFYV/SIW1H2A3B4sM+n
gCErAB5szo8hpi+RIxdAC2YA2GmFgQ7Bm/5tTBVKvsXRj01kziCfmC4aC96ENu1uTWVXWPw8Av1M
ninmcl+7K0OZYUJnp0/9UPEwSIXFdRH2+vNpSVgr+I7f51aXotE5nrsKwcFa5bn02HA1AaMDxf4Z
n7Ji/iwQNP4wjGeorqT8cJG+PYm9mqtz7XI7DPk2oVARtbZitz7rdwruq8IJCWvCcWAchOY0rPif
5TrGP0t6+0jKzIi9A+7MD23ra+R+Vo2+40rEb+bZXMl716Dsd79eY56x6radbax92qTfMxHGHKpB
pcXggocHFw7j6IgtyzKZSAe71Tr2/zu7XI4+sEk7o6Bbg5S5Jrs50h9ofHW0CJmGgHEbTPQUxsCG
UUOMwmEc3m3azFfY5cNBhVvviVlWYF/+AQSH70nSLDOYrDRdhAKXfZ0sxpt39ctNZaRanaExASZa
mY045lhKREfOxigfMUFhjRQNkJMN1/R8K39pQfNXFiHHlZdkvpkJHmax/AhQnF3UZtyhCgLP6RxU
ISu9hNmJ7xqNJjGCE4vQfbVm8AsjhuYk0mCf/7j+CvtFjBfGfTsdg9zON4AEJqNRaYApH08HsjwP
Nkl7nkbjgLJfumlio9bka7+i9dBBanelZP+zgBAZVd1+5tzbUf6rbqpmKlAx0JhFJEWz8sFfB32N
9JnvKhNynD15ag/zHHDFWITvrp/66I8/VB1AjvquLH3ZyBqG3ZPaylHoEhb7KMfIgJZvTw8qEcBX
LJM09ZD4ca1bUIKf6zjW/zfpV2TRzzmOderpB4ptSGglXYSFKzOqiRSuHOSx+SZaFDhC26HRVKuW
sD6aimGTkzh+iicHUOx/TCyBnp8Cf321xEiBDmexudPkPcLYdI0fp8uXa+++sf8N1nRpSh22ftpk
BNvFVXrCg9XLmaRKDRxfzuTV1yH6G8N8xnFNsNnAMWLFlkGLcmVP6VsakjF+6IbqVp8/s61iuVDi
dNbEcYuemM7VSCJatw7/dUXCYzA9p2AfgN8OU145nlbOeLlW2mCsQYr01EIas5TYqOeofuuMMTv2
ToJyPUNTx676a2tjmfozlVB7oqBDDBmNcQgcJ1rCeKeewLipQHUEYMf62aGce/kUIhxA/+kyXkhR
GiRo7PkiNrOMU55lCf2VgRrA4eyz4M3nVmhAQNw40XPQFcMeD/56xRYb78CVwsSgg38X9Z6QNq55
YtP4xQECaO7KFhs41dQMvVhJRCroXmrOdN449PqjJ230jZwmJLZE1ERHfokzuJVxceClA9dbI4ov
pB1m87R+lgrJbyrqa+7I4VOKVvw3j+14Aqy9UlhAv9rrlmI0EFmtKvWrcvOFvUFFrqDSg/U1ywns
Q+DxlZdJSeoQsL2y1vCeXHBDiYbDZGKAms26RqZBNpDEuCchM6hbMphiPWBYqbS+7jZl1X+AzEzi
eZqyQHL3i0SMYlyt7uOpFftW36hWU963K499Cthrfnn5qY1H4a72M40YPvpIORD2cWD5itsGfQcX
RSCx3eH/l+gbRNQekNK3lQUHzKqZapkz7+KQT5GJXPdGPIexBfAGW+4PTdo7UzR5NapXf/PZiSYm
hzP/lHLm0PT17HpxnZxmPcpa+iewnF0itrBBKfM6D65TnTEin8xrZwl+3BYKupgemjQyD2aBjmGO
8nUV/Veht/zEC4aa2KQmSbVwmJCYy3UUL2tojBhmuw6J6Ar9H2MdubqROMtg0Y9nCucRxTCWkTVa
IGIX51clWjYsi6Qmc24he8P+gljDMdk8pqbHKqjS3iVu0ui3yle2ti8vHtYs8DhIrqFapVpALu5T
H0rd5ELJkhsICf0vVtDbS88VtrKX/BD5xnnbuegpGqoOp0eazQFdoESOFLobk6t9id7aYRijANom
EmbHDmWwvZxy3trQzSKC+gf+/KEr6ldktN550CW6CpfU7vEUDxpWwj0taj6TtOut2ojH2m4b+0HS
tTDplR1EWC2sRt+M/qsiavEIc2GyUnJY5wHb7Kx1J7f+0RALAyYEBSf+xpMYhWXKDIBgBTVJrs0v
cQDzqiVR+4dJCGCPVF5HCRqOoobOeBDZ2qfcSwldY69h2pZPpmNMITKQEhpYAEguX3hog1vnbMP6
VyrAkFqqtWnfPdY6ZP+W1s8i60PCHKfOEWjNzUEh+6VF8GFHrdOfNABi70/y6eno70MSNqzVMH1B
QTXD/y7Xk06nHzWdmckfDrMS/N0thkAtwbmpIMY7K+XHP8JMc7+btrI7AzYRxv0C71II8b6rw/so
GmPIi5DrtXquIKMPx106PjsKGK8n6ITe79kWgyQTli+gV+kP4Ai3yVh1s0ZsA7QL5efg3EGpRnY0
pGO2i+Yh7q0dtIwOZPq1Gz7+041IDV2mizBVPQAdx5yWy2i/eaIfVqPYngpPjtiXKS5Gilbzh/PV
w8Odl0NuVN8zEcSbFsR9/dzqHXtZfZjV9jK+QQQSeo0Pdo5u1q52Jk0U79WUrXB748+Lw/hbzwjR
k0wPh2pQ1TqEqjiY0gnFijPgxVIZcUx3IZld8kZiPYmjmuT1/H4CD/6x2BXXvk8cIWc98ZWqRaJs
KnyF3NOtt1vasw3mti0LHEUslHriA86+azW8R/pPM5NjdEnuAFaRTlj5S012/POOI4YOfFd2v2v9
HRvhUADCSCFBmgfIx6RF/deAf+uc3sFAwnsok3xb3GeB0uBDa36ClIrgDoouOsA7xcR0ME0emU2H
ecxdW+C1rppXPvrcDVPbsJH2W4/iz4hlxbxwlsSaexuykVQ95qMLH3V6asngk5n27trfcntUU25C
07zz6McnH7SRQMTy3dRro2WRVcFCXz8TiEwFQDCmAvcX7y0uHlr9HQE2yvrsBPDOGUaZn7nWONAL
39lGuPCMchXtxTCmDpf0wAeWCwx3j2HJeZX/VWnHd0BQ4Nr+fXv7NopmXUWxEoPQDbN3OOwsoock
MNP3DjJa8EGhMT6+gSPkXa4pxAtqNVu2NCnQ0fek0SRQbxBNPfdNPkd8H13tDyzf+WUGmqfiHqmf
IamMiZnlgH+I+nLSx/TxDcRk8X9VwiAwC0A6Ns5k+fzb65cxkPn8a2XMn7GrDVI7qShXnP6pB1fK
04AvY8x2SHgPvSpe2b9awq6rNIRbY2w2zSr3iscgHbpHw96MFxJ/5NZz/0BGFAZKFIlcmsICRzgm
KER2UC7g3AZnBWct3j2uEQKXFGJ5dXk6Majm/vd2sNI71H1kepqNcLxuKSr1gW/URtJC/R82GtM4
unvJegnXK3cWE2QVMSLx4HdFB5L15qzBIbnSrwOhw134dc6T5jmkBVtAlPAasS3VkUwJUXnbyXZc
Rat8swq2gPq8WthsHounXzl30sry9swJBzqV/iZYxIZBxN/ZNEAvsYRCdqBAdFHh20J3rQfY7MRc
Bg2HERt6dkxHD2OE7vUvOp4ZYmWP6AertYqEg61QDj53KNF/ihJYNgIOnzOqzwgxpYqH4+ZLF5o+
Sdqce1uIFKmEYpA09NXMYXSQOH3weBwgqJJcJIxKXgd2fCu6o4Syt96Ykapk8oHHyfKfe3w6PLaE
cGkl0vLobZRoyCP3pypufIXEIaKW+pHvK6KC6S63Aeb6FEHNIBtoD1/h6fmqZY9GfFovkW1AsVKz
3QRZwAC+Mk/4lMzwRz97d4xMvtRIYyEXBf/uRwclf6e6UfhqJ/wNB7Hqem8ErFngWkKKBRaLxJMe
LvT4Ir7PZ+3V1mSFeYHcLlMVbQOMeYhOn5rxD+w09QHLM53/Y3lhWu4YfsQfJ7VMhgd/AOX9f12V
P98MPh483i4CtuvM51coDJbzs48mbcF0IOgWiJWAtLcjTlPmfV+PhCAA/xJRZAftEFoh6vdfpiXO
7VaJULTt7GXyXyltjvDKxWbkjv8Xq/lREvNqXa/Dvuw7ypOmEdWKP2dUxFUkb2ZtXAjWL90f07EQ
h6nQDOtNzcsGl7ACzGqwYM1spIQwRUJIc3laqZoBFUwNx1xFlQEOSu3bVqoMK8zKtqxH9o5qgPYn
fqiFaMn2ZHR89WCNDEmCGFUAc+a46kLj5N8PJ3kllBI855C1elL1Li3jm30cRM7Z4PoAEn5t32vB
mFZm6/gRwRjb6xaBJZnyd+OdbV3Fz9o54OWzE2NsoVUM28Bq81SrhSHeNJLzLKyOPrO7CNBSSwDQ
2qnQi9asOMDE5zowreQ0XnFLGMaQKoh1vZVG5k3n8SHc8XfT5sR8BJ7hHU5cQXeapXji8tuxJYo1
0QqejONqDLJvBELJhr6ILIMoJGrCuYe3lOPO37gKoBAY5zPacrushhYiYLEqfBgDMkV7nf1CYnbV
fEWGVn4pg5+NU4J5d8bsUa4Bs5VuWcVLNhLVJuOJ7cQXrsket1TpDOHiZKKml3wMNXQMwjkiAl2p
dmvuISGYbYZBFvy1eBFszbN9biGw1zYb9aoHEAP26i+AtnBjTlwX0tIgqgmAy8oaHRUSnOEI3Wg/
W2f5xKIGHnFdLDHYxD9p8izHmxa4LdCtNNjfYh9B0Y10qC17EbS78CxlR1uzg64bWdjgy2JFmLQm
Z9uiCilU6bbbhWTXnLjiXmS20VGXiWQOYsxbe6kciaVeViCWo/FLMhQ45Njq0N2zdBBbgCDQNWuA
KY7ZSEKp5jotGp40GANzi9MGQD4fuKiZS30CMJjahFT277BzAkwn/itMuzkuuHF97IVCXAK+ujZg
TiacfHr7cb6JwoLXFw8e/qWcvMnZMiilwdrCWGXh7jngvMl6C9yxSWOqa0EhZ0b4xO6DKfhQ1r7M
O8KW1n2Gwv25sRXiL4HJhwrg2sjBgmdLmHavV6Sz8tg7gYmYtBGct9QY9NY+EuERx55yRqBog/OS
xLj7UUJKiK+faeTeL62OGQPv6NmYZDc9EH1k0YhWvWoQVrN/SBGRLIxTGlcrgTJYGW/np+2akdeT
I4ny66IfdBmz9LmSH2+dFre2WmTi8AAwApHD8i4CQKzKEFBwNnM184511irDx+9X8h59Eza5ltO1
RrAUpr5DVlbIYvw17rV4jFn75ZI6ErIuu0fiTfmBUaywotQnwlq32lt8X7gZAm40rPytorwoyrAb
X8mlNZFsQ3IWnB+/1TgHdQ3Q6GjARk8DEgme8Mlambs+eetL+E1EIUnKJ2pzkSrOUVQZpWWerHrv
Djp6xHP+hEYQxdJyCz527JNirNxieY/tacbTbGIYLs9MHk0inIas4uS4NUQN2cD8BgDy70LpHY6w
mewpaW3Ol4eC1kPfb5XhNhHS7ktLe+oF3QxSxAF0lmh7O3o4IGmPVAEJ+4YuNY7Zce5PNhkXsNo9
NNr7vR5Np+p7cCFYo9pEBOGbqYNQOqULj+uA36likRDgn6pGazTb8VxTrqbyjZVuL9AqaAGFeFB3
Z/tBScVupAkvdGk8v+UIXl9siIOV6MbC97r9FRoCSgPWP7uBoI3IqhFg1JFLlcswjbjPrwFxp+3q
Qz6/Fq/ueHQpE3mbCyK5vshppDO6huShaFyBbuAMETl2ftnqfigcggalDgTvy5eJkqqmc/nSen/Y
rfclienBh7+aVZPf+hguqgooj+G/VkAoQjmTZ8lASPeC5IJIKZyDJgwO2XhmAsUsTQqim+PsdwKk
Jn8WAQ8D/jExxmvuizCD55SBD6tQ1YbOXOsF0RNbKgYVKL2JdniGJ1mlK6aDbDWPKof0Vqr3WMK4
HRJrxg8IhQwCqTqoIn6nBVuEuoRJ+dkvvfRpMQ0fqj2rjlY70z8P/R6AxhuulIpqqgHPph+efmPn
0SskrnVEkgKWZrA5egCfNRq6drN6FNTriYFMkpczIB+Nv+CNt/81FLxPt0k0YoKMrZOKCdsuhHCG
kFp2rK3GbpcG4kCa/whq8penFpQg4l+Hq6vZVzgB2lpo/D8ZFTeYRZPJZ+kpqOnzM/bQOe+re2kW
0ymRCMJERVq0dc8I99aAQ5gIKZZpb5eZceIV/SlEFKmdjvf+UpbQ04Q8wSK21IJf8eJsZZ3IERJ0
CzWDAAGDPkZMednojjUWjj9jqE/gVo8uH1j0BHLc5UnTezfpUocFNwfjtJ99WHvlVaqnKK6YCFGG
8iDnz0yVRUxNwuPv9rz7jmRC46wyv5Nksp3tVbLQvUSnkIAMxvJ9pKpmOyn8gwuG+s4Xk7NtmqnE
JwHe7NCgJEZqstZsTcv9Pig96PhFfoIxNBj4WtoMCV96TYxMikxSdK86Tv0IbaOgwCq333e480F5
zOiKrBPK1MzMltgiGgCMbj+ci4TkILlDBv93H7KftrrT/eYADHWz/3OcH/xhoSyX3WbXvpGdmXSo
8pt09vii1eN9DnQyXKc2hQsWnDkaM7ML967rDlqnoKNvWbUWlvCUtkqAwtSIROAKrQz6jxJ1GwxB
0oTMIYUC+9+mDVCkdO8Pe+wWwESmjYjsPL0bT0BxyFEetbZ8874AB+aVVi8A0EJZfOwiDcEKCU2u
WULKklOvK6UKLa5EXAtE0j0QPDPCvY3sjSLlXyttJN1SF1JjySDta8OF8r1A4x7MzyP7JVURl3s7
6ojDqPFanHgXWOLBwGjGz0UNtFi9uFoVSZbWA71yJPIEOxgtxdXJzj6Rh3u2dAeoXZX1jO/VI+bP
Z76Y7r2tXSZ9iZWIBMwYgvYWfqifkHHVDd0XRlNw6u8aTb2lDLoEpfy2TL36C89/S5uWKh6TC5FK
xNWd4wf3mZblW7FRYYTt2gUQAcAqKPL/g2mPafarxnxut8MhpZeVJjqF65gh4bvp1UJmsBV8FVTn
sJDTVTCjdtTtttUz58IhlWtXieXp/ItO3srVTZvn0puI48cRk5X2hb9fgp/tUH/dt5TZd39m7AK3
+A1ZL4k8iL/1JiZBgA+8uXfPjXPbEWT5//PDGcFYOBv23ZRFUX+7Tr0A0kONqv8y7E/aONS2S+38
NS9+Pyam3Jhq4++AltaLVgULBON4PcHpWpyAnIj8qFeL39d9oDhtw1uf80iJlaUfIOswpvxMCNAs
12U2ZLs88XhM9P0LAPFxEvROejP4mUtFJvayGvAv7OuUJA/V+3SDIhdEPDagn1uRcgzPQfuSwOw6
jUbQMg7omGPYgz1ZveJcfJHBlSDBEgEhc+/QQL8HJcFIzKM6nYwXiFEtjN55uxXeWDAtot0avUIc
XgP0e0NpCLXZPvrdiwi0MSrrqcGIuyENEL7igYEV5vuwJewMFUSntLsIlKNKJ727lvNcRKczHZ9s
LJ83hydLn6HV5HGg7eZt9TNZE7Qhh1c5eGjCp7OwmBnvFhqBTOcvOrQdkiGkLkBV0dKaOuoKr1j9
jxw1Dq5RIac0TXoN/SdfsM6OpZKozuf9A6dzIcWXXtx34kaKLoox360WsNTfkanlGgWT1dCyGlHb
guYf2LtXoEANkW7GO/XRP5HJVzmXuFUThZdtC2DSsebBO6owi3YZX9i6CN7+1J+urcEeHqTQ5O7x
gRtCMB+lY9Y2yXH5lVy+nsGKY69fcY65GCzTQkKeVQAtYeGCSol3ttFfv2o2rm3Jj7RxpjzCibbs
oS615BijT8PWob6NXbaYS91r23i9pw/vT9jDN2ifetgdoxWMyrNNtIClXI3KKZws34nV/qEXjAzR
DzsXN/ajMBhn7vM4FjJswUmuT2Hf75OASArujX2NTr50MNb0QD+XXvYn+gCZ2ZP7ZBUPqWL+WVXR
tt+Y0Q9kC97DejK4Jcu7Tfh6DVMycC1r9NcVad07QMtPPcMv6q0pHYwF+I3sm4AQAL3ektAHF0+5
q+5hWQXJRe1/IrxSmpTLQZybal1So2J+L5PyfC8HYBJC+l0E3ZE9dVYOumxvGQv8/f1x0blZZ6HK
++5sBPFNcegF57k1KosKBpNE5+siswvgXaJyQcVmw75HfwtAtBQFvx7B3ULjFhqNw41O8VfqKHMf
GOkJLYMs0jthma/2DjWCVCnno5qcPYOyEVfETQ/LtRZx1uHfwvF8/xinVpoXznJyOa3/I+0NkdED
EWBiPiWz/UFzBLsg0ZoRBvp/7ouRugcOMuZ93NHLileD/AZQfhaebxGRs6qbBRCR1880VV0KRCf8
B8YnDrErEp/VhloOhJnQD3oXaHpcMFpiD0lmNar965g6cRO6uLQ1aPMi0DTxCxFN9OLYVRYej9m1
a5Oz5wAG93vI8c/zDc3/nRQ02JKfE0QSBY3RXX4VLWaMxKvSDsrPIEWn5zpwywGp768hBxgEmdRK
G/wSQsfCFRQgMHorbAj+osse6/OmUadGFCf3ybmSr7Bj9eOzU619e+A1XKMa6jhUMm0BijWbWrff
zZcZaIxtQ1p0bk8rNkUNXERSnpjYsgnzDDX01z1N3G76IjWQJiexG7gCmsTcZa39RC2wVZRjC2uM
P3W1UCCYp1MfkcWbk4WxxM589k65hB8nKh/k5ZTUHsKZm0JDTCw7tpDRMCxXOwt+oTe1Zh2y0oS3
R4R2EQVjkK3HKbsnSf49xXxvDMBd5i/NhrW3MC+DZxyZ5ropRKxzjXIfAS2DXKLsWgtsgcC4MUHZ
m4ZEO87q2B3oyu8W+yG7YORQ8C75XqmADHpdShAxqU20ktp9sDAbgMvE964s7201duc3e4utTxHa
9aIMWo6Q0GWtMnMpQth2xlgJPEd7wuzzTlUnNRWVrpbkwlfUpLF4kMNJgEKz0c7sVwdDxF8WWYDS
7xZS5etJ92bVdqvvk0RFbRTRHXKv1qQNRXK1WIqIMGitd6THbaVvybZSCROq08h/6yhWWHXhpmUr
7byMrSI0yDVyFVAbI3z6RejiAuRTdzAiXMQh4/lUT1/9joLmTN6FXBEJnRSGO9heP1e/JDmmQB0s
dG0iD+z/oO2QSL3b0MZr8oaB2aStQIw+wIjVzzVoJ0blyLaZO+JSzHlg1d7PLFgV4h/2r6p9xsBI
W03GmUL4t0tTUdmWvpAcwQssL9c8XIiFTU6a9cn7Lw6ZAo3egQUIH+dekvK8JkP5moi8IHczE+Xx
bur4iji6fvEuNzYgUECnOiDQyiSBs+z4vP9hw3WpxCS+HPD+f5JSuXr1J0moI+fPikZpQNr7dddU
K8fa1IjSZZh+Z/hX8LLSIqIwOP2xEr34BPHGLC0mY5w91iSB/D2wWwI1FTJxfuoSObXoOyezJj9n
1SmQpZlZ/iCwtfpKeQjtltab9zmrd4BBMXkLpaBsCdN3eV2C56nSM///jDk3FAyY0LbPj1um/sRw
mDR9Lp6RaLDB75EqMzW0HkBn1U8dLtJegvKlPzeE2ct8b5WhTvS/A56kEgQ5ZTevzKw4b/tzbDzT
KDHSRlQBwsC7QH/LLXJOf+wYm2mhg0YlsgCzTjzJ7TTVWK1CHEcw3r/lgNzFM/kFeH+gTYJidsYQ
NRde8sbk2unVooUzosXsVemi8A4E6AQM8cnii1inczbSjlKPxNjofc/pe0Loeb1vATx3t22Cq+sf
rNGwn9Zn68sMzm3To07K2nBHlcIZKyiNTKY983F4ovempLFVtF+jOw4OMHe2ssxEYPGPoHXxXWS/
yTxEdJm+klNrMnKXQFn8tSKIBY7YNrtwJDzWuhtB0vWH8F8S+JMTJiuhUsmmLTLs7vhKiu4AjBgw
04Bfwa7vi5zlhU8fLytOi+3Pi4jdeGTPGMcjHNMhn2M6Lb37IW8KiKjUvBvY9FVf0qqSnd8ciJ8G
LXuqMdGkk5VYuDeSAgkbRp9YH3vtXB5fU7BAmRaWrWh4HFQwd0vPe2ozygCFA/yMkHStEhF/7+NC
Y8nUXksDuZl2+KQgObgiC5WKVED59doY1HoAR/CMshnv/VxSYfgihLjjuVJBWuJ2xjqk/rPnYffP
AaVn2kv0pdP1J3JKY3iI7BBPHFk+DaTZ/+WbHAjPeeS1rG/dGAOhfWnbZvom1b4+WPp6lcNl83bm
yI3tIDYIaUedwMomaV6una52JKSEBc6F7crC4Yl4ZM5gLfgDgzgSd9uRVFtB4plvVroVDUx9R3lm
oVo9moXRcOHSDXD0hDp3F4tZHNT3myiEsnevrnQXtMht6+G36oVWmAiuTyyg56RJOjb8hNrCd/cE
Ma6+EDZGGhq7NskMBX0tkls7v1qJju6FKFMcXWGd6djl/FxNVPYC2XxuVwBVau0iT0xb8Nc8Yfx0
xHzem+hSveGhH9+vbDqNNMHG2SPEPj9anJSPTEdP+gMxiD/M5dOqunSDzPv+zzdVHfR2eTWAAg9O
u7OVSDAEjQ+/SecDGdrwxGq0zhHD0zQfCevMWXaPoHZo3XisY7Q0CPrcviI3Dn91vG5rYJzKMK7A
RLciqtN3XxvMSRk/JSKkzDR+j5HywjkYz1rxaADOk9mM79243a7h9TH5wK22smp1Ux7rYXZwvLr8
avsR9SbNAtiZuyc0Keo4vi9i4Ozz0Ktx91f7X7U4SaXFDi8sMLrfZJ3i2wxAd9Q6ctXEdOgqiyYc
tl7MFn2yM9e1ovSf+yyCNa9U0ORcopostmz6UgUxbAZ9WEbG8DWWsgU98IpH/cPFFtlG+W2VSlxF
EQBdfCjCPOMfdxs/nWJpJxXd5Kr85cOMOMf97WYMMQTJ2osl3B8LMd4+C7nu4f5WIDvhM7n7hQ6C
3ok91lrL7ABmtI5eCaXNr7T3aknJYApTnlIYZ8uk8A5REEmLYGssE9UBWngYA6TtLLmtVd22CFf8
EdLUc1z1aGiW/ef4pLkVHzFoxKPTMGzFSuVJJcTLdUB3gciMr3rlTLqECY5vq/0nG4sqNBfIdqOf
WiJ4l+rIvXB2FcWshxYefhk28/+cFJFAs4w36fpxo989ZChA0r8+xBUP+NmSfVzIgPBDJLAxEThN
mvqoztsL4JPhI2dpeFklaOiF3dg1gpreGZ9058L2LVQKtpCsJtvNavG7ds+eZZbOCVBJAWG0K0hC
k8H8Kw3mqgP4/f5jEXoB2j2FHRSSDsXR6ljUANwjJ0NnuxIyTieKXNp1MrctC974GRQAR0qZ9q8R
YduBWs61GRHn9nLlD/yt7ORtFFZmMS7X0MnB1EhVKjv2ar6DkAsnt7LC8lG53J84XHOFhaYQi/kk
w4lgx9HxYp8JqLOq75rVXQDM1l9BYBFOa8LBDHTlsLZtCUDu5xddmbcpPCHqFqNjh69V34JNqMPr
Pye/1Waoh+Pn6uYQSgyitpQaguOcevtadd7Kzl2RzaL+DevFKOiAc4TAHMxW/dqUx84fZK7jD7WK
QhXqx2cOBOI5Oi52KLUPYOOyyuIxD+uN28GzBPIC/v30Bl32cn4mqd5QQY3WR/dFzMDfTZ17Bscb
kGEJB2UIyMzJ93iRwvC3JJIiQgfTJy9qj3ZWmT6Ren2blERCMTr4kCynsB8lFQUSLa+nbmojd/29
N1vZelWOSJXhY81OZ9Ob7lvp1tOEsP5kQqfCBQwwwGev05OhKbYUga21PwyLLewiHXMzBrnvqj8F
urgHNFNCPB7UorWwFjm4C8ZdffiHPFks1iEOIV07bsp3NqVaycrQdXHf+m1yffHu2UIE7CLORed9
Gi9Y9+FxSwQO5sWLO8FggwNFiZ1EawroFooSRT8gu/VHfoKwnphDYYlNwIfHU0q6uzCN96GJoaCg
4aBEAXw6VWiF3H4hx5vKs7yhDfPbIVSfPGRmVRXC3NUguMhgrseDGkO1zQgeSVWVlNv45maUmUNr
z9cAsTVNZMnbAn2b3lhraKjqIn+xwDECRaGvcqSOYrrUyWr/CqlgxWK8TwTSgGlktNsov9hSbL+R
VtkPsYAemkyuDnEA7gpkFqdtRfo1OMtqq4Jrc2pXbAMdU7X95fYtq81XxDriIL4erPL8e4KFBtxb
mE4E0qcYmgnBWYo8tLD50A0eDDb3qWBLEVqWPPsIew41lbOQ07INbUYnU7vzSFA+Fe05CTKIumx4
ldZZ2qqvvn/8UPkfx7MtNt5ToNGseA1YmlB/62whT3Mh5POIM45XFINnd2hzpmpB/0iuAIMUhOBu
wiR5+KC+fYUAUngVjuHc2YRM6VMe8rV6O/pMiJaVekq5k0C0gIB0pJanjNsOxa/ylod8EQTQ1oLz
EG5gJbEqkgFk8k1g7a46Buduyu3aWQBk5oaPdAzUaK7EHXG3xNe8Mae+KMXKNnOV7Ba9tlgvcmWX
sHbGaDLhkWk75sJx6MpLLiwOz8Sw1XM6VpyrwKjdukRQq5j40MHgo36d6MhOnhMdaxp8ajq5JOSm
PFT/m3sxaDdLvATxq+jfkfLmXxaXSJ7zZgpq4Z4euGdxlXHRJ4lYOGjih2C+L2mjPWPdkq1WUgOd
o7B9EwaNTjxBcPpsLqLuTnNLTPIvaVmZMI+37tvQSWDTZ9CbWNBQ8OuHpOSXYIVPn6E2BOney1UL
IdOACQduJgvD0H0WW2+cLPCioYyw9G69S0jYH+IZ1GApB0932ozjfM6Duu9hASJ6bOKY58Ddd70e
xUHMfOte3oId9ZWoXC19mqSMFnsAkoDFW7AM+2nSjM5Bmg+UDowETUkpvhoSV/6tgO9SP0XHkcdv
JRdXANYGvI1KyVfb03+lSa7tCQDl9KvRJh87xh4gSmx491IzCNziOXtlhllcbkYAwiwRTd8ZsLfp
nKluubYgPlnddmuUGvTeBJjPi9EdDK5PMUut/6FvgtaGWgO8RQgqbI+nSdLC1+QBwhvqxRHuXRPZ
5N2zr3mjo0vZSQATH6b0YhpnJ9xhZAiPsMn/tVlZcN60I0wV+Ngsc2M9bWIu03AJ7KzJI75wNiMJ
jTV8wPRsS98BQr7qk6F6hi67tLwYPFvNbuhtPX6me52uxQEOYo+zf/zxesf2HdaYbi0cXwlPo/JV
gJuMPecuo9bTav/KXd0ltpxdORvJKE11ilbiADDJJMzz2sBwN3iiWqh+xQjK+MGB+wEiyuTzgd9S
jIW43/RaiBYe2v+UYoS3XitkCddS7VtUUh6qOrI4JHzFW1bi5iwk0mrBYneYblVSg1dJkiJoQU3j
rZk1u+KZtxpKlXYyuMigcjAKOi1I8oiUE6zWPKr/BlVpIbeU5OjlVex4cyG6JJ6HPSgjvkP4vgAV
ctDh8RQjvPwi25Jls9ZB98na0zmIECBbL6TmZ0nIdgEPNhULyvrBhdpqr/X3FszolYStlCS+zd64
qDRNBmJHg6bXFzeWn1/CN1DWnVF7+zSNQ8C5Pg7hXJRSVxO4PF70fkyXCaPco5sT2/8VYYwzBp+b
1YYqiF15mZyvZkcak1MDZTkcOb1/4Q8uFgIqjInjRL/TzPkANIzV//ar0Cv+zd+3jJu4adiUfm49
zGithPQTg9fo8DZ0zWcH9ZKor74Gkk6VJT1tTJL32el4Wmi4pfFEb+wlSJouQj5N1TluAhcn4H/b
hIMJO/+bmPNA3l+eqUB8ZFYghknvH9zAVFu3jY/NI2cVlzbPZPkFmB9Ta9Gb8S0nocDcSu0uuoNo
AuGS/C6+JsKKaLg+F26chmX4f/kPL5OO+GSzP83+ws/D3G/PaiG/49pneTwzk0EpaQIMGiE8c69N
oKLFcvWdvWUP5gttAT/q7iuSBFJgwgDzIThopST42pLscpr3lYIw1gbY3EZuG8ij1h4IyAwWyx9/
fAXb1z+Y32BWd9WcnHQMWBXrNRBUSiml6QTIGPiHeqV0RNMtyeJ+NGC7hN3YwCg+kh52LBwWGv/V
1YQ9tN0W4lrjrcZn8P8gPkJqYzKZhOkPJi+0N5xzdMqNJBvwEjedWMqVVtbqy5VVebcT7Wvf5DJh
oEUijR1q9H/6sfOz2e2R4t+jVUf8stcKh+znJz5T78lS7ZueNjl993gt4dhcsQmDnDqO2Ar0oriw
biaSpqw994+rJ/O84c2wL20rDI2Dbiuwwhpw6TQR6WWdYeSYInBnEbdvDOJOwOgHpRXxVWEg8gZL
/Do1er7m+Nf/TlayLj7cr2lh1A0aw0ChgGd8bqokqbW1r1CaG/k57qdya4m6P18jM8njlHUVuZ9l
/gSI/qPn4RAlV8P1D1A5yPNMsED1KXzFXeUP/Q2yjHyacVrGHpK9fEzEV8/vrlGRHBv3g1Hw7byi
MdZTDmVGMSgAtfis9f79OJUdEB5UALXP+gOS3gydb6k3Wi6sUITS3gOdFvTb8iTvwf+lmKDyvHG3
r5Fd/ZPsCaxXmllSM4aWqTsnWxe49gN1G1ZYY6lh9QRUkZmDjLShteETUKdHMaOzi9ofPbbkmY4/
hSoUGlrt9Zm0jegSJvKOBcRAco4Bmm+ZOw4gERYFRhFDvm0tsMOXHqvsOkd/7ovL7NOA/xI+usdf
LuAaxlPGEuIbvan8n67JSVJoZrLq9iqkqhc89qNgYgaR2Ep9XGCquWpVNxJIgSxHaGGxW9vzhyQV
yg1bnaDsGsXjgx3DGzceEAhp9X/RVQrS1JIBvWsy7XAWuFH1a6sWWD/nmpI29ehEmyIGXQkmLucO
kOo87jgtYwSvdIRuNbKTsEhOnFFqD/2r58WGaF91eB2E1m9M63V34BEC5yv4g52c4UxL0noThRHS
WiVrn1h8WpDx/vGbITAKVTjS/8lBqFxDJbf9byqSCH4Wh3Vo2N/kQHGJ6tsp4Jx4PyCN4fgT5uzV
kTYes3mxNGViDHYnkW9Ix7pb3isG/smGIbZfSfHqLJ202JEuPAHCSZtfbitpwuLexUoACRZ894Sr
vjKJvbk2D1MtDVYys6SckIiyPvNnO235uSfIMyGQkTy26P+6PdTMML0/ZrmGUnUHPhGUdrMDvaAY
NXrZBFEZkfYzdwZWxTanz4D+hABwC30i24YJ4ZkvWPC6Sp5/B6JnrjB+8EUi5p2qkmX5aCWZqZQu
gtzBG4wlHYFrd1AbxI0/Y6SaRfqsJ78DEThJfL0VYJvuV7AA+0rxYiPbFdZfWz9zSR8JNe9vUc6E
I5iArRkFmsgK7tLjih/8YDq48KLHj1juNMa3kTcVlfe7J03+p/069Hptfb5yIt7rh42UlNwtiVb9
XX3Ux4x70VqAY8exbU4Z1k4iBfmrsdrJBLziznZQfBV/e5JremxlbTqkwq112xYRTv7Dg2CRzExi
vPcCvHpyqkTrav/aHlDCsQpfjKnQZWDqNvTFLy3HHIj8HfwX62WwqEwxogKxMMasCsrKilYsfMku
7MSAEjtNOMjFeeY55ZvAQFI5SRKC359vaxcbKHepLOXA8OBIp8zvNT/XQCEo8XOl5EVckHfdEGch
GJL5ic1zlZszeJKxBdjSxu9A+4GSEgn/UebyDDyDu2/QoB063JZ9f0Bws8cvO3v26BfGQdrBdEX4
2F31DmUk4EXz9HunfWT4eqq8BakAHxQnod8uaN8+Cgavt0kRi5nzt/yHwbVNH6TZQTtTp3UWAYor
LNfcL4svvv6n68sNBfVzDjKe+sAkYLaOclZkP3h7WuTTlJ+nbI9q1Ysv3YU1TL/u27MJXLqD+BRO
Ay57vknvtfLtyyGZG1nLKNCZBnbHXBOllRiESoH3hA2Xt983vwybZmzwgepL0lK96NEoLFdnwU3t
XmHYGhmEh/leAEULLr9vbq//iAyYiYbVtmRp0/gxLOlaJoxBUL7wWejcIhvlHE6/ChBW+F7QSYho
XxVrIsad71m5MSKqzJ1eXsH6+iuQ1t8UUCH7V3bs19YWLGGKI4SxMYBSK2XXPiGxSz4sUaVQN6r+
eJYDDHZtuLKX6ux9ixkHv+dmcWgNDbiUmbtQO2kfbacCla7hCwqqXyZuVxeh84JWywMzFtNziX4r
x0UmnpO+W5PzX3KMMcp5o4dsrAtcE8WM55sja4zbdJqwwPb1Oo+X++EWG97+2YfZ0ntVgJUkdUrX
1vBfXSasJasDBGai6TsDVCyYm3SZiz8yj+jR12zx3/cv8va5ugsGW5nvGgzXlIom5L1hW9bWh70v
/VsqpMtwo4IsWXXywPwFEfq29x+cMXuJ210592+gbCuBmKOFdsfpco/yzFSGIV4JNAhGWmnD2qIe
VwAt0wUY5O0UmLwpqBsKREazokDPAQsMFrOfzyCYFa5SOJzcIgz7LD0m5JOwKXpS5OdiSEe5OAYI
JDsiPL4P8j6s0MwQh7qs6WU0IKjMEA1b4K2ea82dmN6kJdcYnN7lt35dkI0FLa7tpb5ytB2mpSwT
j5SOH+obh3+278lB5kqZejL5OpjAsJw1CSRuCKqPEtxg/EuCPzknTj3MMW/71rowleYCpNyxfKMu
jxICm/juHInqlvg4G9jiXog3H7X785o3VT6TOAkJj6809ypwUadf7l04QG05k3Bn4XzUNp8v+id0
CxUsA8jiL4Y+k+F+S3sAnpXjgsDTDGuYgAwbM4uSQyEB1Hp+sVnjVuMe9NLuORJmvwz/TxBiUvln
oUum6ct/XitjdV4okzVL0iIdXAdAoN2iLYWYE91xAB3rBQQtNLFjpsZJOJqtih7ndo2PwJRlNVpq
56epVyI/bGN3wqeCM0cknZZn7sGgssW/9NKiG42W3F8X1pVIuv/j5n3vcUrbO1yr7YbVB2efu0fi
rf1FxvXXG4Yi6I+TAz94N81Q5GEyW7QnNe9p2xY/oXLHg0+cJMgzfTsxuwGp0xVNTfhV/9vnwwhE
HzT8UbHo/3rwpySMbx33an/Z8e9in9gYyfba3y84mFINYAUJ28E8EgsWrCbd+YjvPk3saQR1aGP/
VxEEpRcNeNGBCZx/pdi2gOrvN57PsvpiOLD650N+grpvlSubtg2JNIjCm0Z+KxLmFPTxrwcGqJjo
p3KvXRU5a2wV09lbFALRniN/o5EV4zrt7UCD9C6XOpz8kIoVnSsrsxemTQ/i2Zgla8HU5te96Cz+
A2j/tHtS6wAYCVfVcbAIHxgnHc7KpXN3FyAaCDl6uoA9RehQ/pqE6ADvpSQnrKfm95k/W9C9cNXv
od88a9i4SLccOWflowQy9bo+A/YIdFzLXSQ40dkp8skKYmjhsLPOZjmfWWLCGgIu9AdPtEacybBl
s+/O43bBWqmA5kVoBJli9y2ACTHt9qrmOvJ2fZDa5p+wZwmAZl/Pqo2vvFcO4F5ZJ56NXYhjU5IA
yod9CdUosHNQVHnMNmhI35XT3P2GnshDVRtXomjGgb5xc45ThHXjQ/RH22Yj2OMAvVzCUKtC8+9n
Eu8rIvCii9yDCpO11sNvOM5ga4pUeGW7j1PQHfKIGQbPvR8ZvpKlGViPHWnKDv2H46nQmjUneVHV
I3gY/ozrNQpImxHTbDIhgMOfRfZvxRWtfasf0+LbBGSyI8clqJWHucyC3cOPhck2lH9+QpVa4JHZ
pdWWg+9l6sLEu25fvX4PSKRrttsNlApwWeczwHiMaa9P625mgaGYEco0h4Yi8nMZ9LpAkKLr+MCh
okuBgxpxx4GPkHmko0UMkbmC6othV1iI4K5wgETK8thhfSEAukblYF62EJyYidoA7j5Qw6+lrFZ9
y3bmiWiyGyu/XDAURW4wgNEYTuHSLY69FDhJ22GL42sfhfObUk7Ln0J/ncjXO3GHfdunUCaQN2e7
QEzWFGBg4PPvrgbGEH9MCUShAd9+SS2UHOWChUtQKd88Pp5OFMBplQ+Wh7165XbeymYGC2Kuht8s
Txnu3evL4ZfSdgHFD91eX/jYxCQX8tGBl2kqPMYfmDKMcn8VPcek81hR7stLLucdEyF2TeD2+/C9
ks+C7xvN7t8abqJYFpm4Yz6arsnkOjzxTSn0ciyOA5c95AeHNVMhVZMB02gu5j4rR63zuVNyb16H
O2qIKQTciaaZss4EWrlXNUQs3BaA6yjlHqsCawJC+n2gBktfHeIC3EKPuU49M1bEPfI5fUo1akHF
qfe/LCQtsXV7mGlwiHLwCB7Lm9inlWnEbCWpSv9YITEm8O7vqZILcggK017lGgIMqaNQGNrmh1hi
gRdN4oe5/lD1TUChI/g/YoPISnovfcQeNEHg4DrKJu0XM9ACWk8RX3hC3xuN9eTvILq6QY1UaxGw
68bf1AH2kXKsbyu3qjdMfEEHe6JcFmgBvo3riEf4N0VfOioE2UATXZJWOBAxyuM7PRnoKnoziVd+
AdlbJE0kf9VTBypX7KXJzMChRN84puueCIv65ey8GnRnTFg6hWZxGdUkArxYkm+1GiqYPxhZcL6F
b818/WzBQxjajX2YoV3SMauX+Yu/+JE06AdDPldWL7TueBSawhKK0mujzwSpRX6ba6V2NyJI1AuA
oFJ+7m2oHDDu0ZIZi7zh4Wz0bob5qkCEhKN5R6RNZ+4VRT3tdk4Ym/yDbHgr9+FSKtSGwPucCZQz
y4z+r8IXu2M31ZdkfwCQy3ygVUh2FBlYNuF59XjOWsVzk16RsdNmxwCEnvLuYETRigGwTeQ1UlVw
mHscUVzba0a1S4R3av8oiurr+VqiCNlkrQj31y22WR1TPQFhcFJ0CtZzr89Nd1K6J/ZhIbwgpJuh
jXQgWUcnzVh/lLr6YgmEWc9TNSmKwbnyJM8Z8wxPZCxp60Zx+KKa4UG2qPLrm+XWw9PRii3UAhSp
xNNHsVpl1Vngy15BwedWZpmoomkSuFnWhjk/9UOYBM6MSRg1DiS0OVbmLynsc79+j2cbeLVQOZA6
03XwC1UJiWj5MjvGmX53zR95mChlrANN89u6LeNun+/tObHCPUkCG/qe49kUc+Ks2CTvHEzptUV8
j7ez2UiOamB+VMjSC6i0yCJQGkQTcdkvrsLNawwUaDE6GpmbBZOt+aAIcWNOq6i82IDa6B4d1JDk
gj9bsRhaodT+K9MREknlHRKesb/rKht2LtXYu8c8PNe66ESErI3ZHH44/n+OE5kHfEqq1Oucolyx
lbeWz2mUJzT9weUZlQDikzfQp+nJFbApBRt9Gk1NJNGyhNtCHskbcfyebIqRnUbrGTMiMosauDxo
+RprVSd55gA39MscBnuLOjheeR8FlAa+Js5NiY2oz8KPsX1cT03or90HU9RhRHQMTP1b7oZ5A72j
GlaXJtZLL2Tj6gPbb9j8TA7sxnFiVqgW9F8W5dvvmumXGKVyaW1JRGgOa/8Uhm5gFJkfflnsJXEW
ejs9A171kXQiVzGlmuxHPA9MpaNRrGGdL0vRVpPD3H6LD2x/Omi2cJCiDb1jiILgTAuaFAU2ElFm
FKCurkJmM9G7/t+KbzDHC32rZPI5XoMVr6AZahGK8qZ3O/KfNG8uMHcaoEgq1QE/AvuysH1gwmFs
0bfetf+KuKULqHLWhvr7RAHvXo+WU8GsoD0pjWcoZ3xFycxqnbwMz0U/wOO91xChOXOV3ZsezbJh
BwyBGsVzc7CMB5y4L2lxfPBB7fCVAao/GOi5oQchCjtOXOtjq8Xg3hcORX8mVIdrsRbLnChJtutZ
T9e75TN99wMbT3ZMLEQ96xiMNdJXC7Gscz5L5QYQ5KTOLZK6gXP3lnQjKdoDTNoVxreigRbxR2l3
7QD+HopsVe8ULAkOewWogcPGJc6B8HW2gAeDu0GOsqWb9HL096ccovPiFKdElARTIZ/JUbqcFvgg
4SOWsoLaPKFpr8zqpvCBo8PQ5q6aQM19Z6JCe+opVHWzqmpATBFrlqiYmcU/umPQ/IExau+lAIbU
3GlA5inpbZC8REentjTt6hkQhsDXO8IDFO6beVcCKpHjkywiWmdgWfDFPaj+soiawC3BAN4Gh+ZE
4nV1c7pLQrNDuQBCWkbAuLDRQH0AyASEywPU52NHhIR2UWliRkkZntxf5Ely6xKHNhUrlzWPcXDR
Pp8hm0/JQ58yxt/TeVEgnmHtnghxx6oQ/nlnE4MUO27jXcA56gq5uK0rHucql4cV7KldFYAyWe1L
+xo2GnNaQ097IC3b0Xt4NeLkT+JGfleOuEBFnu02+4rcRqzmOL3WD1wVHEIie+315ONbesZ18g2m
i9+eRhKBleI1bSbISuCzXHy4RQxSHNLFAJsYm49RGjvsfrw4Q4VDcOZoYuT49VwM41citSvLhFwp
BoXi2Mpmsw6e/0uMAVO3RRR0YO48mQ2PgyY6N91KNBb+RnyVEMEDbZF/XDZITlXKijsht3YbPLVU
eSL0QmpxisUTfi6bM9pksvgiWoy1X9AiLZFqGXx+7OqzD1wBzn6SLrNZNFRrae0PcodA05QhinSt
dFhLl9p5sIFFo/vsWl053UL+McXFvfyt9b3wdxxs3D40UxqZxanlGcXbiIOKP4qJJOrPTZ6ZnZtR
KYqBbsPCCr2znBHf7+Y13GMFvXhpMKuCJfsav98IiNSJWObgJbqYI8G+4NVl0x79rqQCTdadCHoH
drR18VWxAJm2tWgPLsVNcT+BRUWMQjJRau+dcA16o5VFP2qtLGjdDTunZpXPPQtqSMwQ7O5mGggA
Zljpn7or2FVAlj9fZOqKZeX6ytOzYCb12uowh0hk4GyXcFHPotxIFKFoHHYSVT8ltJGe2HRSOU9g
/K2wv3fjYkq0L/r7CLG7WpxiCxf3NwD7ILiSL7DRzPLH/6kkiesYoIkz0XuOLhB9sVdPY2gOa9h+
kZrR19USa6b1gBigr/Koed40jFS5yCGHNpjsjlJjKNLlKNwj7g2B9yPmTan4PKbZUTsGJ7BchPq9
E42TIYPwpd6+NGHNLoO6Te3BMKv3Ebpn/FRWrIcGeoiCLeoeTKJi5h5FfpIO1fZKmpqs3NhpqiM3
906wlLNBrqo8zZpJGl2BaWaiEr3H3yW5VDtiSMioYE/s7Xj9Ec+cguq4+g4JYnfFjqNKgr3SjRqc
Wbc+TaVN8zxaBdKPG7q5Zi1qliPhP6nsqJj4cf6FH3ONFVCD3RB0sU9hiS67nArBL65Wz4j5sKnp
eMrP7AGZCQQ9o/u/n/1vdeteDX0HwyinSx8g8z9WEqfeDdiDPXiOJvg8LY6F7RJFlzzdJwkhwcT5
jNithWjiRl1Fs0sPU3Tnx11A7WpwKNWgNCyL1LfmJm2lM2nLF0f+hNbe4EWKnWmLve23B549frVD
/HOtE/m4YmLg7f21LJ6vrdA/2DCAqWGLlihFUKp+F7knWaCd9w5/oCTaAvAidy4n0jvFlYcpL3nG
MQuBm7RrSHwP6iMHMHMM5CUWgfWyahrNAAyyUfPv/BsSa0TReTgGg2cdxvju/Fl8D0m5AMHBztJS
W/s8WcL4YngEnr1CWTdX+PGwEq8HPq8gKiHkjCG/OdyBLl+g1C1y6Dgt4WdJB7IYT84VIaOfR8Wf
tEXhIPwbhciFLYSr6JzldOQ9Dqsp+1jZVwLif+KLgpoBTBRgIcLI0jQWM3Xk8Oce0Vh7XLHrEXXf
8RbO8aaas7KGAuFDrxLZHtR6vZwN+TyjWhoAZyXcWlnMjihGXF0KLol4LJKp9ohzmLYkQAgsalZd
HJ1rH4wYj3X9X/djEzwHvAXY/DowWnnvNF3i4cQwr0g6CxYZ+7j9lfUbSytUzQvD/NPdwzEPszOm
uxO/g5xH1iPX745i6bi9gIDbmRilS1ROOyB266uTP/gFftj7OpoS8wMOFFGft37NetkvA9iRDSbD
SLTo5m2oIFn8Uzr/zPcSNtgw/r0GF0D9pIM/B8tV5SGC+P1wSoYEJkFavCsQM330RyaDkCX3SU90
RhDQjoCb54KXmNVYmzGnc3l0/luaZtz7L/NlAdCnAbLHJFs5J1jZbED7fNpfyIyfYBV3sZyOWjhe
NW16OSEJ80V9Ug3E+ZcQVg4zfhgpUjr3IAbkWc3I75KhmGvSExdr/ndqTVYVl/CcG68bgzv9Io7g
/T50RlW3aZ+Wurvh29H826mjFBQq/bmpyfkCiLbP32H19mLHtWfo2oAHG5aaVXZWm78wECMOvmEc
bwv3wnnPwg2RyqSiMinaXF4kOvEQd0hVN1HZbfZ4G1mK0ONeIzS/jKJzC9TOwsopjk3Qyawqtxjw
TrWcsilUnaDSnQPINae4H1EZRDvF9n3Jg6chFJsuOUnYTQdUN4xtGRKtptkdxmcbjIoga4bx7WOK
0t1aYkOqrCA6nd1NBjr0BKarsSE1hA4irMP1wChT7A31/b93gE+qRwnfxJ/7jGyHlxZlwrntVqAF
3TLvgHn/XMbHNKh3Nv7W+9L0ORNAm5D6yYvORhFzJlUNdeBywgEgHjCB7fAphUzHwNF9zyOdfE9+
3MMF6I9ThzpCm0yxybehcD+NiFz/GfedZRiCVFPxEn462h0UBL3Qcg6PPefxam4P3W8vnA9fg9s3
D9mvhGcm0Gxh0JsCe9OyRBVB3pV98VwpGyugqQc/xKGzbDFQDntPEHp/GECdbOXuvtRvKuPsBwH5
1cyQ+gJhiBORbMNqkZLSyBI30nwTerOl/aPd2D9Gb7DDda6yF27EdXLeyYjWX2qG1uL3D1mMwSD+
32dFJKqcn4Uk8mzAzNhs+XOZN4z/AmSJaN46DdQd57dzb0G/vfNBU5qNMzPPopgnGhbYKabalsbx
uF1+TevkMugGTFnaxsb1tEmE2KWPp/8pAO5nULLFqRmMS0R4W5tAaqHq7UJMUZr9R8HD+IUB82/z
74Xq6pLzKYze0owze8hN+FeRUNIL1S4RaNPVdmTwhjrrDFO6Fz2Sx0WpM/N5O5GCEpLWJ3OAU7O6
svFhklnMRzvQc61b/IlH1Hex4bhgO3b8iw0cfBQJd+9mCMcMZuzS2h+z4zSCOTJbq4fgr8bR38mT
rCjDCG2IG9Y4RpIfhwPMA6Yie41ZEr0+3cBhWqbXUakq+Qjmb6hnzHcOBk4zwRPkiGTiG2XNVjNH
1qFroi64c/S/uhH7Cug7WiFbLGWftVB61y1Us+fIIQorDAW/TTGaOn19OTX+fdLuV4VmkVdcror1
aMcNU7csQ98HR5L9MmjrTYzkM/i6CAG5LzfTBi29HVQCIvz5FSKuzH5HCkt7L1s95e0gCEzJ2jnf
5m7Xdw7mdxmuXsm95Am6X4YIlW2c1l1HNbqMQ8SsBzmBwowf7eVZiUYuAX0BDfbH69Wtw0kpqzam
7Y1V62w5tIBP3VN3lhz3pgg5AOZINBcIoKrGu3xQm7D2DFR3xFe3nfjTzHcDzM9InLg6493y9WpF
8WiXaGtkZ523UcxSgyU+nJyMcKFzh1jTgHA4sT2WQ3JdMOzJPhq1qfmBzvAwfbqdfQY3ZQazjCO7
wpTcJkZDAPwu7ZqZVfijF4u1MStxEpcS5o3Dmmw9245EddlMujvlfBv0b1KzzbYUi8kMp+0C/0Ph
qA/KHYX1POUmZKWO1uZ8HmVssqrvFfY4WCZw9cg6iGA+NqUXmiBQnZomcu838rbeaIER7B9rjgh8
U4iR5Tihoj5PKh7LRkQEDCvqxwzjVzbbfxuVYz3eYcIz2kB/wpzJ/sgLu5emaQMvlewZ6WHzaisX
9DO3ZHV3tx8lWQnEx/DvyvnTbDWqy0D9Kqd9Sdhq9jzM6njktpp4kOlV+G19pDX9du4WHWz+EJKY
wfbFBEL7KUyuwqp6/IytfvA+vCjDf1LfEKHA47/srHUflFSexL7cN6hhoUYjN4XTNSOCx0QTiAI6
GS32TkfpFtz3dG50mvj1Fd6LyH6v6fVDqz9fcrP+tfC03FkbmGK6Yr+FdYk2Jj8ALp53EOD/wB0C
yN/MeZ8BYXcSGi2qMiXl5Cz5SugZHOP/ZtA/+Eajabg6DdraRapWx5YSq/1hGUimmDLD2c2Ur1m8
Rm6eTGJADBHf6xbk6WMyhmQTmgMg/r3Ik56DQwRPhT+4UfNjvteMliDQtx6TU6JOawwTjl3mxK/D
nLDguwFLYD5ndqS1BngaXzke/dykKHQMtkXvShdbx6P+95C5avQ0Gr+rnEE57FgegMnll1biHOsm
qrOd2i03DmcR6ManuMZDf3o9p7gyaIpO4y/avk3IVH7jSQRQ9TvThob9N7VXlTZQIBwYQbla4ILw
GMNPaYgLGvl/efW9E1Sbx+jSSBM6uxhvm/huPlVxJwKNbJLeBB08/yYqHH/1nU//zVWE+Td6oOJs
qBAsdFqusFB3KP2E2F3ySITqKyCSnmSQdWrTA5+ILDUkgQctly7kISATkC+40oBOGC55qd5Pp7ka
EvOUAXvacwF75T/ID/kyQHrQDdj0N5RZFnRX96UU02bZM+xnazThjCCzUC2uLvhvBmhtESSXE55a
C2hOhIYR5ORoRwbgY6oS72gdJ/bZf/8s6Z9YNt6dtk0q70G4TepbxYeFcvvaSr0WDPuYzHCpUVTD
PngBInvMU8tZjN249+mM8nTbfF5paNRCEG02cBYl5SEQjIWf0XuDSjv5nJLgSI9r1dl6JuRWgxRN
iwyNdJ6zfVdQ7FGMCXhvc/VWm5xd3YJiExUAKhCsRFwNJmbOU57j3N1wTK0rSiebE/G5YBojgJEG
ERpfeyCk9bGP4/etc+uEx+hehyhS0c8pJjLFxZ4lxe9K/K5viEVCehX6+8VUXEmaNDregihP2pis
WSE+6S+7X8Tm3sSyIyCsD/WjOpTmPNNX0FPPct3QrsV342Opc2U+jzh5/Y7zg9IyAlP7Lj3bHghV
zhrHY0g+XtQ07MZNDcKY3fyMwAGN2UnEHQkHhWoSZEqWsLXtW/DR4OogMfqaoIE2vz+ukqAE8Ygu
89vpVS/ToPea4cVc58luc2pl2g0yC5mUPJj+MO4xlGP5lopl9tWVrEFdAD+oFhcYraEKfWqXz7Af
lDI1DgRSpyVvpxxkQRxmM5QRQw5ttBydlOi3g5kE/DOZIyRt7p3kgChNoDsO/hOamoHQJQsVmGLp
ViMXdFrwzT7QaUUOqyedv+rPMZ4tA7KBiGF/G0Tg0n375Ik0111PxrDmzboLaBTOdikpChWw+haJ
pxs8O9xptz3e8VkY8ADR6b2RAdNDOHhF4MO0He2LWwe0XAZp2/7G5TTIlBNVQKGP/YrG5PLrD7g7
KkYbsxItKmVSse1cvR1dvxfpqGThxIG+YBgmwuDzNrFA0SbaT+K3np352C/C+zSbtvfffuonQHT+
eirhG1YMr8w3kUPkTxhKl1U9M/FaJ06sukH5nb4lYkBM2dJ/zAQLOC4Gakdx/YR+3kr+R7YtaHjr
6+GvopJhaj1A72R0jaH9gTNk+moou6XsWRRhpab3zIm7Gd9oVaf4A7NDcIu8Siu2Xyq/wIuP7RDQ
O1k+R9WU0PE9ZSBKpwqDH8L7+ZpWGeQEJX1Ka+f6VwvWlmjja6LbWAFiAwcIT7jVkbR7QTdXSwac
QYF6MJWuCZduSp0yklx8uZ8wy5IYQRO8LpTjqHFKysFupRVl1PXWdY4bEtewPaBoQGswNeAYYWU4
lbKpzREPpRpHja2d4vRzZZGD1WQxqhw/rdmra4oChTukIsownwyxmZpw1JMMBqlOu0zUquWioMvB
1DC6wa3Pb43mv7dGoKH7lWS7Oc4PTDCRFBK8XqK9j+k1HT154y/AxcHcdKa4UBpdnl7Ub59W8NX7
8lCc7+lbFw9EusERI+csisr4KKpsfIz/R5JcFhQYAn75sAcLi06LLIlVYGs8QHC4umeHpyCRMdzg
/yYRKNz51AIfcGwQuTvv4tzvWQNrbs3YaF4KjFCbhGdtchRdQBLWIcveV5eJo8YbUCf4Yx24D92u
k1VwBF/lrshk4dEsgV5TQqRwAGnfIT/Y/2HpGXnNad3fbQ4Rw79ffuUbvkwV2tqZ2eT7apkJzdwb
bXdXzr1tCqb+y7kYALonrwjkRa5XGDS3k1VQaZ8c7wuawsquqjMPolOvi0vz0h71fHBoOXYxDk+s
fnVceb0u08s328g32doJDjzTl13epmnR/88v7kY2svEF9JyNBel74durNtbnkBg9cIvFU9NFoJeJ
3K7QWTNa4bC+MutQFBu4gROeOWlPqJ0nZEJFlqsczgkVpC2l8MRdjthTKCwXXcsnIVKvebR30E9v
P/DjxKd3VLXZ+cPBjRUapGQSIxy5LH1s1PYX/jF/VxiJcIHHiLE6gH78WewS/ROeAeXfLRMj9xhM
ecWOO1UDI14qdfoAn5UTR3T5QkygC+zWwCJWhFWCil7lmsBeBDnV2GdwTxKpkE7RZBFlQd1VlsR7
3c3oDZkvmsdYuB9LI9fqbJWComeWUZQXX7Qm+EWpvDctgUeD2e9e+gmmIv8GHUlEiCtujHHsEoRs
CklM5hvsT/04F4zg8ZolC4xZ7XiT4RIk8ozfwRDnwXPwzHrzZdv5xc32MeVSLaTShJXXYuzJy2VC
IjnEZVbq+/0rieKIwE4Ugs3KTflhYN4YKZZx05u39FUwV0tTULg61owoxjaKUB+QpP2yRFb56+rr
mcFpeSSQl/Pu/qrX44Hu0TTuWXLDmPSk38wFX9asEGfkRhEdhJq0C9z/1+tvlkIS+3QZlpaK61xV
o0KRLtU7v20bzelFPoum8edYAhGHC7fqVk7Wa7i3vtCIyu3hFduIRZypYEtE6gH3eabF70G2puFI
OrPUx9/LZqXwUQVbVbB+/yzIY8YSG6sfiL5lnue1ts746c5W3HamIXYcH/BIHa20nObGjgIsdEtW
pHAkt1jY/cUaV2v9PPjCsOAX71slUrWYoeZSPalBwiwJwlu9T5EmWfpYq3uU332pMIV4xDPBGkfK
QdMtWkAzEH0VAt+Q20lpe6dqCFp2NNJT9PaHw/YrXuqOJesTpqGKAQRjI15OkILVsbsKYeHg+kdJ
ldrUuf1j+OOYHTXQmnK+E8HKBIiH+ewdgZGggF7VDCk/w+p19jXsiG9qBrBWjzzwL8CBVEZ9kp5r
ANrXqP1NuaZUEx7ffBwNeqtDQ4BVbw0wWEDANJCJLpTuqo2FTh3XqZ13uBm9JEHaE0vbjHLTaS3/
Wm9AUcSSfSaRUJC30qEUmcdOUn38vsMeweK+Sz4v4RnFb2Iw8SGcqJtko1uYvL1JtZmtGRIuJ2y3
/qa8YpO6FZ3mKGKD3E2BZjgMMyuOv4D2lPSUFCvkIEgCMzd9txeX71DGM7zsbjnuKC6kQvWZVvma
TLMlES4061rlE+aUHQrNVgxquejD+ZacUq45c3iwvUx6Wq8NltyBYnJTSy44yMXvNh/F5KdPa9qE
40dDbxcZcPvucSW3NkHNRzA0CZaFQbigSw8ELvFVWUzWvjwxbno4WfzFq8LZ8whj/iSKI61DmyYB
A6qvh6/yOpT/Pnpyf4gbK6DDIpcfRJXxkZcMqJ5d82+j9Ee55Fl8SASGJFMlGpbN/pOLZdxDefpO
3i81CSO0EtjJCLhIfpMX3Df91yBYYSqTNP0+dBMTv55MPw3hFtUTiSzb6MhogY851+rdBS6G07+r
LTCcAINTq54yZefrdIlgIFPX+tDMP30jvEKZ8qNDHRCYV6L5e5zAQvbwrKxTkv5itv1FQiZC1j2i
vGtJ7Mb6qCN4Wu+7k9ZQ3ocYz4eP8nOmPgMZC8gn+6ZdqRKpoA5cZtvqIlv5DglqxpMzGgZHOVSD
muTGvxgMtZWTItnFRWAmT8SdcoPfSY3p1j0H6jJ4sy35zTCxxTuH0qJ27vwQs4AjqyAviNhjDrm2
mjIr/yvVKZ4yzGQ+Hui1JsEwb8DbqIphFhS/LCvOBpw9wJPO01ipUBNPJo4RoNMhwt0HxH9w5eGA
bh7psklFvewBgchwJhegZduaq3IKrRjO/dmEzMA+6wmRzPkeJ5o62Jef4IAkXNRwPWFc0YIJ9Nd5
qOBHkDxul/3o3FNuwTj5R0W3qht0gCgK0XJu5cWU0jQEy+bQw623zSFgV7G6suFjXBGR4JUognpL
U2xxPv/1wOc3PPmuudELjRyl0lkjfh2UMW7zqrzO1QMzz5udkopjhh14+q0rZ3qjBl/iZ0uyIxkR
vvFxIQflwWskHnaX0Fx44s2mEB8mwy4Tb1uNwBVMvmTJWAS0+xBxnPKQsEgE1iNIcLk6QQsJ0+7C
XtxNNjvb2JUVKu5TjmSc6gVaolPO02AB0NKjonXZlVJD3PIYjqX248oMuHVModbZVuIeuqq84CKv
GjrlhG440hsrGZoBxPsOaMOZjuNOEUpvS8vDqS1xpXc8sIVVcP9GssG6RA1X22UipKcU85es7ZpS
timF69EJSgzoCCZQdd6jKXFbdB02DCbZVcly+DwooH1Qp0Ws6Tno2FoTGMRCZaX4awkN5oa1fZ4Q
8E7h1zxVNUGnEyDJFOjepMYaGbojQC4Rpw1orPogp5EiVScDOILtIkUJzPuJfLE/cl/71+AFxa0F
uhhVjiYdqw655VohcE2DNK4MK53un7icZvypnlTLffRP6PQsw8c6Ja8ibR8bs24FgU4MCFce7NaC
ci9MJxgzInhW7fIyhT2R2I1MSXWl5OaOIOdBFZ1DARe5S72YlFjg34k8+KfQChJ0SzrfTqPtUvNu
tobI4Nh3Ao6uOo3FF1zpbKDC4I1+IGZtGrwabdvQDCfFIvqwykKoPv4wJHYLd6JhpfhAHX5Ma2mW
A0YhO3XhhVvStluo1YZa0O6ghYTnuOQ5yuVOzqbOxhc2RG8NzRVGUcd+7HJw3+R1LNe6JLG96PsY
SONVtWzyU/2PKklPYPx7zfb/Uz8Yfiw7m8ltG2Sk3byPJgB7LsimadHdWg8FNIizIzaJSa4AlSPQ
i400qxgoasJffXKeFixgNJiCfsC+cb+9FZgX2WKIOfywv1Vx/eeBE9SDeJgDavcwq8jw2Lw4Ou4R
CVvT6/Cw65SFx0rC4Y6qATC4aq+sV+qOYG4Q+FFHYyBW8fnLq77zc6oTJ6NL7yhG0baO1Db1t/xo
EWuSBo5B4mi3ZfTuWltvNofAx1UnD2mTHESoqVyM8SOnhF8VBZLTuJ5IZC/eRCm9cAxti+Pl8avM
oa6N97mbybabmQsDWcXKi1Bsp0HFqRUUqVFGRgFl8GSs01s8/WlSYD84LOm5ku/FHP2ZUlvQRabk
PGesJh/TpnkmiL8+BVS5nmpW9PSnz4531xMOGKvcIltisSW4NBihbRkjhPRztTgsgHBgNfCOzTHe
EaMq1rz/5vwEOFl75zWjoPmp7XoHBIJzUyVAs6Aqil0WEsbYvw0aJtk8rHhHIv5lYEyCMsm9DXo1
d9RdQtWhPnBs0tu/dp8uMs51p6oxqQZYWBjmoSc1Bu8U6+sWpeNq5t/QnqEXrkPUkjIUPo10pqVC
byRCBMMaCHl5cDZPEgpBkUS4/0oVQajHQ4Fv4Shsb4dnNBIyPHyGodjlMIH6g4Jz+d2nqOMe0Pni
dwH3tvAAZ8sdUzvW0eEZgsxhLEO/B5ZlEXsGcGs0OF/eKcKS1AKdd7PHHIQzwPh44xKI4P9es3DR
h6uZgcR0LyjgveD3aDT8uAuQBbT4ol/lJ4tThLjVZ+3CD6L2wDhK/kXJkeTCQlBb2UBDTL8284GD
5q/qXdKcnn4IITNn1scVkhZCFa0MZ7hEsDhIPLaBbEOMYB09mbpxPSMYfeD6ATBbM85oMmTby6Nn
hZ5XUwbYm6cd+51SmcCfo5kmM1DpC3hs5yd77DjBQAZxuH/393QVkrr6tbrgiOZAymmfCWohIw9e
0DG48kYdrt/upo3KP9RFmcg/5EHOk62ZERui0K1qT6Oo9tewpS3We41yUawphFDJuIlJGome6E1o
i/FbDHgSMTNMTpUblWQ/1lV6EJOFj/TAE5a/pKHaC6sqMuDAXcKxpWf6InG9nT39OoYtTiq0Oye2
z1bPr+nJDjVtM7DwVkkzBqeKqDKSyBbrbV20LCHBkP49Kqtp7ZrDFHgqhx8l9x6+UtvMT1umbPW9
be7ALIYW+h26dE1crxQ9AsdrWD0mlr2b8jDfS2m0wVG+Csq7qkitD+yOtK8XJEPvWCinJMcQRnuw
9DfDnCKC5HFFbuY0Y5w/Wy2J1hXq6iahaeDz01tfVYIHcaIBtV2hZyzkdCXbhycJeh404iSg0EJH
tFk6NCyWKKSmQBYHwrC7SAw3OdV3F8vv16MrTPcie6K4BLe8EyPi4p0njx+7mtvN5dSddSlpBjhv
yDJydY5AL3l7UC5EKHkWYrXOv6LNSjR2L9QDc/N9vofj8gJKFYwzZx4buO9pwXAh654xRSl2/dXY
0qH6b88nYH991A3X85VnNhF3138vnW9AaL++sopUxWSGkXxFLL/LO9nJRug9hOPgzoAC5ZJ8LUhX
bxxcG656qDnMGLBuPONnKwbNhzCiqUF4ldkJODN0mW8/IPnMTgzAT/gVLyy2UPgfBkc8iFDj0PKM
kAidymKex6JHt4GTkSypV9QJz46h8hsQ7Ld4XYkGv3E/L5ZPxjifXBTwyR1YN4v10KsHKs0Noerf
lZ+veS+o5bt0DxZdcscVdG4Uroy8QMbQFVEU3ZfpOiN7w2ePahzI/WG1Nzst8qF3tT8uqEBRTfZ3
8K3Jw3QdsxFC52KbauoUqeK64bOiY+hCTtlUfGgS5jZtEf0mo/K3te5z682mOuQ/glzUKEssGc26
QV92xLaN8bbCOMOJdv6J2L/MMk1hjZ3lBDgVmotA1xn4ugafvD4oIOQocGw+0chhZLLP/2eEE+Da
YYfIxqjtCBAw4of0Sqb69/pwNtoM8xdq6oX+dDngnnAXno+DcarR7Pb98fo8TKcWtRrkuHSK4Bp3
isaHT0RW9yh5ye4Wl/13KK+AufHf3NygQbcuMivjj+YNMK0NAg1sCeycNbQ3y2SiABC/+T2Kzvr2
dRyVr+F/i87nL5m9XEcDe/hN/y+lJl6XvME77RKJcKusbO6TAIdsWQMfCufYNk031da/I9zTMjiG
wKebgry9qkSmSQUvYBWpQ/zWP5pFw2Y0a/ift3pMmIAllJjbp/9/VEbTq/1BuGUOiY5r7zHK19LF
WoGWEFjQRj2KFjLDvwycVdw5VGH3lVg218RV+sZsurihmwxqBsVntVnU1KROOQ1o3JseTtJJaHBQ
/xS3taUI7xeBI1QmT7FJ3Fo1W9YQ4wf9/m2CuMQ7fmyYoOo7FzMERReZbmOYc9aXPN6IDAKUW7Vk
W82ZtI97toogs5L5H7mUnVFqu2hOiu2OCN3sESTCl0KQpa9NQzDxCTF8HzMRuGDbGoc35Zf7aLQQ
BSsNIZdnrjJe+Olkq7nAXIUD6pCPEoVSHn2wXdyhQPaUMoBMLCRnWXwoC1EEBb4TP64G2L6PwkTX
u/NpfKwAYF8TCuXjxi7AInrcQp2edx4KaezSH1Y5gZUKSPgXLpmDv3nLFiv8dFxLCCru5NEVqwsK
BSMQZUUE2C1vd4zTev75pMG6C8Js4IG5tU+ePiYFBNJpHzIfkqAuf3A+NksyVfRHENoe4o69msPB
XRJyMJxArAKUqGz0c5udxuIl3K6aS24QdpLHCJAfKFRHzCtNTNOlSC4sy5IkUWkgIIp3CNxEWkM9
fuTckeF+r11Ulv7KZ+VtBqy/iUsjEkFIzrkHgHHslfpT3b3YWotq3ThbBS+orbZRE0Hm36Lo5s0i
Ul0DuakLFtBSUmVtDjkcs95wj7TL6jCzd5X/RcTiJ3IKzBGTifloApg+Px0eTtDboiE82K9dwPAj
yp0RF/qk1gZuXmXeKILv0dUkHIIj38pEIVfXW0yHb49PcSL4HY6c9Nd2z/1+QRKutPJZ5VZjb3W8
6QULoWsg9/0FVJEIF4lMcd/9ySB04TxmHH5VVIS/1CMEH+k0uKx62R4t7M7De1COJDHsH9QL354j
Wrkkqjj/VfxwIqwaLqXL9IQHkg5v3Pzl/N+taiFQ2eMHnrWwk4hJHfR5YZ0KGne2V4z/A3+HHoyy
34Yq6t5ALXfSiWEO1vdVEcEdNgbyWwX+d/9omGXPfb0td350ft3fJKXrGOF3T1GC651wbmw+KnRr
n0vokcZ1oB2iLJxQbbFrIBj2hTZS9iQMYo2q9Kh7V2QI50A1oV8HeMZKzQ1goSL/mQeEvD5lYH/2
ZurM9MBDZiidLCimUW6uCQFp9Wj5oC/wUv9NpZ05Mh7hbZZutmvXRAU2X44zkk+JYkkonaw3YdJc
w9UO4Abpva66IX50HIyBZRfQ/D5KWEkMfYdSDgnKbitN1yyCkSG85f5hbIskwVFpTVJ7RJqZw2UC
TmyRz82pB+SDGqw+/09YPjlUQjaNjYOTnF4xQ1fW+/oyH2FVVlth3INTH67pFpQ5cDOL4oxv/SOH
qdXWnkLpb5j1W5Ao8CIOd7gPT1ZYzNBv/mkLvKmUqi5VnEwA/cQAWq0nWKIXASstlV220ZSYyXbc
vbHRlXx7Fj6gUdPjfDSh+HGcwQZXtkffkGn4MOyljbDjg5BD66Ylr61cV1cWQEzII1QBWF7Wownz
xflxubwERyWtBYHzAS8/5Q8par9UHh0x34x/7jti/ScIpiU0v8CU0UVf8yuwL+P87oy3GVx2eZo+
868fpkBbaEce4t6t5mT6tFOTQtGMuh4xYsrU9zOhpGiqaR2ktuAQE29OF2n+JIPMKFSq6oYHs83l
vuj+JXAz6pC4LY3qzME5xM9uN2HiTRoCnHvrgJL8p//1Vai02/JDqYoNjc9MRUccjUWRRRTFpwD5
NzaEx2fOB9VuM/WnAmmlRHaokCRpgqy3VNN3rogVBe5XCypoLdBnvf1Md+p8Y9Pfjw0IzNnjIC7E
edydDrlj5CXUb7mvvp2SaQz4MS1DV0rfoUgPm48J40bK79RfFfpjIjBCfJAMtbPIXWi3GoATJBQb
k9R5XptWXQhG8IJDOGplMRCa8mlI4MnxW5QBwjkfmkS/xkb/AqUZOhsOMFxVe8ZWA26Z0YwStpkt
4Xh6YlNP94E0B2wC2JoTW2nv7++Q1wfgzFmq3J3x3oG5AO9jAQwvVUjOEoiRckwh9VGjIoea5p5/
JxjUwzBG5iAzgU7n+wT5apvxknMV2TV8GX2h6Ak8Sv0xpyxlhkO4jPza64wD4slt5T9LooyKGVrF
KXiKTEvxpi2/+aXcwgvDqARJhE/nCAv4uMecpcPAjFi6aSowrhj/zn0EqC3ih+kUqzqarE2f+tTq
RKOBEXam3Tb3ArndA0MDqoc5qm2ls5IaY+3ii28uU2wwo0K1LIMjZEpWHzdfLHgdAo4GAOAbJVVg
5syRuVGMPTMDAQosPnj6tTSPerzjQHAdN0IMOykixYBjWkjht9VhiqiXhgx6UgXRJ8u6qaDK7JK1
iLnHreZsUnnkbWmL3sjm/MJzT08tTz73u9IiMYqo9PmPzgd/5iV+JzjqXWXksjyN06ybZCaTTAxG
YyRruJp+whXO1Uv629n4cDwTTH5DmE6pl+SC8jP4zVPNkjSzHI1QCimYZXhMkDBIcQCrkRRxurUK
c1tXPC6cLCUoFSu2mAnkTIr6w6vKKZjtsp1wFOxtyAGgvhPpZE4qVSb5qW1HrUa3flrHKPLGNSlc
/Xvttl4hx5VTHjFjR3mnUXxrdspyFUASo671fPAnrabWJBzJDtl/432zg7Jh+dU+1GvahpPpO+/3
FPdFA5/8MyN2I86N1znkAK7fqEX45YcTiwakzMIVihS5Rpwwgvui6i59ZIz3EPXwQM7GMt1aYb9Y
qkxRzpR1uSBQ5hnmWYSCjolI3sTbRHHkGemxzqvhBp2FXGpi/Hf1pAME073kIx9X/P3Lag+ZA3Fr
ImZR8CvbrKXV7gDFPk9J1uxeI1/XItG9qbuaUT123wjg/91hfYRMuWyTauhBUvnmB34VlrkWfEYg
QSNvE7JtjR8k+rQPxnu3/1DHULH30n3S9hQBYVV0EdXqfwYuW984vdyEop35hHQwnEYsC4ZGkPO4
HrPrk/jHatJyBg5IyhUBy8bfBmQSTHtjR60n5vHxOmiwHJkR2M9kDc7frTA1pkh4vfKnuRu75Y1r
9WLLiRphJfFxuzKaw1qQ1PiR5pAY72CUoK3FsT7SWZYZwiC6yUIKJdspq7uFMj/OueFlxO3sZ+m7
vV846GCaRFF6cmUXdqrfAESUcQfG3aL/PwRawhmF/SFLMlARJILZd4XRm2wYpiU8kjJIs8UQ/5Uc
+aSmmk1b4bHUEGP3mQ05/Qu6ZtJx+moHGPV9W4wAQOSuzoTiGbZLpQ7v0Yx0AEA26+zaF09TRiCs
GkIJwvX9xT7DD4HLRnOunGJ6hV+fkhSFFUj1uVklw1gQBVkhjuT5XvsMIoHtPrTHUH8obLB9F21Z
y4gHjXtX17yQ1UuKr8ZD3/AMMuba8ZH+ytERp7DUbiOi7GRGrpgPnFzHiS+rFRmK+t4PQ+p5Pv4n
xvjBLJgmW4pmGGMPf2zYkXcXnbEd6cavcYMxyQLoZzrjjmJF+3LAm/IX92guHz5V/OAqRgrBoUal
oecZkuXoFg0IJ3vY69QeW4hwDqP/HT6PjRjUVciZwmuAKLVrVeUTJ7tIGQilmG2IAj3zXNscMj6F
TUAL7wUy2uDKH/EkOFn0tYi6Z6+Uag2N3tDdFUIORoMqHtgjRJ5LkXRadHA4hakPv7lva8hF81TB
IofoAWmx1zG1YlPdjiVmr+T6LHKksRUdt5Wvk7K/9kg83fLH6m1qeaoalbrzrdlwndLVNMdrwodj
hQFsRUw+ePIWC5wmGVFdWugdapJd8uutWVXzUogsKEVvpIbg+/Lyy6HYHnvSuGMJ+Zwg/EChfccb
Lzier3dqiGQfPDMbawWxiKsykgz0TmaK1ZEPKcCGd3xI5Wbfg9rEMe9RYyUg6t2CNx7rxDxQCRXE
yZZ9eXEu2Q769yCoMMSCOr7zwOiUVkpcFczSyYUhqMaYVFJzizMqJlmU+JAN1WFXVoX9+xqowd7H
YP5XOX0vYkLYFxPKgPrx21omnwICh/xQDtp80c/9+whJt2l+PU1eCQ4tIL3WJXmysBoSOlKWYpJD
4kDnAO42EYKAhY12DGSVZIDiikZNXnjdkWGleBOIuFJZM9iYnihjNLGhrKCrPwQGQxdc0c9IhHCs
B5BKk+ZTRiOZPONgGPqPyMNDhrQAkdCd2BBEDmCFAHe7CizquzkITNcBxZ8AJ6ZhkN9co40E0wH2
Fq23ClcQ91yq1MnyXqD6Q15xMHjmnp5lXsLrK8v/z12bkrLH8hQ1z2p9zyuErnBQryMNm7DkoZLp
eNU+zbjiVaETf6NRmTjovVUT1r5Yg2xyBEp6gyNBscGyak8s6lJ3Vvuk2+fdZF09iuRmA7gohjuI
N0cwBWjlPY/IKXhpNDeR4qGwu0Xw/HtOE9d4oAgyPXjauGbVKPPeH/ndz7n6QXvB9te7aN5vhPv1
/l7Wm6+ABu1MiAAOYn6ZrKXgDR/dU7LqNSbYzXld+5QcDquGQFliJkrjCYVqLixbu9clNe3t+a0q
GW8sO8xChQ7U05UeQCP5UqsBjsnmEArT7V8xN1y3lfhcFByNaUGAoGaJTF9HzJIzonGFG5gv/NxH
ZBNQ/xHkRRyTknp6BD+CRUm89MfbVA4HnBFeRQTAdrWO5slZxa7ayHVqVAbkI9NlVco5Os8v3wX1
qEA6Mu8vtOeaJPovEGu0oXShtj4tz+vhKQDoOsdZ6ra9Bg5KC7NB/ZVK2Ygeiyqx1YncE3lhwjj0
iIGTANNBLfGFM2Lym8vZvFqJhT05+IOfTFIPLlDof8a60pwiX9b14HNYQFoCHMaPQfhVkdAZR3X0
O3PC3m4Dt+wOqRz2MobI+XDDiFyiFVJGK1ECv8a+fwMM9+DpG1XUe4072XEoJVbeuvO5708fid7+
0tE/8Qmf655rwDar/32w26z3GjApTv9H3oi2WFD8kVJMe0gIWPI96DCuKqRXOLqfzDoh4FnAK8f6
/nqyyXbTAOIBYZTASV0BP3OfLGAInp1FzXCWJt9Bee2hgCHspkrEmqJ5f8BHOV/05m8faC0PPETP
he+n3tciuNhw52C1+2esabcoSsYORy/amG2rT9r8FOwVMPMPRSPOjfjQY7ZOYd3VomWVRSOVaQba
cvOLa1PNSstXf+GoCaj9Z3SHblXw1oYPi7Xqol4CWkZBvHgmzQXAmnJONQRuICHa9z9nvAMK49yw
QZwgkfpf2f2G8n+QqCjqe2BTfT11ZVIjzFCElpzzTQpaVSpublLqtOBX20BTHFivde5LZp9eKB75
9qXTcSlchCbg6bX+ELH2SPOhSfAi966/F9UXKj96/EoJgBVlbyuoPt1fM/FBqrw0JAl/naqLyO0t
+XYxB5xtXz4gjyb94g864M9YC7LeKX9JovKLpGF/z8beTAKagHhef35i11ctWMl0JRT6YAg0YjWE
Wwa9MwlNqKLMbR/WRSAKVSXsMjn/5XaEjhu7J6OV3zj6mE5RPQtUwTPnYccthATV0NKTV6B+1Zc7
3JcJhO6ubu7ccnVKAWURf0xWVOB5tFtJYuMIOEBOtzWbSG+PGY6UOKWXECl1BopytriTN+sc/ZY2
S1s/kcPjkOiIWKQrWZABHz+7PHbMbszt116Ok54t5x1U1HxwCF+qjCv9m12+dcZltm0f6D107ffD
MhRTQBKZoaeevDYACtbZMNtlfpILusrJQp3LNHnpZpYwGpHLjFNWvUfO/FDmOXBjUWbj+cQwB47s
cx+yNvLp/Xj1z7Kpaz7cTRZJIY9uzAcwhOcMGYj65orX4JrB4XmWudY5mqOis1xMJAFPFEJ4uSd9
5L1G2Wt8t/2Axu9sYv1xpq1WrGFyGeYKixnZLdKTOr8mrHiWzi0XmCqmXnzgnmjyTDIY3NpwLFHr
8Tymn3tZreCK79PH+/qkOOMJhU9AqZMPQ0DUeJX9zsZ4HctLHFW03ouJigjbrTcrQKfyvqG4q24x
ytI479piqvD1SRvG8G+EACHcyi4XnNhT/aClN/5YU4WdR45DibBaBM3Vl7VW1Pa7KEUCoz/1mj4+
rjCV0VOSDIRmO4BN6InHjp+gzW8qM2mFhqqZzD7csWHwN3jsiOn8c/y0mDCtlLHFOX0gW9kg4fT4
iO3zseQGNE9RyKUj8qhn1IZnR/86IJnHU7ZqbMkvqHrG7KoyeTwqCnwxnsGkt814ntZRupVNCc7a
HJf0GHfkKV8RWcNYbLeAbnhkIIUBvrUup1dp3TNpKo/64CSysgRdLaYsF948rBse52b92cfRiG/e
53tQbJsLHud/70aHzq9iDBemhOBhzLs5R14weluaxcA7NEmK2+cUe9PQXg30vH45ZyBmuziP3vq9
4teQ/iEX0WXqkB710nv347DMgkcoGrlZch/rlxSWG7zv+5XJfL/y9NGIol8dVDeq/FwqHmwpTuDu
G1MRFwR5r9Cux6TzoJhJRmigwNbCB2G7o31CCraR2TPjsBeHMZiQofr1TfQWUZFrSFwk4VxFl+BD
qCPJzCtgIqsxLdJAXkdOCq7rjxuSU5btulXBh94Q7S7C44RyShGXR3x2fchuWEK2gaNWSC6IxnWW
GGBY1H8tzOyBwa13fSZgtZ5RLoJwamOZ0w2sjuSpn/u3LJ19/EsIR0G2uaadGp9eupiaM+jH4RtD
7NJsT+lZ+GGBPvdEQotLyq1TTPUHgVAtCf29QT6Zoznh+pEadjC3dN65sOZYV9qqxe/G42o7/1lq
y1oyLbQe/i0aBME657GX3vZCc5n10OZnN9ufnDjmt5XQJwMwhMm3BVzLTK2W9Ox987GRlYPVL/Hp
Vj/aP8eIXBZudHH7DB0ujE+Di76BuMSUNH6+s3b2m1jebTlCaJ9RlbRF7I1j0I2Rcgz47SOmZBym
wS9wnN/sJLQ26pQi2Xyig3gGvZ1g/+zxNalIcouLktiHk9onl8Rgp4KXB/fnmokOKii+x/5yrcax
skpDo4H5U24pNLokfwZXdx3we7q3wZs65N2PojU3TSP4lUZbWvUCwmUprfuBdLuqooKM+8IHpKn6
CfHNzApvYETv95X7I2GqMbDjiI3Jhglq6ahhtY8WqExPJEcfWfzK3IX8nEXoOhOt5rUzeBrF4dv3
6SJUEhdgB5aeatGRKIclLKk2/w06ZnwO6sA77j7v4Ep/l20ATi9Na3Yq6gVmL51H1Xc28DzXD3oM
GTmv8QISyxJ0X7fLeTvBgz701okwGl3CvytT9s5XaQ2tnOdT2QdxPynJ46FO2aeqxfAu0qA3Su2W
Tod4LuHL6evauW9mCLi/STItBRI4AgnMyN+uJoyEjG8kmgLKVF9guoSRm6HT98I6yHMmtLS5WTYz
fXkAQiKxfeK+4Dn6Vz5Mc9xOsGve0m4O65E5mMkkduciukuJgM/9VDs/tHSryI8WMgcpfWdcdHTa
SK3PrOmKvGfs2Lmjcj24tPsXBUlJePL6tB5Ute9WnjNOC4TikRrpCPAi/jG1rOqiz8cKHsEV0lFo
m1TD8We/4kRbxDei0IktZDFuWEeDstvNF0XPq5ilzLxWp27CjLmh7BZWsdUEcLmAWkNnjpnOpD/J
ZUBTKq27OyFag//1pk0CqZAnSCM0kP6pZ/VQ7NHCywpaDNgNeijmgOvo2xzJ/1qcS2FnOgmRrU46
baH9Ww9wMGLSCb5B3bjVfx4jlncmBL6yf8r9oEhdLqQYGLSo3ljB5KB81yvdUHFU9lI16GO/2Evp
2aY/xrRcsw8A/mjZnz7WgiSjAVGg1ELwXBmEvAEJ8izqz8SPIHmqZWvBl7oxnfeDan9LdKVSoKpl
mJ73aMm3v7P15Jq9i6zerj+2Ma3968ssVyGHET15MMco6DMyi8m+XIfyyF4cjzuTmzd9LMumr9g6
bwMEoN92EQ1cbJ/apos3YYgaoEZ/XV7Bw/CyEa6axJryGlCAUVLP8MrnD6SsRRJerDUZws2RItf0
KlC7llfeZx/vLvOkLlwplHPXqqisT1Le6XpgXWkfvKy28m2ZUHJGGOgrBxkYkYnEfuc8i2JNONKx
YBwZ74kDOxohCfXo41GYeFsRzGcCX38FgfjTHnJuAkM9BbH3rlZe0Z0y3rBbarRhCNORvm/ewUhw
TTwoJzHuaMwtyvXH3r4XLUedzwCpICxw3zEEnj1xopmGwhap8apBfDisTpPS8rZ2pWEpRnSbNYHl
HYNMd184k4Q/WNU63lXQ420EhIssnhSmFZxhX64aDQLUyGUtVqffslO+aGEoF4G6JUzCX+2kWfon
xhtG6xRhVCy7fhu56bJYW2Srb+cTgCtwaPFhgChrG4RAGUdjhq02tEg2IDnLGNFpENGFPvYejhn6
LuDwWxNHEVRLe/leBKbbQc0D9LU7p82rr6S0Ao0+DFNMcEysOZLJs9GPruTvH2katElRYNOneEVS
bvBFBy1duhBHAYmbTV3EbqD42IEktFY3iwV3ldCYoZM9h9JIqu7qGMncGBbmLJi6LZ/v8BEhqcUD
zesWkN8L1cbLcR7Rd/gY+aN05yYurhl/HBJS/nsUON/zJ/VIpw15JO5E5C9CTNK6FPqhjCmbVvvy
Ujci7rabCE4yr/dbxjVsmFFETASPzRVAY4vi1WTRsY4SsIuKTGGhpob2I8pUKi6GZW2kMS0BDU0M
krCBX6MKo57xjKKLBAc7cVbBjjf8XWiWh9Cg+HWz9j+Jy0X65nC+VMK8qRe7HaMxviA5UHELGWi8
8S2yZo/uulpCvvPKvUqzJWijAAHwQ2Lgneh4hEF1kfglfGVqVyMN7JT2qyiTRtDt389KcsccBsCm
RYICQA+XCbqfZELbl3UIvGbg6UUWvn5GlXAhJiYTSvjvkc2VUo5DhZfu7BQvF7WYXOg38UfTLwTD
O01eIJPRGRRe0HBCsqO0yJLlezMuqjJ78l/kbFQ8fBvSr1pFAucG1NxzirqTL9eQuHItDuArdDzx
9ECbpGKVhDKiX9uZCCWHXEhSkYk9LHQyU5oCYrZEtxN2a/3r4vMd7jVEhboLCvh6JJvxK4+qxvGJ
x+/k911z1jgEr1U5JpMvTePgOPS+yYtLhYvi6CzOQiMZvMbU4+ZSTok7RG1G/6IYwi3ZzmhSZgmi
xQ/J0ZPx1tVYHfcUQLvckoKgIMxMkPGRbX23W0B9+BLtXijN9ebpUn3HWDl9pMyBUNfKKt7i10UK
FBXUvdrC5faLmVZVYiQtaM/zrFD/eEBr8OCE4epZHzcPMFuryTiHjnvVZuVeBkxo7wP7qiVMwyws
OQf7zTbfr4x98YRoPlpLU5rerRI4IxpzRIlrBbl+KOzwl2dk2T8J/aLodLwqCLCHLbKY9Q6Vj6mt
5YYOn5VhlV7b7heZGIVyJMZm7QZlyPv422vEdZc7pOxs6sg4S2gGPMz3FU/yUzgdbdiAxTnS/ecK
G1U++ptHz1+dAn32steH5mXjHqutUhtLgQ86LmaZ8zDyZLFXcjA13yNoFQNmwCkJixwEi7bB/dW+
TE5/1cEloJ5gW2tjFAEPqo8nyZlw4LHd+y8BcD/KE6W0klubTF22NhhmSaMbcZN19lETAVGpJC/E
cpEn5lqf87cYRSXiJ5UkSjXfpAMzvb1nYV78xQ65DK7/Vg8KJDG16RcsaV9nuNlyn5OLfB5bRDfn
W14oAe5+ltZXRfEgsjHoxAYLSb7IB8RLB7hIzMTVK1iArDLFO9flLO8NIX97KbjZJKJsYLkQ25+1
mQR/wQQvZTHVIlRbbeEE3D6gtRbTeViNU3NQvUtTFxFmydVqv7cexrDy2Xp0aSgdvdf2R1Xofmmm
pviJRb3aBRbUinKRPLsz8ZqyN/eFOVx0b9iD5Yk7MUBxcKOgFeQsU8f6rgqaIe76FE5g9kgcpxqH
yaTTZGfYSJrY0bGI+g1NHoJKyzQKDOEW2JkqZSQTmKfpovn7a3bAT9NF6sj9HXbGoGZlIxkVHZcX
XaxoMMRhCprdK0Ct/rFFfJYYNTUQiJMfFytZ8LMdSJ74PjyjpZGA+XQEZdgoyBA7sDywquucrC20
Kn+ONfmQ6AmrOQFycbzl1QQVP5i01PZ7M2addymuYAphdQ9xiIha/Shk9Wy5hc9V8XZAZ7oPYIVj
CqKeli9zlVdNA8NOBCUs1yjd/3R5W93NhYsCld8mi7ZaGcBkKW9iHhbYipZ+A97LgFUbPY2IACRf
BEMZQilh0E2gK7z9j/3RRatS4LIioId35nV9WyE4Ntio7Kb7Q1s9tEZmtmm1aTrTHwEoWsps/fa8
swRPxi7LIa7u9XjB+H+lAiDAZykpsjW3HYohikiY2k/CEoB5kidiBTVfDMDAA9BVRl+ZRklF6Zlc
LT0v1IWFxcoVQnfB6WPEzp7pvN8yLBhjGfIVSR7wCpuiQeJ/ixQh4TpkTHF63i0wwn32GU5jwIb6
EmA1XZCPmLIl4oW746umdoJRJxY2Yjg46nIEByBMSuhKuV6VBlNnU7EZlO48BNGfyeKXlgMSWBXB
Y/wXQ9LTquBAzBX5sbfKwG9+onIyJaBVmON1g31Gc8iBepzaNvvM0rsNXvxT3vR1iw+Uf4x6EvRI
RHGo1pqDidoMTjObucgl5Cma0dfRzwV6yX8pwAYeXw2sSmX2rFsYn1B3Gbux/JqAF9o6aC/sgbOZ
e2aoahoIIBpHW1njDO8jgwROoZNwH4715dnft7+b+y0eHTbgFAm/pcaxR1sc5u2gA5innPxfK5T9
rUwXtrMqG4TfMcBkJUF5KLL0HX52VvmknMyymS3cB4DCRcbl1BObIo5Q9wf9/RwYPt89/CmFnTT3
mk6TO5Q1/EW8pEC3llhNl+xaR9cVZYp5TXeahpGwGO+Eu3NKkBGVGdcllnBRHgXxhvrZCPmFMQ9X
hRLzNwPHpqN6XdEAJIINcD5bXPFRsKLoXNWbb10fVmLxuIyqFarlL316GnXXcwqiutRmTZBv6Hxg
EgJ0FllCLtSCVHYxgjFpqP93TGWrsMcj839Tlpy1YCfF3STFM+VktYBQea8UJCQKRAtvHWSZ+nYR
Q/tXxqldJk8wrNXWJrn4hwsS/OhZz1vtYkwAB+X9JJGFwMzbveoTjneOK7evZy2D5Pxtg6PthFcA
d0On2Yd31msqGokUS6sB+1rXwYaguIkYNIXKJrtM4WtEjucgkDKyN6o5fKgPqN7wLyUEyOgq6UjT
56It33twrUshA2JM14GhyuQJhXYGAcHuv4xIG8AWtbkmvt7+enZ3LHfXbXg5LYHLlaK60MOlxQm6
2yzGL1DTML/Z613e/8T+0hkIBE4VjoUP4c60qs+AE6zEa+jpzyJFdpH1icvfWI+3RNlA8YNpzVdy
haOG6yRpByrAsM+9cOMEWO/S2oOm55lwcoQJbW0pWoc6oEoOOCC9A9u/d3OT/2ICPdxrsso2C9sj
7IRtC470yKzZwLHzemzGpE0H96yQpUR2IAInjZlbUw9NhwIJV2UI2+g3tDQT0KAnFv9M8u6rAyGx
unCf4Ox5fNIBg1Z2w99+1QJ/K/r7V2+1J5B5dx6hn8eoLj7Yf58hi53hP0MMGkCw++qKDNxdlMDY
f6IHeGejrPtKlYLsW4+rld4xWcEqkWq5jIzb4J5ZcYEcOfZJY1WUQrA0Z7a8sytlBKE9btqeL7mM
hdZFeRcHCdKWTbjPAm/9Ehh4CYrpotG8LZDa26a5RnT3lxFpwdxdSibs6lUO7XB6ETqjrxZxfCQ1
lhs1tKG6IHdbeOP2bmxeGmlxQusGMw6PmbQ8DhNK8qs97avTLhwKlJG6GXc7yEtIsQCG7PpAth00
beZrW8wgKQ2SMGYktFyy+18z4mtBCRO/nuVG47yFCy0uFTXp5q3in4EFnjoHI9k8ilpw+8Npdq2B
Td4HsE2eMFbbK4iZvhQbWwSqTtufQWzPFhhqhxPN3bIbPmZk4jBA1R6ZFvS0EGUuI7NfRcAwNiSV
U42JPZRSvnyCF3CB/iyg7UkBp82/+JoPMZddDaffpri/KnmDUTsbFgOpFpBe2Q1apO9eJnu2vQPj
Kab4EafqLFNN5Ro4Pn9hNOnlVjLbHhh7vRT5+y6JrOOnprBQAPsgR9U9L5cb07OgNcD18m7ngnFc
XOw7yXy3dNaTWyIAseYfbCa/gWcql5ZlJymJOo2OlkBTHBsjNj06aeDCWJENmS8wRrYNQ3cccr6B
zbOjguvkhwnfwJrR8Pg1c66kB3WtHe96WTj/pfanforBQn/RTDoIeunJmzT93iIg45OKJfnikVJN
/hs2lCU6qIImxrSK+5FA9/9jkNjmmrtQ21cHrNyDF57fp0h1n/78t2zS620fwPDEKZwabju93QPH
W+hW1/Zlpc6BiWE31Sr4DtnGboOjHtWZCTbBk1wKjme9NHrBotnF4wnOTvIgR48+IZ4kKT7o6eNz
5LZuJTGIEgJ0PLNkVzrFGuH61D3hcV5fkfHHqxNjFE2muA25YEsr98d5ob9ImWG53yQOsyJRTrBs
mDldQGfrJP/T5qQorPyE8sBRkHQKybLK2WD/DjrXk6FCVnFXpgAppnKgjMnXKL1w+48HFOVGv3y0
fM3/bgMfbuVD0NHG+/c85vnZeHFVM2fJ8X0OFsh6/ocAdCwOZnCxrxX7Vtmzle98VR7U82NlzDaF
hNhL6KHQeQO3n94zBbzKxbELOeVoNwGZUh9K+pdgKQCNeu/weAU34uYcXHpI6sluGR8eNbPE18PO
ifJvpsbvIGrhq5YtGMtpgSp+6mTVB+jstvkFG/hcHhPEfwyWvtmFbN6vCVdVT6PRG2GkByFMO9Li
J+8bX/lhEs6PT+gnwLfWNvigqXVKF660vbQdgRZD/KKx3is9pkkl5fa3EiXO1u7j8TySjJTE+RWs
av3y4JbNY70mfZWIqRu7rhr3CJenfxe9Xq+WCGjCHwqD1ae/3bP/m+QWI5N8nayqhUbb7FwHoL8A
CGrgOaIsGwPAu9dqSEQCFIRY35UUgrjUgC1ydtoAX4KXQxK4HfOtQLJTu36KSxpbYtn+IeLVSbqE
Iaick6Am2HsvleGzWCUC0nKqQTMSecV7xfsYdqkqsiAFE2o6mJRpOd3aYEsYbtihNENM2Kh7RGv8
CtdM7Odwnt2PzJO8E0apXY22hTyEmIKJfw619Znh3YA+JxDdrGa2/lY08Y3CyLxsgCsISOqc5J2z
/VDe0buaP3M5/9eflOdFoGX69CdIjRRQwuZgaHGPpQI3RXvVtJdsy5RtPX352vMTlYkVqfIGKNdi
TmzbzyM9SrJvM0xYnbeIxvLTSmscS1aRbx6/6MEqEli2MCi2hebJAT8GyzPgr3qY5UwlQW6x1UpO
3mE8qO+BwEXCOXHAe8y0xlEE+TGI3TDcbkrJNbHDUf5Pr5wVzHKHy/r0hVtK2Dhz3oBW3Ko8mhwC
AbyjpjGzqxP52U75GLkK+0sOa15Mu8A1gIf1/HCafjao1DlgO0yEr9ECD25lkFzecZPePMmeXAkr
loX10yTHdcVX44DLbGm0fEC8sp4QlOkYW/Hc99fVqkLZzw7+jLrt9AzWrhiNpIdaYItq0UY5xfSC
rCzorGhTGKTYoj0nZyFIrEaqiFpOPlbepcxQtGfyTtILe4XNstwpJu5Z+yYq0S0cxhqWKkoY3CsK
PvFvAYhPKmjMlqBBEQcvjqDcixHTHrmRZfVLekdsQ3ErIsI3v/+jJv+lQBIEll8+dZOla6u813X3
eNksQFtz3kpHWCmyMV8pj0nOPnlVI/4Tv5zLkeeVBmmjF/0rj0vRR6gO2PKUY+UBKcfYrwtR5RjD
euOHf7FayOV93q25pH7lB4Bpqt3D18gbXD2aVN/Dm/fzZ2j/oWSqb9CH2d/HLMKRz9hTZhp3ochM
1lpQHWhLcufzJtivEuNyv1td8pVZXXUvU37nqv2dbWnYV+GEKT/U3UFVejzUpB+FwRVrsvPsN4Vr
yx3D2nXBkffQ3oVtxV+UkdmJz8ohhdeLXvjMA0JgE9kkTgAXhFsZZwg67E6VvUCzxaxb/hQ3CIMT
69i5JbUrqn0AW8+NsJe1KpfrH9pqLIbQ17PpDogoAA/gzPqNAfOHjTyPib59oVEbVcgdfHC6Dsu7
vduvBMENqgIqZyIweffUDwAjMtpjxU6gJoXCwDkth0/kkw7FYqSR/v0WVWpGxTwXS+YBCMXndWxx
lMP6hm526cyKfpV4AruFRh0qt+ROhlOR5KJet1Sar3bG3VVQ53yxVG7mBtTE16kxIB+bZtERsLAG
3QGfwZOBriS9/30+tCMJEyuZwX4e6N1TSRqPBmzFSFJspM5foh2MXneVVCr3QGoRe8VQhpFsBz7n
SMr/Mg3Db+BN0W1TuoHGRgNjjGa1a5PfujoKkVxVcVdNnPn2t84W/IsouuMQ2MfrW1y3sxFiDSb7
ciVaOUzPLOkpZH9Bdyn339v2zMg6v831kMB3wilV7uUD533R1CMtd72kA2fm2At3nfb6q+S+dyJN
05l+BLLPPwt3JseFZJMOxImc9VkphwIQDKnCZ9BwYfcW8TSLgD3ClJTi/7CzfdiKEegjiC+YNZG9
Bwyzjc+WIMxb6+bB4dIlVI/4CDzeGFMiGEQ3m++Pskplx9ggCvzqqpmqVYGdKsD/RNoO4D/5faMK
50B5tOainl8/N9viZVpm3oxfd1F8oWO5SrxErKsqkf6WmhHDI9mNs1n4xOKnvL8VlaXHeHjVGTCl
LUQM/5Rx31kEXw3x9ypCmX3jfTn8l2HLpRppforFH5MAodSms4gRVMIWECTlzd3WONEfL3l18ZFM
486VVORwrBFynw22Q89Upt1K/FKbFUJID0C6HeiBkleAKtBW2hUDuB2M/YlP0ih8SUknQKca+C+h
IqKYu+iMnlzZrhhDpCbVawCHzbHmB0R6XMSWlGuOnRQGRTZesb+SvwBL1u8gD5lfVhN0poLigpcE
n+dJ0M0vqvGXEVWuRtnuIYGNzYvlsXQ1Pk45qXZAbIgsDhwhYo1SsxtrS88u0TfC8ux8cSuX+tpV
1gv3XtL5OsAZeTF/ha35XNng5g34vp7Mv7UDbNnCFTLzWZ14W7BgNX3ZJiRTNLGg7ez8Xt87Vyuc
ntl5KGbkDfOPlLFETu1sJysUB1VluCMMmA2DTa/M3yjzNxmM4axfMYwsjxT/qYB+4YaYoGmVA3oi
KVZVUjfK4d2Jj6uhD1IrLra+2lQ2jx3Hk7VRu0zYNK7ioa5gc8BNRtJgQk+S9iYpiT/hvHSOfDd7
LfF5bmYC8cqi92EuocdR6GQtIk0Mm9bdYm8RPTUCYRjJFphE+J1UwaZh1LvPYGWxxeI/gLpBVt20
ABM+KDNrmqCCj4h7od1aPKq38JZBGF8EE0lbBeryRyUZ8T+HTAPzvjN1IytHs2wzzkPNQpV5ttYg
YmfvjdLoULBy5mwLeJRj3PeJSJ1mjO77FOH2nQVrC5Z/QR2fqmlABX57pDisQIX2A6BrEwBfwTGn
yyc7R1HoPuPMhn8MBTSBuitF41WrOaHjZ5t5VekYi/XL83tiCx9lZpJ+5BYWmy6cQLfiLgqUA+IV
HPjnL7Cp5dC788lOB/3WYNcL4SVw7PEMtDyHDbU6Mw21KcxoOjc63WWDLcXGhneJ69kXdbLmABru
xM3Yw5zmOL13bu8J7XbgAzs2NJ87bONoAJ5VH+Qz/vfzyNeA/zz1ZRlh127doDPiIpIk/91um8x5
1ZYC2EfdC0HW7HG9fqVtPJu3fVp8SEtWu/+FVNRR5iFw2Fpti2KTx5CnVaf0XhnmrwjUQvww9unE
O7jJCIxHCBtyG1e+aKfXsRy8hZlFfiAkcuT85QeG0GjF0vlhdQqp5iRoKJ+PQW6IXMCzo6mgkS91
WZKjIOFCprK+jRjbp0VPcCX2tiiC1y20oUiyecPOI8GrTOqpxdZrB0cPvS4MYcLJH+QFGCxkEjDc
PcIUMIoLKYqizxhyCNy9P/DoOL9L6Taz1tkchgso8am1NUVtrn4FU9NSdpTPoTK150rrU+aKKe9+
Avc6bIu0M1CZiUDhfD3K+eX2XGUBk6tKMwsbspDxd0tfNOFOB/+smMGzUMfAGcnb0H3X1YjReaoC
r5DP9uFw8cFzUXnztKddqy5AEUdPwMim+Qe/an4U+ZVl4LOqP4koAuBHhivxHBBloKHDkjX5z54H
WefLN4RGYwt28LSH/qvw1j/LAiHNl7WjZGRMbw45DVelf/c/FUm41o01okR5tfRdFbmr01AkhXA8
zEKN4QRRcyhfUP1eJXQzQpWp4kR3fAWg/23gDJl5pog1EODfD8XrGgx51OIIkkjYB6Y0M+Ct+utw
MWWPpMSiaFELIPQ2FyhtAdm56zWmFNz3YgQHf1/QUa00yR6qxPf9yt0OKWJ5mOWy9rXnD2IilnQF
GnH5fLCtIPozZ5K4sX2vcwGE3y4yU0uBhFHpX1o663xaf7qkhXPLiFSNryiFDXde937MeCYinP8I
rkav7zVU2vbEO8lgFBa0WRhE4k4HTVtIIQVDrpcZhD+C87FyGn2bj3bjX+/4KOAQQWsheR683SAq
9hN0oG/mDKaf43p8ykffcyIVVc8I16Z2J3ss/27rofgeKp8vq7t9Wp0xpzvpVdU+vuJ/lo8l/fSV
nMTmA/xnNloyCCYtNvpoPyP5cB9Ogp7kJXHHKh0+tAkuyRwqnhKx+Chf0kkJiXcIhZR5G3NLvHLe
uLNkzWht+1lenpJwtqVNLRYj9gjAS6jHOMSEnRm8NfE8aHqpn+iy4khBzg6XfMJ4J2JQtq4GJaE0
lCCQEplVNXs0JpuT21aVsLSylRQ5R4hqG5Zaabybxy1KEmQeub+0uiK46ZNj2Hc2hB5kYEU/TsSr
/j18462rWK5PxYr2OwKLLIwi931U8VKPv3cgAtV3bvUcLslGfDrsoUVfZrOgOevo//DCMCaQ0sXS
Xs17C82GdRGQ6fJ2iNC6jcCv19LR0KTQacCp+YbMX427RPITzdWEM5wRgsy9uZ3DGJ3N9Y71gUTV
OzwB70P3nqiw7JiEdjIdFfNXzldaaymNqAD8Xpw1vjFvGpikNOp9ydU1nRjsffJa1jG2+p6QuPa7
tjHbCgzdJbOEp2yeQ0maMDe8B/4hLT7BFK/fzeq4+HDO6k5XVrdEv3pRpeteEFtJK0+PKHga3VXa
enVYAaVZjkuYr2MVwFXputTiQH2/Yy0jvHLJqoSAaC3HuFmzvfuff77AKRYye2FRmQeraCgOGBni
rU7/+qO8kA0t9Xsdb+zpRPJB022KOw4kSGYN6RMUOMXgwjPRmTxlOzQrju7cqVdH8Vf6efv755iT
makfXZh645zIpGllmReqOxUonbkn5TbzyEwunE+IRytrLunFN2DUHKUZvIxDexe0+QDvONHLX5Pf
AFTtjpZQU0Vy3UKFZdPQbqCB4y6EqvmPW4FGEHLW9rTkuCh6xoRMVxyl4do/CtgUKCtUn2ELE8gI
Ao26WuwD4E+uNAtourliqH97cuma2AeBgPIJiBY2iFvCwRo95ehcsHEg+AXl45mlaMGqsGTNDjks
FBrCqQzqHsOF4tgS14MdPXC4Q3/wpTFNYFFFrgnUm6FY3QJlFD/rvoRw47O2SnL5J++k/T4eZ269
Y5dUQ5MjXojxLNuWLYoYefE4Fvk0QrsU5k1pP+7vasB4bkr+nplYcMY1YZDmjO3UI8f5dc4Y8lra
m3NgnRb1D36btgkJIlQ6U5bHXaurnqgEqU/ZVOyS+xnthqbWyFXNxLh76zIY5AbZOi3wclNyz9LO
6IfRFbz6b2cp+ilUb/AzKYJ2j/qCy1txAwrO6xlndo03ZKNFzm2w1NiUODywJdyq8wsTqFcJj0mS
JK1FP/Bhum5ga2rjChCt2xk4h07cl1vlXFdqLSWVhuXPvt8ec3LXhhLfPTPcly9Tha0iQsGoPhai
5pQoMv8lEh4Tc+hlxxBeJwGnwJJbpHbb0bvUEnkyKYXsZICWmbBkZTWIUQjWoE7GYa7oLUCAVNf3
lqp1erRpoMnd2NqZNnIrfG0SQOJ1QXQOL8zNg4fQE4ePnrSLavlFqLfgNsS5zqp/Lz2yhCX4uOz5
YQdowMkiwXz1v1JCtCNJGDTYU6nK1+qCFOkaQUwA3He2jx2iUXCqorhVTKSRq6mo/Ac5WASADeRJ
2sKVgBx1V+kdrrPjq8betGuerR1ezBFfRMgJwJMfU+qSM+2PtoVD+UK8lUmrnCBY+OEu35UMFmxF
Rqpq7hFu+VGOKlfHqRFq15YEXE43ik1ydmWNa2L9kGgAowNES29wiXaG0MzS3uKpt2N+SVSwTNkU
HoDde793yphfnX9JvU3W8Wk46tmdKjBCzwBR65f81ufRaGo+MlPZFsSC0GqYjT5mKh6/iu48atkt
N1prdJk9TNy686Obnerk0qdycMRwKClE0AP+lbGb4l4f4B+vGqwA/dTA49mtuQsoVWC3Sw0d/e94
nPYrpKfZy3nGijDY08DyPojcLLd+52CTOUuyQxYaxIN4/IZ18DlYm9N97GX2AL7kg++5Fgqg8l+8
HpDAYMVPHB/wtU9qCay6aOeK4WyS7ngyGX5JoN3re9tEmoG7C6g5OhI7NA+3uqeL6htKBXN20VPK
pnjPyWzkzE5Y/DBrC67iewd/zLIwZFt0VEeU8AWbteRkaYKnMwj9urwNcJOyZBetIB/i/Ktt+2aI
nrzA9dgWDwWnxlP2g5Lwerw+zCtPTulBurtHTFwEiLcDOyzKcXmOFuVm60iZiyQ6/ThFuQ7h6JWE
/Jah30TyhXxHNCZ1iCucd5sgTM9AgA9EvrhXjPUh/wcDsrwwhq0NwTgzIo8wXFzD0aQLFvSY7NAu
a/VCPGFlKo62tZuT0imPGShsncbfQWjHZhsD2QZvSMhRZLcmY7i56qsnHyqcFHZVROm2b2J8v3N/
Ph2FbS2WttsWvWOPvjhMGfs/Crs2PiiHmK7rgVheBzPduUtwXUHKkaxZDiMFpdMSaFH02VG9bmXC
va0O76UvZwcajrZy5G4QfhgyRy73P4UdgxbJNCDZ3XIPcsKJV0ukw+O4IeT5O15sof+ANkKo6ruh
fon5JknpuB9wtXFHqa2l38vkdjsy161DId2qGw81oH5bUAh4l8LixRa5CQs0aoSsu0UOob3HN4rV
Xf+3WdUCFoSRXhgJNOMaKnlJRJCzrUfdW8XsxPXP3XJEUAK7/eGVmARCSysGaQZYBQGMxHggBxIM
KAyjl6GO+wUqJYlOZgMobgpFjCQRGKfVb8L9puKM+fgKVS1mE6jHNMDayK2dkIUKUf/QjWy0zETz
VjSkfGmHoh7aBzONE1nxdUbo73P+bPKqW4X33ghQ4PEY++BRimELtpHzWC4OV9SM5iAXZ9wEQd1N
aYeMGW+oMnnP4Mj4WHXhyrIKugdKLlZRRjSh7y37deuDc8WhKCaZ4xYOfveFLeyBKitQh0Ca6xda
Um4SMDkLiCNOa/xbBkokSRdp9ZmtBmUpAmwsXWL26wZ1YuP4T17JqsJ0JwJN7JVC/Cq5cgpc0Bjx
z8Bl9IvPEmk0ncrYGZAVZ+CM/Nptq3qhxWeeO6iVC4n49pPt/odF6I7pUiQiJO6YLUTjVCL/3cT6
BJ+zUY4K9gTbEFsLtc+tiQQwKT+iP2BEMJN5UFzbOOoG859Gwc2Ev1yjyJ9DVGYuQ8Lko7fuHYzv
nUDVedSR5FNItCzSHH3Yojr6fPjLf/L7reX2G1gT6W4CE/K+vbU3GHsrEoaS6vfxDPMsoh5zysx4
ApCgxcqUeBsAYbFSD++gaJdfxajv7wMxrPfYbj0qKjkZ3YHOeZcs6RIH6x2cx1qRvRLn7sljXDvJ
vGz7KKKOkJ1knofUnFPglD7+mtk9voYDnddyrhyKBdbImJ9cAmrI9mib/6F7Id+fkqeDm3wYPN9a
RRbWUTqenDIgCcTCWbfjzEhqmUUlCorcgiSG3lzBGvR18CmDWKn0NtfYZIEPcy8qKmYSvxMqZe/C
Cgu6aCu51PUOltQs12JeSyp5+pEtyyV5OZCH92kRVVgH4PZkwCRsvfSo52Ff4FzFygwFBX/FkPW1
ba6d4N+TlnrE3/bZOg1r26N37L2C/N4F1G0N+dPykG1ydK051boyycWUMuf572xAC6nKeG9Do00V
5duZ5vjIfoRphzICSRaIUztV5c/7wwf5zTD+qzFVRv1pD5TrakLUMJchHWjlszOkVPhOGpIkRc+F
OeOqxGow9xyhM0LWiqsfqYmMtNEJ8OtR0yNkxG+b32iI/2Xl+y8DjLzmFAuQrc3UlfjTxgCGMWdo
QELonjAjd2aElc0SGZrSgc6HW/XJBOKDUC9mlG+gnK8lGG0dRpO93WT1IC6akRZlwS3IXwoieO0M
tyWeMIy7nXXXWiII8dXHBf+zwDeHmN/1mpK0zB3TQsHfKQlXCEY5pnaqDX3CAEPtLC+zVQvyVFp5
gGdbfvzXTngOrRE8Fayg8BVkj9rVEhCafq7mgmg2NJMtirlqHpXKnhJsfpCjzBHVcaCl1pGsPb7j
nAja5QTrlB2alqTcbOc7dfkVtGpm3+jJ2pZSjIW304LgRZKgqH6rbQQnB9GJ34HjAIcIq/wOd91I
10MPfQzJMC9RzrM9OUgl2uu2THMViwe8wxuziC+AGyybojlrHcPLzecK2gsxiwayqpwN+d950Dej
nM5OlxZwDU3kxA5DFRFLeZfgPOQ1GDMqsQKwmjVxs3mvta4egJ6jtYEzGojA+/nROls/PhNjmD4E
ZAcd5fRwQmxRjKkVOCc8GbGwcNXZUtcHwScjmhiOpJcJ25qPe+jDPElBs7Bgt0GgYW3CD7QPMghh
ogcD272CdfiF2P3Nh6uojLLEtP/4B6hVCcVrvszh6PL17sgAjGttKEo4e5qbdyGIaX6AY7HR3gGt
MTC66SzhNQXDsEPZmlQ/Hc4WZjOqPbjh+lxgDy7KLzJcmeFZ62yVAVL9iFJd7nWTY/dBSYF/itX+
NHDvcpg4MW8PUBI7+3jHEieZpkefsExTeSqRQihSsJq8aQDX0VFvhtMR9yh4nmD5i5yKkIOPPoG/
7yGGtZl9MM6V12UEhy12Eyvsyfo/d0duB7wbxguBH47tM0t2DNgF0+9TlHLjRDd3adYrmi7Sd9Dg
GvHcqe7WVKixNLxz9yBvLrtbT2Jks0eknJxHtVHBahHMXEXUWepV+3f+zSQPnRHLOwkjY2v8zhVG
ioGvaBa5BSPKPHHLHr8TC0wmCnIIrfM7E/8v4NyFSzhvDhr4isf+BB6x927L5g9F3elk/hTml6Cn
uQpYsLfZBUzAKNSOAuW9WMqucnEVXove6PUf4APg8Q6yLp5FoyyVwiQHtjCQp+m8ccUsCiRhR16s
buo/0etIvdWbDXspgCBUKy2K7rJA6ZUKNKaAIKZnr3hLcgw3UZml+TAWFTrUmP2B9tNfGPerXL1D
76+lCoAp8LzfMnjX+B5HgparKBc3cn/oeh1eZ6FSiSDauRLLKWRduhHMQ7PS0VMJ6OpX7dO2bg+W
i+HRWrGKsHil3jaJQ/4r5ao+74vvolGa9C9sH5yPJumDXWRhjjDJNM6J/z783RvsYqPGKLoKZ/jp
0N3MwXzHFuSDQcj40DWMh4ERPED4Vvv+fWL5YDWPFyHBvPsLuC/pm8bEgOugiH6Hrii0Uxo3vsjU
tSNvxUifLjmhjvVsSWeSrka83i+H7frmUes8Apv9JiuYqeEN3K8XaWgCFlrZUTa2TYO00+0cTRkL
6ghdL3VLHFQLl38CCyqRhncjA4wCfwAc/y6ZdblBLHnJdTUyjmi0G1yk8uFVPM9od58Qm1P35gGc
7ngnf+FCAOQ9QeHQa+3wh8CBF3QRaaq6EWDNUuA1gF5HDAyFqZiYuP9gepdxoqXQ/tgW1S5ngQUm
HYlr6r4rg/+VFCZYTq74A5BZi8gvjNNSC5gBF6D/1QKxYtqL2F/LDCl87kVKZ5ikbPjkq7Xa4vmm
YZ1vRle1c0ejBV7y/+y/8faU1vI9gwfmmaK7aAuzzlu0cctqekmRytP7fnLjamz55q5jm/zsOGp/
u7xruk71x5jvyvdKEqkPRBUVBZvI/WH+NDlp3nSrd6vbdxKNlQWIwNGz5wsXL6r5GG2SfanuXjeC
qUqWprIANTkUhmt+ekMH7WjNDh9XlyLemiSxhpGIW2YWO2wOzPUS4SyvPeb2wkEHMNWzD3unzps9
VEjOxH88IQcMZTtlmrKgIdqlueZSW1/wJwMh2X3BSL+sQGk/b2BUzXYddxqhYeaH34X/hPK4Q6Sd
u6R6NAWudz9qlDlhOY/tfVhl7QoX0PCn+MKfnt1zpBZhnLuCMBxNha+vGA2p7cUcb+B14ap0oeOC
H66R+CJRSqgJYnP/R9w0NA8esI7MSWxkEIUEdnMxgpl0i66rVrfA1Es9jPiyFWUTjyBPtPgfdB9Q
/gbcs+UlR/WjOSvggxRw196gEAQlZzEu/1aP85Ap8fMkrJOS3tzfaEdIcKvg6/tG0qmyWhjkoF+j
uJa9TX+zKUYIF32Qt23oGzOcK+Yl+QGCW+12Z7SrP4ZSRLevzRDToH45T0a53It3/MH9KAC0GPVf
pO/S67TkGBF6mLPCxoNz38dfU8SHh6GWSh7nOz2FvViF1FQ7maGIrvt3H+uCvAko9w0kgwFkTWI7
s9d5hj+hrQhCz3K4CtNglObjOrUSUYG8QczbTNgPw6TxYejg82Jo0n7IFzLc6KtFSPdsJudf3U3p
Rr4TMMJX8gKI2VRWPbKyyI2z3Dsw8A5LNGszpqNIunxig2QGkySKOtyOu5rsochWm6vPahlyxRdX
YzrZacY/om5AdTPCWH8K5kK8E6infW1jbBT5bxlbxiAwEOXoiZvl/ufySD63cwj5q8CdX8qncQwo
ihB9uf/GXWDBhtppUo3fbAy0FGQ6bJ2oWONtz2/KYUz+otqjouqNjQynFqYfYtEa+vosLnoW+3ig
BP9QzbvaYJ5S9AmOUa4SYom+3yf5NL95Acd1aJAMkrejUJQxcWg2vuDeHC3zL5TlSyLg3QKs8H0h
tGT6cgkEfqBxoqp9y7KSjZnLFOmDn/9NJ19Zt0J7i6+WOpXpm0gU1ZdHzkZnxQATpEn1F6Jg1XvQ
H7Q8ICFs2wWcfloLt976r+7aXFe5W9ZjlggZpFw9s71EZwFD4Eu1hA4j2P4Rb1CRbLKczSj+yzIs
RK07V6yiFnGxEdoESR54UvboOjkCCE+9C2sJGny4DHvORpHEE0mCy3Ws96NSAXB4mq12QGUAWh2I
Ge862eEdasLs2zcU1LS9+O0XGc+sGmnhB2H3pESBGZM6dxXB8HVovfR22BV8Z1D7ISrYiFJsE4FA
7XX+02pIqm+RrhrN+lr20TTlbHvvWZkc+yHG9BFwyYSEXvbGWwV6tr5QC3/czkRw88UIrkGvq2nt
gOkkX/Az1BzY6b7FE4SlJ1tZounE/+rJnT84gcxXHKQGlEwp0lNtz6TNlILZWyBZfTvuXR6MrHol
0f7oVotpRDgbsX++qFN0J/43dmJ2b4JUgWkv87ITNLctW0IWHblNIJsQtb0Sz2NH8g0PZpC7nQEY
ZjXvDk//fzh0XfRJLfHBq+YDlhDv+QcbTMZ4IHD+ovCANl9ZMYndF5uT4azOAGhUnNE9ZJK3ba3e
TPQrGzAav+8LieVuoe8xM4+K4ay5M29nW31KnpM/2qahPS30V7vF69W3Ele6LLoR4/79rt+3Cvjh
4yDltH5AdVPXix7UCrrnzlPeXDs2u8RQBApgkfZ4w9egQSragMW4WhKZy4euX7hPIExDvtHZyjXx
wDU00ke/F3GCbwbJBLH3LQkpp5jUYi1dZ/IVZhGo1UVgClCZyHSwB/iaO69iBF3DoZFuwrKPosXB
50cyD8I3ls+qjAIYNSM0bn89a69OCbId1P+YtVufGa0xOae0sLc7U5r2AkDdtLWThpDpvg8XSoCV
tQ+0XviJQfKk4GjddiNxDD+xQ5Xa3+wkYtwS+l0xyuwgHpatfmn484lh9hX9LSK95sbNgkgW7zR0
P9ds5wL8wOKTuW+pIwDKfHZTgOzh3qUPoIPHPnY4X7DvMi8/pfQARJRcMf4dPDjDer4w377WrLc/
ulJx6+IxYatA+7fKUxfWLLan8pemOf3idW6lACHs02jGKInEq27EPIVAhG6R6iRKNhaWNgnPPN+T
QUnAfj1qeQIE7hcqJ8LXesogoZCp+aEPK+MQUya10D0JSmOrh4kofstgyTLOUtObmqfKTp7VGtjY
i65ykpKXO8GgikOSowS0VzcM3N8Pdsk9YJP1+GZ+EGVPqbPhusTKpJGT1wtzXYy5BbzQmng/pnof
qQqHy02gdcFsKT++6yHcJTyLcxtu1pODhxHay08I/yVmTaIROnMAcXR1LxoRcfEFeE9yTnbRGFCm
rQL93H1/aL4uPe6cjc/l35OYJt2m1nhQc0kMO+vMYRwaVCxJwTUZc6pYd34HjE5VQ9Hh13Cqhp2a
D1CXIry19E64BI2v07+JlARcYa4jhMt1b9BuhVvrqBSLYK3uWCLKuEcycj6EmKzmdlXfkY+KYDpL
iodB9arKHbb5cysP/L70n2D1lXAmvaJHNAV/InbjxB2OJEEeg94j+AE2Ze77MgpIPMblXDZyO1c8
67/28HLH8N7yk/Bp2bJIwg6nWZ9yuNLvJwz10Xx2BOZ+yUWm5ISSQ8ydIfl07OmgtbAlqJRiVTZu
yc89jpCTgJ7ts2Uh2laVAqn4DpkLD8QFIE2ePOgNyypdWzteN9KOW6iZK/HROI97zwmiIHbmg7ZE
J++LESOQJrn42Y0WdLn8fbV3G+mcii2cHRHKXzMboiZgnbczPow+UFXDpskzqIEFyPvHo4HlLcw3
opz/lqjihHSSVUYNj31sU80w5321EhOblxUpSm3xluZvwt2VK0N1O+/F2qZL8ucNrx9i+TLR2tPJ
tVn06NWMdKE18Gh4OWmNd/fksaI9880L/RC2FnJN8B/6ugK+WXcW93XxeKiKs9V6K1nQGI6dGe3L
SWwBMdslJPW24byI2OpBwDwZ92nifYQE6HiQPcxXcAWgLK3uOnLRwpW/KB9WBl5XRiCYeRO9VOM+
JWTwgvK/KGr4a3P2mNNx779Zmn3S4/R9UcihZsDX+XYFfrBM8h3ae4P+1Z9X6vdtUYWKXIqgLF6z
tLLWBqdoMAxiWldU88/UjJdGh6XBMFA/Tyq2H2fIKXgpNvwLXIahQ7hwiBZiaU1rGwjNt1GFHVC4
BRYhnooNziNAVId1zxLjicGk/2NvJgzJYw1CICuoRG/hLJQQczqFUM77iML17cYJqD2CQxUQqQQP
mbvb+8UYh4Y0ClETztpnEV2Ua0+zIhK4Nmyv9SVwNhkGJk7I+xVwV9EKDjQS3uStjUslg5CVxY9V
NZcZMz8gu3+vY4KOGVhg3g/A+4LqbuOiHISycPFFX12xg9YnwXwnBpKSqamC0QKbQoMlwQcmVZEW
P0zckYPqnuE+SKDX8XLFxDY40RQmP4P+vh4+wG0v//RyweeBpoRuOyi306j5ULKbg6vNntAhJu7n
RqRXUEyTOrqQ8RGPwLwqBUhu29hXBiCfxJH5YaEkyoEhelDYylisEgycExsLWa435NIBzkYoe1eN
MzDBbtFB7ZmqMqVQCnBhzY0/turAtJqaQN3IlAhJZmjdvu/ntqSioygw9+yHq56+3LMpFpvA1jF+
1DRri2X4YT+xW3Tx57Paa5HT3ltavpzkEIE/Eg+GTqQ3B8CxwVPH11Xtems1wO6P4tWf8ahR+Vpn
8rocKR7Y22PI0m7vjoUS9CUjAEC+QFh6q7W7nWgwikS/1alwqc0WiuLR/FozdOfC5JPqkkbwVib7
zEI/jzOP/cUSXw0TfD2RPnXzRl5kw50FDgQEH5GYGSoWhX5+j+CNq397kd1avDeP9ggAje/PMWmY
dQDwmpNE/8kfFgBuexy00u/yzZCiNhsvt+InYmo/6PeE4TXF0cTaL/rAONOhlrQBeBJbm3WZPD5S
g1FpiLgm/X7xcTOnTjea0IdGo5rpgNWD2n6jF5p87RZ+n6SJGtJ9/tlnnKR20wxmS67Zb+j8m6AR
URk5WoEc2FyKXTX99Tg8Nv5qyfm+qkaRV8E3Zfa64Fzwtm6xeh60xdD8iKKkibhYXrU2OS0FRTSk
vE+ZaTPLFmAh2osfxE7bmJ07yL+uDeMZAOfpQmppNjJaADszxxu+00K2hRr7FJ20ORPn6ZPP/46u
gSfG4v7DfBFe+w5ADfX1/HFbWjtHm2mTogX25bVgg5qjOVF8u4i89ue6oWOTOhiU0HaKUfvKwgLa
Cb0zxsLPgD8pl2lRC1gc8w9YHtNv+uKD2YxHcnls4Iibm4q1mu/spWoN1OwyAWspN1YHBev+ZHRp
5Yv3/C6qZ5+r3wlOkrkkGL9ZSTd8ni0zurervTT02dg+3lLwN3Jfcz7El9fxR8yqV/A9SXxhcI2J
ukrCXBBc2sj+BFsmrZ/yrOJb/akhJbA29+jwUYULY92XryOa7gBeCTzInv5uI0VcIIigWx4WtANk
XB7q9+psOq9OcQ5Vm97hVe381zJfOXG48fyl2whIgBZC8AAML3E0s4XFW4QV/TbrozBMVsRK6z0g
qvaHuAPhewMGbQrIsPSYUX4VBK9DXpkL2LpfrRUb6mZR36g3zv4h1J1hFAUU5Cv6oW/3CnpM1Nx9
cL01bVZFTbv6FO2DSIx/yoa/HL/ZYzybMJ9tsn//HOTrDKIRrLWxVeNqGze5ZVSqdzc/csbtmCw6
B0uqYHuubb8PN85zysPtW9kBQScDbNJaDSdYm2qoIS0X7muzfQ70IZQgDjIKtGLCRYjPkI/bE6Pb
8khUX4vcI6aYHqHWeyBm8SJa36woAxQiTIRXb7BMbDfvS5smQdF4bM8P9K11ogKtbyGq31gZAcEg
m2qX74P9KvujG72s/WtyECsxLywmEZluHvXAxn//f4ja2WAeYiHGcuTe9fKwer1kxpGXmLDeNtXl
tKBIPFkpUvnz6udbQKpLLVfQhXVRwH2TWjYOsUJHAkmPWwEBmgvEqqtd5PZlyPpCV6CuNYgP/bta
CZSeXvqSk2RBBz/xZ/3GmGcnk2UzUc9fX5B/m3mNJ+GjDZv9fxcVuo6bw+mntt3cKWLE0cW8j8/8
GjUA6azL7+ALOgdGWXC49msrxuwjBCycRlOQBLI6f/aaBe8YbzIjsS60vnjizSo0pER6DhBqAAa+
wBXYOfmAjkQ9EikOHImFK+R8inhJ2j2kv00jVxfySHHQgsFDyyUbkZJ6G+3NbWoou9IPgFSBvKnm
xFmnTLFtxFlupOrE/rLUaSA5DzlT6wWhq+Txk7eEKo5WTIuZbDWVLOrRofz5bsbJFwFk51ECisa2
pr6USMHHa5OJWUzvVjPFOTdW7fdYGP4/opnp0wPQTojzMRw3Lv4y+isYAEoDh9f6ReeVw38fFyRl
0WEQkQpphH+btO06Qb56vRYPCWRai7lir67ZAqVScdcG9Chdm0HB91+KOXLWnoHCG1hgPCuwI8y3
MQSi+LYG5WLmLmOWoc/ZOfhDNJX6ci4JkVPxj54aEglCw5mjgYiWI8fnlx1PydiDT1ly9aG20/l0
bijrqGjXhjYbk3deQEVMNhf2DbtDHrVopTTEKaDB8XDIJ5K0w3MAzYK84VcVQz3lT+3fcFPHfcPs
lXRifcPtT+geOJ/lIYLo/j3bgdkbkXKu8w18Jk3C9KO/Q5ea5b1GeY6oHzLEuouBcuKV0lor+92p
ycw9dQ/ytf5/rlbtPXBfBEicFMReB/GFoqa2uS6T4fTwjrFp+JuHZwmOX+v9Smr4ZXpretgiFEJX
AyJA+dTMOFt3rnNo0MJl1QPNyUBH+YIqeLqngsXHl916j1HY3IgC+9Q0KCSvKqSK+64czc22ik+h
hbVtZU7ToqaQlwUIR5ZC5zvjq+ZFafHH0qFlQFs0ogS3SAtRJQofYyDuTBlQ8e8S/o40oqtZ9/Nx
zIm9L6119XEfN8sKU15czi51E6Kb8N40j33XOoN/NtBvisSLY1AyxV+RrOrB9p5xM1sLODsVw53I
S8lWs3P4Suxcz77/7AW1iurvJyOrj9shFzfdypK81Qc3Po6kS2OutMVjCzTiU5IgAcIXjS5P5MlA
GA29YmsLVaLJX8eymwsa21kyVGFzQpB9YKIRYRFWlDtfqsaMV7JcK9UvAg0ZMB48eF0AImCau4WV
zjajBdzBbSbdMFR9GUdcHVdpjItM2UZJ1bw3RspzhRZt2MBarj2ZwLs6FjfwER65jigXSp9GKcnA
uqFp3q0Eg4xig8YHDBIqJsmSJvXdhp7iAE7ABtvTPw4KEr9kfaJELDd13Iauj0scPvwkrRnFOTza
46/h6SjNF4ecxqBaqOaeqOGZQLUhMcPZFSmFNPR90EMZw1nxlCjAHnwUVF3nSSyzsZ7YO0tZrGMh
HaJV16DuZRaxXMMvRCHD4+yRRusqgI6/cxVIFHLmk23xEFRAhjhb344JO6XWmmy8tbjKG0SqnRU5
oQQ5COwjOWyq5qZjMSSET5L97mbm9S3UOjbR9jTooFunn4xYO363VXoeXs/+EcKx+BoboNeln7tc
D1pTYrFz1tsm2se5sb1M+qVCymsjWahGkkHdIV74/2HRGES6txYFJ73N5dj1nT8WTK9WvIk3RpHh
wAOKvuWmQgNbXW8DzfGeajgcxZuIY27nCohJNvFpN6Rju9uhlUIsxUSuP9UGIRgHtnYLxDb+giwg
joUPWk+i2iM9wItAbjyRUchQ7ExeCc+AZjU6l8LFR+jZY0OLZ0UhicscZtBVaN9z19Srx0y5CoZL
IqKU7kERCzKKE1js5Xj1acVClCoApz1AHZWvBTrrOuaocEMUqAlT5Vmo/C9n6sg9B3MOpTcXINom
UplKSc+EwPF+Xx8UCGo1IjPvytLdsAerp60/xgof4tyZPfLVUJ7kXJLwZbFVMyM9+PWv+OI3TOP8
Ib76LaYAsKlYrWcgcv/ggr+JJhfwczl7+NMJIUxUvBMgh//E9EtqpgpI1gRCIeURrMCH0V0u0wyp
R2rVFKGVKjE72H/16HzY+f2GSFRnsfsULsbkZ/oj0MxRFevATtcwdUzhXajKDKTgbRdM7QqI/kbQ
hUe9lOo3Wq3RasrxqUD7ZMouDW818ub69pGExhMJoWSDbK+iqHOCdiyBARaP62+itQgo5Lm6X0BV
64P/Q59hFZaFdMkhSmeJa3eke8+ofNGEWmhW+xzEzr/zNSJUtCfHKrQklzP7ffjuKt+HQSvektWJ
VSUqpCZevXFIrbfQ8hyLTw8f4hHPfu4ycrJLcLni3NF8Ri944QjUBabtsLE6a12xnciG6FV+r6Bi
ADl8ASqNG5vy9ahv6gJXu7q0b7H+9bdpFMBY3jUiRzMfkhp4MUBwRf0v0fjQQ644+ZIh9BiM3z4u
BebC8RkkM3vGYCh1lnob302/qT7nmZ1hfn3LeESzHmL02EU4F8rpgzLrTchV6Il6l7DK3a/Aedou
agd8I2aRbqe5agehR90zolS0wSElul6RYtviupXOm1AnQYD9WyiuunQky6ofejtaVkcgTB+vxE2w
hHVaMFMDM6HNRKe/CqLJYDB+AVAX9LQWI5qoTqzeUiJQiw+l0Mhq+RNnQjxbQHEEzUQfhhngjKsw
gSGxtXyAvCDUJJiv/eq7LRELxnkpRaGbLBwJk2Cr0vUy8thrCkmTul9Uk4pnkXZQMH3sfyKJck4K
mbyjE/xKvR76EOmTfHyMkPQnVquVPDLGur5km9ZuU+U8k6uHGLVUysWWAItBtw5F54IxlkLFrTzj
SOY4tKckxOLNWdOYA3pzRClm7g+rYk/HU9gIXe7+TI3tlxjtrQG/znTrcIo6g5UobDNYC/SB/kLi
fEK3RMLA3pWuO4qLdqwu7+bHUaQlRVErUq3CWhItTKgbdbsi1VRBGLCCsbvpMkUp8NKqZLLZBLxl
km6eQ03m3IcRs4qNfvoexR0iKrlKeXq0J8zcfJEKwysmjAfLz0l6lNYOzT/OxdLyNKbCXNdXPa24
cF2EiIqiPw9ZJ62Mto7WR/crBDm7WswU0q9w6tR8KP1Rh7RntccLsiPRuhBJDExrWu7G0388qmXO
YomNQqeWXMSjjGZgeNfhKShQpxzUqr3PMxgKZSpt882tZ5YjJr5e3B3Xcc+vMwQ1/YfWN9iu1SzW
uQqMbX7nuScc8CQJRSBX4pnFuGyNQVA4mJ8ogEIfyK4qNz6QKaGIkuaVcT89Aqve+MupXE3oBSHy
Q1QZCj9zJYb0B7ygC9qeyy7UUkCGO1SFTFrggWXm99ncECI7tUHoB7pJRG3NOU+3Jx2NQISl+8kP
6m4YvRvD2e1kqBZkh1hDrygn1YtCqLGtgkxiO1DxS9hOFfQLMXcbHWl8TvoZyaaAL618o0j92q0E
KKtYOf42gyB3Ra0cAI92mnthD8+N5NEnRmXC0d9SfxuwGg5P/ORj9NLBnchzCKnkjPM0tFx7M2ay
4QvJn2CoivSGFORBrttf7vO44pkXBOs9qUs03bzcD/UwhFwf5Pb9MeHm4yCnG1s367OLL4O5bjEg
bH82OJozTNauG3w9W8SxoQ2KA7DLz7ZOunRQvFre3TzD0vmaq8mj4Tv5LquXgR3u4//OZLFIbcg3
aD7/Eqj3xBng+YVitz/6djoz+WYLQR7VBw2O5QjL9Bo4esH+5uLn3rS96dN1mK1EX6Jjd8Rt3Iia
q2vKJ3qD5PhVMPLuMj52nA8jckMlv3VRaB2v2BOfwrbTySmgczNzf7LRpYk91fMtryNyC0kB/Vin
+neyzHjGsVFgDNc6bFrNOjOlAF9m1XXf3k71YQ3W4Txrhdiwqz0HhEf2Oiin85rqTVi0YFkmAM0g
bqJNX2wXLBEtJR4kUFXMy4m81tnjdKtgW2avmcTjHGHpo5x5xgvti/Gj1JiCxkguigp6N2xLsqAu
CH1B8ZD8SphGTZXn1NHRwHyfsgqHwx7/ACG5W1xQFTXso8WcAAp+SMZU9LAZ+emd9Bt3oBnilV0e
VElTqqoSKcXqHmUGnfT//+VrFeFaXMpmB4v61ATvWYT+kSZ/CejCkPVFr+OtnV4TDRcjYbUL6n17
kXV2K1tZvcbL1gTXuOR+YHTcSYRky78DRcFfWiLmcxq9JLbWiTflbIz+TtFsGMTc2FCA7WNIPc2z
kBsl6O2lYuQj/dcr8gmi3yvoOy+toWaAQhhHdWQYPkQBYtodCC+M9GCjIUTrN+18ZbBhQhxwtTrX
EJHeob2FMeoBawTi48/zkNMtK50/rwuly5TUZ1WXkAZfU39BCKo3vmuHy5agu1zt7ByAD0YVKkZp
bhzL18CayVeQu0QcW6dMfTpSGJFVVKPk04xhu3u5Gv9PZdiFGv1S0eLnDC3yPEDmgPrCE8RE5KGm
iF6Z3bod7Dwj/W3BL8FUo5nGvKjXvu61tVB8n2kgq0haUG5kxNKlzjX+NwLdXgumezdyj9HDcKH6
5w/Ds8OSuMh0OH4YtMQ9lO3XkmPk7p+08LFKNKgXTJ+JFMRk6S/v82fqtCZ9vv3gML5YxGT4up4Q
KqjZNofNUXSXB8IJyHJWieDqPcY5zHc9ndyrJqxSeZTKuha06MW/zS4Xo4jLX93hReBK+aPr9q7a
ExjDOV34rXsD65wgoNyqp8cSU9OLDGH1LGIgLK1EOE1azXYGoMzu7aWsAdjWUUzGhGXWwaceXSuk
4bAnp0DLqArsRcfRRC3ZDsoUGd64ORwUImbuQhyEcLcx9V9ui91gst09Zz/GDVmXuIcwi0j71NNP
4P7Jre9H+LcNu8u3Xs9Q1FzTDaN+jiQNKV6kuyBySPV84HtZ8tvJjXw+o6SXWolH7n+l1pngZJ4/
u3hMwugNYIwsjXNCadWcpJ3QXLEqFQTvSHC2CxjfqzlNG+kkv7O7BxKCIrEai5rl3n/PWG09mQOZ
aEYKY/O7pRP7+JO3nJW1fsEB7j6Nw2h5pS25/cu9PH0JE1XamSj2ewkVvEO1JVImWlhnfUOG2SCQ
/VRZi7FbhguuAxOHLt7fDe/XZA/X8YRUAyEeJCYB1JKc9QkyhukIz4c3QNAPGdnoaqQ4kjf07B3m
Blgdcc6Bx6Td6Rs9OJqhPks/VZ6FHYK7klU4pujw19mVuu5r4KeeatD/c9j8nLGGZDVsjTcWS0rw
lSa/plshQVz+awP/5zoEBsWqdAy+WWZU+YjL38zLSXqNgPpGCP+hyMhl4hwg+oR7iAKS43A+5a9s
CzR8zB+gNOX2gCZB91nG6Die3JKWDOfyb6v31Bu/bbacygZ0Ss05Vn4AxEUCzqS0pt88WVihRHbH
DKl7jjhIIoZOcSwfuMmnq7Y79T33uMuf2xuBbcCW0kVtV9OBTb0xBykQKaoltJESCy4lxooYp85B
FO8vLaNZlvEMewuEvYzhAnibqBfh6a0C4M1lclm7t0TqPsbTQGNHmXPKZRa50kJvhOB7FqCm2Isb
oIEQuUYKcirEYIRspaPGuisZyRyBWVa2jP64B7hziIx7DaDaO8PnamoIthCU7hZXud7zwKoU99V6
+bTwVub+BaBWfi95pyE2IatAgJIiyE06cLxoBwWmjbVC9OPowCXfE2RNAzitrdZ1ubKRPECRtjz1
v1pRljRGE88a1zEhBhDYfgWAXJ8kfZlxdicsKIP/KxTT3dDiYGjmd7E+ss/cWfiXW4vqtaKLx2OG
ks5JJ7CuXNLfBmNm1WGyjUZ7FZayH6+eCq78c/5Pni9HhgfBa5qNP1qBC2rDNHmJEWXOpPv5ay7Z
V/BEdwC3SFqzSmOxn17Wu9Kwg6iHabeTblwB1/vidf/uYvTgjkBfMP/B8rRYfC/8eWdTpNkIym7w
Bt4naAvdSYcjpPMcO22WAkNXTTMBQ7YqfZJmTjoRfEHgk0zKD258uHYRWcsB7gWdXbDVeGrfkp95
aleLuU2JB/VFUZGors5zGTyo6aDAZW+bsRPUa1vCwTDhyyeDXWAhtGGg0GNiMsvLWZujmXffHTNQ
a0Qhy1Ze6yUDV2A11w4n+T5xgEcCwSzy4Tz0qiMdWW5sOjAm4VzbNXcPVbVQtFk08ocoO1wzU4Ng
5cc4T4jJ3wuXzodAKpOPPv2GMgA9n9/TsfIs1Di9JOIsFr3Kw2YIKSzG5rn4OA9pesShGiFmQxva
lmf73c8Kr5zxZvpA7m1N2b2MQ0cZZ263YiRyDgE746fXXZbS0b/rMKwR6yHPm1kJoFXCmQ+OsCOX
pW9z1Lq9BB4xN+vQjbnv+JznCXYOCiIsB+wTYnOKZQd6CJTT8l9ydUq7flplHmmVk3HUbb+CAaqC
M44YRogSdrahx9OmEfJEpGv8ioQjo8OX/T+xZkGfkZW0RgsiWVZnTUowgs8ZO8fn9vHRwYiNtyQa
cVmr99QVk2lIXPIz4JjA9zX+qx9MoUgDcUrvk7fWFX5n2fWMVddg+01rUgRaMLgK9cRxNGuBS7n+
HP9pU830KyZf7xvU0qyBXBoCmS6Gcrc74Vzx/GYkRFqiuM/PkUznS1GshhtQj9S56Ac0QQvoEI5m
qBMBPXW4jCTvfWbcgOqR7aBfRLCh2NSLB0yeDBkQsU6UDAa4fsPvSWurdNfQrUgoTv5AWVCONuAb
5Zi0pTC0IwaXG3v7T4s4W8tzRhqFu2iAsBOwRxwO/bGo3XXutf7CKKEmZTawv5co5wNpHAOcVYGU
LTI6G9QNqxjZSH5CGjSmmuC3q9IGG6vcFMsrYc/mmwm18Feo3XsacRFsk7tDl/t6ez7UROi7mZG5
gEyTcqF2s714Ur+Kx8V3xLNO3CkbtFqr6DDVU3rtKNeuUFhEAGj4UGV97i3xfInFLZ91hpom/FhK
tCaotY5e3+d/gYXiPfKhsja9eEFLOUIBfqbiU3pLEZuUyN0x3+2zSzv6L4/PR8UM1aLk39A7ro8/
kMAHcdhka9zFq9Z1ifAjWoih6qSOAQ1PpqvHPky0+NJWeL+xmEae7S3T4JFnHIwKPaVPX7DzHLTf
GMCL1Bp6EKQS5Nf86/CNRwRbzqwjQqS8K6T/JJzU4tQwBe6XantguvFo6g8EKYZIrDXgcjYv7mvp
EYGrjmBcu/SRISNG6667K2wLTjOXkV2LaouQ2DgBU6g65H55mh14qbLVG+ksMCr+tfsVHkvl5Fcm
uX5bqvHQsFa0+CV6G8COdq52l+VFQY4ILGfmKiGmoiDIjCh555kb0aIl53mQb9y26X3Rk4miMA2m
YTeNXCon1XHjQKmiZoL7Ob6xJD9vlP0dsqdNj/frFdNNGN3KgoeQJF/vbhHDgUz68UYJjvw3Th8L
2HXV2URkV4zmcP5xrRDJhi7kf7eRu29Zs8JnsmEnMS26ZUFxFAIokiN9YGHVX39/kGl+HnZy5diE
W7i+bD4eqnZ5HAm0ll6SnjTQuA1HW8cx//p3HjCxgW1BgcrrNPbUfyQYVUz5gD1lcr6lC+K7yGPW
OT60U6CBewf8uTo+w8W/zdSvVEYoDOGTNqQ4UHffsCHAIbqdz4P5tiZs8XH8x/EzbcJcBHAl0yQg
tO0CsEpO2Hidckw/MBaBUVJwmtRl3p76anUZ4gf7fIF5/pXJQCGprcwsUtE69/i7ngrSWwuLULrJ
vv9qiGgV4b8TM6Gi8AVo24njJnAfMhEI0XXIHy/ASAOotrBiSdcmHorGPfkl5zCJ/3cZHzn3TGIW
9vsN2vIzp1XrnIAKRPvsE4kwKHo6GwPntAUpNCPLTRGXR+aE077FWRg5/JvXXI6D77izmsHdrWEg
SPSfy+X+ab0SDjPgc/1HPuyrEG59EERhIlgrKTCApdfg2RvuBjoYIR16bjjrElUPj/pqpcIJXeNN
keot9PWoRMMhbJun12A6tBvuJRdP6HF5fzj8XNK0Q+I5m7Cq0W9up1c2IAWiGzaPeeEzyTDJifh6
oWEL1FKw8tf5mGo1ZG1+EBNJx4uRRqVLHhjsTNoFlBNtOPOHeYBh6zs8niK1xhezjy37cxdDVuV6
rBLAhaOxK5hNbAm9Ac6/6FZHBy5uOlni8CRNw2XUZKFkzKOzdqSeR2Ydvxcc4J4wKqVDouBnDF3t
HotQLmDLtejPrEeAF1/WcZP7WwRL6pNNnPUJ+wHJuQrpLrzpbk+RkZmM+A8CGlRe6M54CrEDOGOH
9q4OCIU0cqu4S+8mG12T4mjPoFvEXRAIpv5U2nMV7KnPdO0Eem7dr6wX/dJItNP0ny7GzkJZVaii
E702oNnABAnRVhMv1Qu5fva60Nmf94a8/0N81TF9U1s9r5m7A07lNeMxLuj8B+tX+X1Vfhj+QN7U
61U40NYRT7yXW4fT5mnHMuMhqgL3jL1giOqXXKxoN7V8T8JqBI+McY8ALTUDlBtRkldnvg6i1srE
8ctU0+V0v2sIuTcHfsgsyp287SNM02uNimkqtcAuTYfwWan/035eHQBhOCtz/aSTdMJgZflyKXQs
hD6U0KiuA+094gRQkQuQ+ECjPPRg0gpi44uJLnN2jGMjSdMGetZn4iB35J33AFaX9UApt4eJnQdm
BfluUQNCoWRr1z6Xja8TTmoYbe6WKcWaiCjxqL89auc7Dg8Aa2N4+wK3t6bWdr3l7xMIC61MLgp4
8PkN6Gzlzlyrl89QFa1BTRa7CqT0hhcVC8aShEMG5C2oapuLITigmZgRgmDXN4FZ6SGmYiXn0w1/
LUmZVaI45FoY9qgSxbqPVhkp+VyDWRvpmbsiVjW/OcckzST8fYzI8vYs2bZ43saW0eH4Fq5zxvXL
G2lCyDYAVdo80280po2FM0HGsvdJFoYTVUzwOAhtP3IRXIu/PkWGDiD718eeodbW6tkj9MDW/PQY
zUtqh8Fq5mZrTeE9dV6laM7UDhvryVUTL/o+lfAQXw0gkXebZsUl/rQsePILUxIWvYqoReXxFDRN
xETDzkD8x+tcbysie8BzmaMAU0HK+I9KOxlEf9SL9iN3gNesq7L7QncbWvAPzoKUJNR0rdEUcLyo
fz3fHW/D4CZc4z8wPC0iX6/e4ozByp4cJhwO3Aj9bYIvdDq+E27ItefnMmnhgWYXmXoV6brI4nxG
WPDkreVkdeC5v+/67YwJvWwgsR/4sDxMp2uCD9V7Ti8cYg7EQiSMuEJdPjkI79qaKBwTWJMwtnzL
hr6aRKBhSfMUOQF2fH7PBaxVVRlys71ElNW8NgR9+mr2KcH7Ru2ZqQ9g95iQxwOrWXkJ2ps8n9Ps
Jv841hq9A3fNxPNn7jcMTjgVDsVHwUKfFnP7QpSncFzH4XuuO38Tf69LeJG+qLVCVI6Ie6qqVbR6
wKE/NcJhkJE7GTOC7Gb0VoJYDwhFYY0tHXFFymIP2ELsAH0LrJViTupNvgR8PwDjM6xM3jmsgNHT
KaIn6wHTQjzwJFinRPygUo12QWp/SWsUmxChlJTs8YufV4B6l6wEOuGroAvsYQIT6Mw8aN7I0jhF
TwDVW3gYFpq45QcjU2U/m+xuvDOT5lfHCCxbCqXEMiDioywXchxAHa1XNdBiaM9FXtrY4VnuaSAA
exV4yhoUkq0kMCJdasrBJg7vICrQMpulRHDZcNyrMktRLlCExdkZKB8EVIRGJ5nd/oNp1Rxp2OdB
vRkak43Oi4kxfLDYxeQLMkamiuXMQw6wtByJTQRTyPxoyKieLQIz1j390CLXssu5C9dhExjLnOYd
w2ivtseiWgFv+7w+ByfJKRWiRTQo6GN/OewVcJpl5DSCOQup7PB9tQKj/nNm17cZWIg7EmYtqcS5
pPmQXuSzO2e6kOJ0GdImmEZ0NNziXVuVGWGVrfjgosrC13M4rY/zTJjf4YNz7akJJ/Mvi7Y9ZINy
WL0Jw2FWzargFbSadPeFDPZ19UXIgiC4M5FT/C627ppWHhqSJA2UMbXIP8WgvnieAXfP22uMBx4e
Jov6fw801InXHDgxZJKFrypk9byy7tM5bSr4OXP3RBAV3YO2+odr8mEWDJampfMfaLkRmgGcTzYL
2xFmYkOoS0583AMaX0aggE6930v3N9TkBisSPB/CV/LHSh9/Lx7LSiMssJFHQ7Ju3kPZBTEotkSm
Tcn9/5aEoHuGsicK+FPGkUQpFW2g1hDzzcwWhw9B/C42lANIt7VvQfh5OouUHSxfAsOaeIs6ylj3
9LAfPTteAVbCP4K+xX6Nr0olp2ekR5hD5Y1wsyaOdUmxgXvaA9bTy+s1zBCUoy8JAVHzCCSDx3md
qUrUDZJqmKdm6WDXjlAQ4yo3LGw8SKC09PBmPNur9Px5Wpg50X0qKrWghN1VVfjRcPDigMHucdJG
WdAVNsg2Sd3DeIPdOjFO3xe8YH9PBMxer7r8+s9Q2TX5Chh4Ck2nCldhr0Q2ePJChUSeDqIo3oSJ
mB37V4ROx8XC3+58d4oxNJauBjktrL9dx0A/z8LlZuByj87B7DgoEIIcr2hHkmIhTCkFi9kYnfSL
zL1LC0u5/BDSsrA5FkZQTOXLxuW2zntBDKrLV7xfrdaWyUdyp4/7OK4lnx3pDlVFMM4V0VomBg+W
r916mYK7/93hJJ0AhUT27a8x5Pd8C2nscgCOWn95kuN5hmJMSQzhCc+OP5L3ec9XWYm+Vakp1D2L
+aRBMTcWP/tF2E2hZiQc03fKwrvbBBNF1Zt5spG9Q9rsCRRImSQ/Ikvr3tdz7BXXtHePoqzoM+oB
idcdMQiAcOwCti7Hz1aSTfMd8WGVZ90i6wa8PKSsxYuEf5MVPqYkn8rFmw/fnI19ChopsQSM9DeJ
AuzT8AKwYnwLLyG8xpPY9+e70SoH/Voeu4uMcJuP2ZD4uxPZd9OZy1cByDUtMlI6tGIlDdJmvRXF
5WAboUnLN52iCp2/tOwNvJnQC4qfir03PtD8TItU8bU6R56Ftq1vLqJdf+qFV3tqeHt9LHYcRN3O
m9CAx8Zrutg/eyAIAd//OcX3GKDrs/AZ7fMnN6R9UTejfYS4Y68zG9K5WxHsF5vTy9RMAxmajpjM
PgoqWDnqmHWs0wWxu7UWo0Tu5HAGYuaF9m8pOEbcAjIxG/+1JCJGSDUh1jm1ynb4bb+uL4NenTew
7vxfBD7ymQHUKTC8yvuXCN+1Mt0LCEgRRLYGF4tbpYq906Uy/yabxbZDB8ukD1XbzeLEm6D2W52G
+JoXW30lU8yrI+ZiWmP5kpwewbaXOkvHxDct0uK3CHFVQSiGIi88nf7dHYnsQAYjA21sbyF2RmTc
t8+ZCZyy4lVub50jRkQlla4NoIhCWybeaZBrxdX7FcvReCBo0IKkQsOQZFD99nKemCQIULHF8zyx
oZTB7jzjGlD94RK8P144gaUBEwn7FfVwqFmZEjz//B6DoaJ5WT3EcfWcsgLLlioIqxPLvaQy+GSE
meZCJEF4gKcjq3U+4hxFVA/7F8CoWC6IaGsgwSuj3HzPB9qFe09WZZPga+TBx9m3/BMtwrUGlQe5
GjLImpssCbPubQ+wdMbzIEt2fRP8JVE8cbfMtSl240DaQ65Q8fCFxhm7UQXy5iyhUbLwQYUQzXDD
JNbNPGMoJUhMQG6VQAQIgJINtpmj/BrBbJKKWlCTC+NgU3zXCPuBazjiuiuYfMmC04FEi07zu4KK
gjbg036wJQvDVWZMuiMv1TvbNxDhQgJVXNPHiWx2hGuDPfduHPXAfWadf7Q94xu9hIumUfVne7qp
OA4IfFSatlMI7DAK/cNQeiuP9Hro3pHxol87Vq8C9Es18jaZ7dZTXXQhkQu1Gdthnh+R1IHFDAVI
6AZApvATgMBrqUoSwUKHifPo1ftLic8qYF8h7RZiqgRFl5swpyL5GIzFqKdce/M6gkHZl69pudIO
H2qamLlj3/3i23Yv2S0Jydgo6hdR20BaCcFm7I6SKAekwsLNTM87BKbdQQhYZFkvr79Gj5krv5c/
0gwPYT5F42NzWGXWMtPdRGfmoUsKqoXubcVscrkbEH6YQoU741OAYrP0ow1Pr1O5TkwbNVLs8bU9
RQjCs81W/ZUzUGuBKNy/Gcw6O2/IHlONy8O0LjKDvoBlHvhIjX/rSxmtoIXU1dhZ/z5E4SmjqgMR
FcrarQ+9Tiq4gJdI7MEb8nmt4I7YkZWu6+OFkheohtBSofVL/ASvvUlNWrqS3IMLFzxQJ/99OGRR
RyT42GvLijoxr93JJB1E+xbf7hsJ2GeFlJ/U3m/pT2GMRY7gsrjds+c2QYduwcTEQShTUb4k8zG+
PNbwdwhjSw0tyUxHwURT8Ef30mk4z1ntGVUPRReyBV0XMAzdJES0fGYXkual8f48xwxvf2OKN49J
SRPSvgykytbWTwZEiDS0miKLv9E7CUapKinZVaNUwMBsrA9h2O/Dac2Eu+5LEYw7CVuSOj5R5poB
QKoBN+rRyEZXmFGiKxu/w9zOkziZnOSjB7avsOVWrn6ygikkSUZN+l/C+rSuAfuw88PH1F3HXdJo
Uy69hqTRNetm+0DKSFq1H9fzkbNfI2hmyycKJLCEtfHsHK862DHGKlVXECVTKuDVfKTQfL4CDX6M
Hu84cPDd/pHd1yhJtZcCuuCB8oRxzzYxC5I1V7VWNi6Cr1SY7kPdfoJwa9+OvNpzop2TlrtZVIYU
dY0ie7tMoWNEtmnwre4UR4I8WYDg1pv3jG026kq8RfLFqasvN0ssKmcDg+9OOm7CUUqfuZUaT91z
KjERUwHIhwURNzk2GRidgBahVpLKxGz5eZSQMsGc126Nk7YPEwXVVPuclUfAsTg7W/E5ygcRY1H6
JNAD3dHzbe04xV9CvSetnfYxDeQKEoFbJViCEjEJHxrOg0V+pLLFCwexs0bQ3WKwWemabNn3alXG
DTgkETohs7tOa9wqyqPzUa00JEgRH5Ru6atpuFDimcJ6bCmE5M/fBmnOm/uwJfrxI1GE+9U32mMT
hXuDS2nt7Tu4yjpKKhaBlG28JoCzQ3rHhFNu76m+lz9pgRvBfs1E+XXwdfcXyAaaAYt2S9h7faFA
k6xpYtvlc1HptTsWW4UHKVaQzZRpqEGLaxm25Mezxud0iETh/Fb5JblCOqgAbe0nyF0UO46Eagti
CUX8DrnPEWAsdE3rKUUHLNX/Oc6xQRaBmtOurAIu/NHiUb7sENJo65wudvaFlu1FfgA30kbnTIJo
kiLMPlPapDIDL/kwXyfu/nFE3gawrW/rK6zq9G2wYDPFUkR9g6Z9V00AluVOffPj6hXoFuQ1Qv3u
nciFQC9JvERIv63IoZSIv4O9SztSdZ04ZVa2Uq/HjTCZQGJIQJDmGdIEoDp/TGbCAi5B1bjRsN3p
LXOKuC3WnV3KyvuVDuqMS6dgGIKtej/w0KmYhcsC52sS8oWCeY2dQGiTqdiERlwSQpa63Jw7UrOo
mcTkdjjhiOEkv5lzU/7id0r20p4KO+CCevwFBO9jupAPLxQcDqIM571X7+xpEtI7gUuvOWfgkd6y
CJHdatmP55Ym5s6rC38t3hyWKI5DAmP8XE+hLk4zz7puZay+Lkch4OAusAfh4tmJG2Vd8LbvjJAh
cJ80et0vRFeCaYl9CQseC0Zm/uUROP4CWIpkTZ2/YbgEZjFxedU4UgZ/qDZ3hpODtDWuqRjOvGcM
mmOZ5hyQqDF8ego+PlblQkTZZllm5COhnH2+TGdz233poOT+bJBvrnq00/iEadLIhHU46hiL19th
cmyBNuwztdkgCmMcgjkCq180PNXKcCNt78TKGxg9T7dcheebwng+LcRkWeSkMeucM8nOGilwUurF
zH6i5dVBDimw+DY6Y1bZEbutaM9KyWihiRJRB5m7xr4lpmxHtZU4C5x4X0Oc8HMVz1rlbIWo08hH
yBtImLgrHcqsX/ZSKE8jjvev1tePTNPEpCnvvovVZloS1ey1CF4fYXl/10qOCF/RK+xh/TWlGuSP
kftMJHUnbsQRKe47OAUPWJIomi5+5ZO3NmPnpn9B/xaXJ9ipSEBBL1/CITIX0p42e8VtLnxWgi+n
KaQdCf4VFme2tHG2mXs/5cFG2LY1dRLA+O9XuY8wak1f2Q3Vo9feDyFCh4DCLLAREbecv2gLOofS
yeULzD9QF3qdqoaFyWesJbU+ExuBmoG8YN+9B3+V5Yu/czazrcWb5LNamzBTgMYmlFPF5Y9XfulW
gk9f0oL9xltr7MKz2opRKB1fD8vDLU3z1RBkdJU0ZibL8MhAzi+hwHDIreIkqtMyRJlj+DldB+pv
ZXxtwWWDlriNv/5Ts/fMmAiuo8GWOGMOeZWslOjdzOmZe6eQhNtg8ic0nDkLPzMCZVHGnYTKs13t
uqn9qGInStEI/TbPDynLfnEZfy/+2m1pqxAEVufCx9JRtA4YuVGPU+MQ5XTkyKX9BN1yzJlZVO+K
1ArUMjN1XU+L3s8jZfkCoXmICzoESpP5CHP7IZlY4jF3tbOmOutvsfVyAA49w0hLLyX5mefFjeGp
+1aneCUw3bSW7+H4y+UH1LKT6bNg9X92YXPDI78uTPjxfYU0BXcAUy8oV8HAU+hMsYfxyiu4IDoH
2zdNnmpAxM7WChjXBTHQYRPExnXuAX7m+qfisL3XPKkDPm6mKx44W7EsusUQIIBRw5nUbui/CFaR
vbHyl7vODqfNY9t9/Feo1BmYHPzUQ2EJib8Aa5h1Aqw5yK0b+tYQp2/0sxHhAenRuGfZRaDo9ovF
kFhLophqi/lV0ae2SHhWPcbjjMMI7fVbDeIQWjoSs9lu2ljXguo0i5Bw9SNFdile452YieVUYKBX
YieR4jsNoBL+gcxojcpRSTsqUHHH4/Hcsq7/7fFq9Gkq+S0HMhkJV74IMWFl66RR8YryUtIW6pPY
u8WBy2FbvZ1l48908ydz/kUzQn9G1D+FYJb3NVC4FRnthCXehrDSE+fy1iVaoT2Uhnfpm3UuGnzf
4X3Y9e3uNJMITILWN4jcSqWR8ikm214qneczU2lyKZQdNdyZTwG9lhw2SRlRxw4O/2CDkzW64Not
yXVK/w5hqvfxhNhDaZIOJ9t5GcYWUlgLY3odlvnspfEKuHCK3wrvPYR5VSwvgCWXG5YkMQBSsCYC
76VgMqf2JksKNuevF3IfnuxQ8Xh4cg1rQaWdIivJ9E0q2mAT/FMuncKWZ5SnXaApnNYD6h88NFn9
cRcNz4er1h4TsHu/ZZbMhMWgzfrXZraTeJkDSBM4qgnQ9RawZPeqQQ85rnrrQ0eXdNYW9/DMpGbH
wtt4LSQBExvi/pQLaA7N9IbPIPRBJnQZ/g9AZbx1NkKmjG+Qx665i+li5uvxZyrtPnFdLkHGMw5e
M4SwJ7C7ftZWa6qci8tdLAXFwPfBwgHo6Xs0mrI/2OmDjoYXbwHIHRa7weHxTJwbeBow49kKgax7
w86MbPDcX53f+sCytjXsaVHPthT1Ya4azNhjhMv5etDmyvVkwriXXQAJglbkQeRVzXbayZZuTUSi
NhG9Mq+3AavRmvUP+til9pMCLTv/na+cuI+KKqRZZpGlCYZwRYfR22bGPWye0tJcCXt4K+62kHRO
eVg12GnWLrwhmBahKW0iEpruuyRoQ7SNPYc8RXS5wq+p4VhhvXFKD7ZK9jp3Z79U9EvHhy9ViL+L
7VRyZAlTpzOREzeLGqHqsUiA4Z/OsxCMva5fVGZnkmjunjuUvdq0IW/8VYtqnQWGufZUMlAGp91S
uibEFi+6ojSS5yasQPOkvY8ok2mfUlxDp52x7hH3G4nGl1GapEyBZ5PsLHntSQbp55MTN+/wLUDj
iXDkkBjzBX+23yTPHEp9gRwZEm+kipSYjN0iVVH606C35acl+RSYvIqZgWyv7rx+EwpkP7J4Rr21
vWffVj8vWEJKwtcFVMU0b2v7RkqUAhKDzbGCulfZH8qJtalrm82XiX6Jn9uAta1CLoQpqnOZUTzT
sWnwPGZCW5dFEXmhWywRVvmzChjzBGW2920G7ETKJpfFJQD2mGN5uFAELeE1yNQ3WFRP8pmI9yc4
Si21EpbWHzHgXTDhbxq+EPh9+u7CU9g2WylnqNAJuXrKC5x8N1idfN1J/6eOkFawQVevd8ROrV+Z
8DxypFfPrsNJwm95lE+a/AeBy+lNl26PVH8TpX3TsBPA2FcqwrVXyK3KHJ51cRtHYR+Q2vKw9XaI
r0NeVHpo5OnOL15Mu1iz9ypSqJV8sGPV4nzd4kN9xh6CkoEbMQJj9lF1a4uUV3veE9htnYmtUoVJ
F5W7zD/9rmuSqYfyW8E0/vetZCXGcR94A3Euhw+kw3XarYffaSdO3SGPj1r+0CvZmclqLT4f5sZz
6cMTGXFEemrmtzbGCZJ3+N73rhYdQsVq4uTciexv9Fy2KbWKBvlSTBgkhjM9W+uG4ZTq/xkftpbI
7my6KlJmwvN9ADksaudKwAo3Ai+QmzDPwgzlICx4p5vXZZWvL0IIlWL7SYsEKkZCyBmmnn94Z+Dh
5cc+vtAZUONg/RKbabti2Rvc4ICpqQhFk988E90ZUog+NBGfh4lmvv2FIKIKhRjFt2vKwJekZa0L
XcXlo6UyaED1Bv3o6I4Rkm8Mn/qKd/4KAxWElEb19FBlIaHFg6NIcxYnKXMAz4JrWkSR0T/CJUN0
RI1Ph8iVqsdU/CZgiq9BeKKTVJp5OVtvzZlkKEwaeJ6oqEvc+hAp+yicFilzEWQNSIbdritk5ZN7
BOF/udQpFWGx9vH0S60cEW4fwMk9hSPXHrcdPd2vJlOb3foQ/wo2QLIFRdq+t7+1UJNDo4tgBWCH
Ai3oBYisHmdf6Z2nPFXiXEkTigZvKXaLEnai/GPhLvhO0YTQPKLTDaysj4DKdItV6adHUjvIpTYA
D+4ocxnNB3wJ186BoqlgmSIjIOlku2gC4dpmlxXAO2PyaYtephfcbLWvUCfUMxbkoz6d7pb/EhJm
fQcA/jxDauB0ZTIzm1f9XmaUOAP5gRhY3bfeUJjVp5TV1dKrVdFQxnuymAA0qxE1nwO1P57BnOCe
aakweiMQ0rdC3/3i7Ki8pggffmiDMSsn/F1/YluhatzBQYcqynr7NeyTDO0U7mBZXrT1o8hWqOWu
zq/mUfO8eBRrVNspY0Fx9otGereky84sjaAkJ1qQJxqNYq9WFAZ2JQp4m7PdHdm0F82UMONYBL+f
/Ca1oFgw8XQkx6uyF4u4PAZykU1bM/2ZQ+VuyqOQWjW5/LpyfWfo9nKUJGpUQ0zwojYRA+Yac9zz
vZu5Y4k2ybKQeml7mE+OoY0RWPDIsxOkz3NPZ8MWmptaAuecytskoZCvTrol0J/LQQVoylyY5Hqu
wfLPh9/B12tuGHV+I7iKoZ1egIijpMoukruZ4cRhaudpDquW0NxeGn8/NTI+u9JlRGjOuQPNVc5F
EbcwWdQmtQeoGu8Bsn9flfkeGKZaoB9IZWayE1KO/Cy4kdgUVVINC1bJFa0kqfKFNN1ghwl3Q/Ln
nas/tYxz7/fjDKrxqNeOTzJ7Ir1wWfymfRPDzoXCgDzFFBlcZixJQelCpKcZdvI8RxsUbr81iyyu
n8FAQPzd7DYEwhtylp7HgkTyiKbnnMz/rv7gj6E/Qj3IqgYPzz5KsQiPuZV2Vj2ezIZnAET3d3zL
VKYZyz+L+uzXVHfdSc/NJmxcS9TPD4zVJn07vt01J3oO44uoRHqfuWiRpA/i7p64MfzeRHOUxrbc
NkgXO/ajmlPeApmL//0s9czclU7KeXo3No5D6UVYXFydeLikTaCDb/3eOai3d9jMs3od2irnfd15
VQvdUscIlTkMIoFEUpJb0rVX2LrxxS7SPk5AzSBqUhbXlWgwKxXrLmNgThPr7wezSYNANzriaDWE
sAOv+WfMLfrb+kTShC2tFOJcafS+nXISUv8lHMyh4/wI2DqqwSIbQ+ghz8Cpf5T1tfYeXPUGIKmQ
c4BT6KLeXjZOM8XgI1dmdTWREN+N+AAQVrNa1iJnCo2HC+5Rpb6r7PbMhBPlvQbAK4nXF7eTDSbA
8j9m2z1JYjG6rcBXMH8L4vyDQgNDE6TU77bNv6tCNxbNxbROiAVfZB6yoh/dkkGebY8DEMOdlIRV
J/H7hAHpPnFGsBjX2anrAHAoq0hWa3SqTKiN0dBc7SNUelFCi9LbkSYhf/vZnBFnFL+oebQlsCK2
/sInZqqF0YLXufkkTObxTHCsfpRg+Ts4W66NWbqI8uE4XbwrA+UXGu+UrnfcdD12F4Jv7K4TXJZX
gQnzptOSy/ge24tDEpQ6+FHDRG51n1oCQvSeBBxFTaqKQfBoQpU22cDoq7EYnvD3qNY31iHpOk1s
Ksag0lcXUj7+NMcsma/9/0/N5tcTXzirx6eZ8GL5Ok0cTHjxhi2oEjsL74YAnI7XieeH5WZQYnQ7
ayiVubfwhdKh69bNWNHDUOo3ItoOEKVDGtSD/79Q+QMTw/qRAPZqRd88DsA//UcOqfO18v50np3E
ocrSpG/SU5WihSApmB6WT6+5VWC6V4rP7aAw7IQ8uhKrpQRwjfNfJyOL3fajY1iTLNIbT9wsDg5T
e1p+889OrUxVIaQ9eowdGb/mq0yTrPljQDVD6xrUDgKx+5ZGJhEvvCeDka42st/HQWKU77rpkTrO
dhnPbWSnCC4OxmQQ62ITMJxK9UVDyNJsTDcvhoPnbwlEVRIMTVJ+tbhK6RO40Ns2YDFF/Yj3YqoM
VFlTnWupdkXNH24RCgQeKODsO6tIhs4Iv4/s27JvW6ZROKGPETQrh7bvLLKfIzYbsDcZWIBtfQrn
j57GPdxDiP/VsZji+N4riGnwG2hkIAX8be5m+ijehPs1/2wqlWFfc5+ioxgEjsHc0Y1ALUXTKeDC
awyBTk5JfW+siy0YgCiSC5yNi/Vgy40uu8YSsXx4p50WzDN/YD/YMkC5kDddVrpUezwya9M0nNct
eou8uVRVzcgcMmNzs+Bdqqh74pwgNOJoOiNDRVLfw6KdPCa7CcpyoFuxafe3K/VlrNa4SLD0xICT
MXkDzQ4OZn70GeAKIXpHFRbicGkqVY+bY+At18kXfBD56w71xYcxkN8pGvloZIvZEw+w84P7X2i+
v2cfwcGeWsJTd9O7MTj5B3if9l+ptS+0YDI0DUc8RTqZ1ShQkDbBZC4X9U7GIJu4GQ8FEc4m5BvR
9f/Q2lhCETuT3Eab8ttu6rG+abD/kNXxeFMx6+DRxpCQRVNz9RXnspncPCufnwCxRWl3BxvgbSDz
2S4vanxM9UsYluV2bVsqzhsko4B2xoTX5lngcbYc5+/Hkwiv8489PGdu+HhnefdZ3zlgeWg/jK1W
y7qdkS4+wOOnYRZpCE0C+IU84b07SL8/abQMGP9sTVcQTzrv2jwJJhYpZP2SbWBekagMn5qh9xYH
2GcUONYxCnD0/5xXbOW4mhdWYQthM39XOQckt9pULQ0g+cAyScmB21a8ns9z7uyhmKBBvxDMp26G
jF6JtSAfcuChW3zXcozdUrvliv2Q6UufsNcSRIVJuQXL1hB5qFBcRFJgxXehLJgu/aOlXdEU4WKV
SKpm+Awc7J/FjsPf7aLvcJ9NkfW1AQzOIImcvPfCk46NfTnwueQU2JCrDbozUUVz/PvC3tDuh1PJ
7G+6Q03UN39KKMIwKd+ZWtIagkTgeQZefbG8jz3OgaPAXcG6KOHwQCbTxUSto25vQSeHWaKy/BcH
y6FMRWFCojdmhtkJMO5SSgEZViwt5Gg32mM89rhH3X/TqLX4RmUq5AU7FTG0sSOghFJovZnCxWEe
Dal9vramkcfQ7PDHvjqMTNuaqabZXt88UOsB0Lg9uJq5B7JQ8+u9fzJl+KrkKrW2zfIAHYYjijue
QCP9UVJwhRpA6pJjzIubTvkfqb3O4s+kkr+8JIlmV3XnN6b4ZI6sLpKcEBlGVy1VWWasOzn1M1i6
U5x60pb5SUmQbnQET93vr0cI4UJa+q3oz+6OBbcaelCzIGr4tr5okr79LfPbBR8Q2yNUrYW0VtFl
8qkTCUKtfUnJ2AlV9np3B7EEq1nUY3aXBqc+KvnJW82znxwCf3ebg0r/GpTCN2NgjLjUw7tp1uGX
Iih6J4YO4qxJQRCgkVNQhafjP7wE7dSOTZWv3JUKmdQeJIrDkTpdMuMlTUyjiwkC25BQGH50GAaS
Jhw+V884LK1cqQlggLmweU5W2/FDWIVPOILwEXjyd0rAdLqK8pzwjVPshjY9of54ov0OwY/78ldE
wROKqO5FyV/i1jRLhJroSGPD4tlE+EuuIXUh5xoWM88OANhcWeiN0xL7eEWEVOxT5iMLE08FXhfW
KUFjBCQubig2cOSa1mkYr9t7FaYjNkv5rt7ib5rdMy+pkSprTO9fvPH/hwjosLzAhrhb34SkdvnJ
HQJRwNPAnKVxtnPsqT0rPLZn8JzDKFo8E7s4W5Cf3jc5jq9rGk1CgYtsPjQYkyny+YTAO1IXdPV5
GSLsjoacw1uT076QN5r6W7S0qSrNX/K/KkueyhbGXRXrQfUPj0yi0oUo0TyrE5cwH8WmjDk6W2jY
ji8PBrOdLhy9jRxzBZ6LuGxDvlWqDJujJ30i5TXz562LVX35wh3CI2xn4T/lihjOFiYUTr9SQ0B/
2Q57vRAkVw47LImvEkyvyI71M611OSlh4jMlBiQpFkPjeq2mdRfqyElt3TXVLxQIIeuHfNQizJof
HsO7cdWmlpg64IhF1iyevyvQjM0AFc7AfNsQjsS+0GOD6f+FIjQo+2C9tGvnn1RXIAWqjIUwX67n
bAL2VLUl4HvkGmaf+hFtHHbEAQkSmC8TqGomaxemP6OFsYQS+MLaq5sjYxSz0KT0XoIGkHLWx5l2
aNyUe1kq+5sOVbs2S7NLV2MGAa95KR3W/bPoxuWZc2BJZmxCSFgEfrI18+q64XGQEH2SLBCiMlkC
OSswTGlQDDhJLyvETFYsqy294Cp4ejxXf3CZValQnCPyRfwDOtXax75ZiisyBKbYgITwSdaifTbk
l32pj3Ocv5Zpl2LaWOVfQmFYi5BA5nRHc0c7AcYGvGWJiJNQB/MvSdyh8cYIKgcvjRw+ykEFrcGW
0M1Gtz78VRKSok1eHx7XjN+RH5ITY9wrvyvMKRV7EYTvUCMg7XmWUAV3l0h79WkpQAPEC0uKZ3TW
FqQCZU29SO/oC2WNKwQMDN316Nb7cjmuKBD37+FtuaOK8IJ7S+ZjJQFv2UoUXzwEaDK9LeDbU5iM
Tb+C/5RsQZ5PKuBa0tGXiy2hNcsPbwDaLbIkrNzwnBSkx54GrWUeBEC5ZJUkXyrLK4Li2n8xhNgT
hYis1SHlTbJ/JTzoiM66i912bKkvmNUczLf/greHQhqrlUvX6LAM8DNXPs5/NnnEwXiUiang+TcX
yNflRgiT6CWtAGNSswwfqShTXl+VHgBZ5XEOZl3pTX3aC0KhSePDE41VFeDDponl76GHp3GsKHCP
iA78ijm7p9x0Xs0T5QMVgbVOVmxUW48ipTIqnjsbCWVzT/FB/c8JI3a6kjJLJZpBYbbK3vGcIDCB
aLQa8HvAAUbApDjvBySTSG1Ok7iiRlYahKzakT68BpeaX9p8WPQnaBAmJsxoMn2ib+fqYwYfgYQr
v3/ePXoiMAEFD55i/FcWzAfAQn4TifscDaKVt03xPEuDQS8B417ldtMMw8ArOPvJuW2U3uESAYR6
ZM4JZkcpSdwyFQ2BLCU0AzEed581nnm08z3JTYZAEtiLd4Ao7ohyT18h1N68FinafDnW2X5aqfRY
ghPDyVs+YnHTKcrsa8S7sAwseJbJRggjljSm1bGWRzilK3BFtryQQ52tzuflqmqgBziG+lWmEuBn
Dv0ws7tS97R/ZfH3rkVkj/E74+9oeKpsNCqCCr//v5s6VF7ZeiVcPm6IRl/00aNFSF3+LRuc0sZF
HF3gSs8RK0y0BCn/VFBMCIV1ojD4lyKOMHozzfHwKJ3m5fQArRlezpCx6oZzjvPrBOiUqfnC2viU
TW8erInMO7hc6C5zIJzraQZ9UWEA62eTawZj0LR0gqIDBXBKW5JDBmmWf+S7c3IOSJ6JvRfFVPd6
yyWoW9238E8TO9QxlKMhEsh4QpJv5KPnhSLLT9OrQAxI7e/WKV30rQX8bKHe0H21cyAIUGrlT5Oj
YM7Vy/+8hTnSKMLu3JN2UPJlIUdRZrq2JbbTgsDiCqTOGwcV2u9mFFks7tsws+SYBdwfZ/Q7b56o
HJndmZ8vyJ566Mu2qae15bQODarHcGEHkbJI0g8I8f2RqmdLgh5vPkpDzIYFnB4V8hvvMZCoWF/4
9YSCW/0hGBWlT7HWc7kLlJgpKrSnLNGin5kgpF61sORGWxafz0ZaEVFAxA5fvl8ovbBZAFSHn7mX
uTfUWxK41xRq+okUZqWc2oE/dHiczwvoLqSiovXPMG4fsjhtyilTi4fKtgVyDmuyT5yvjmAIW1oi
lQvVMQiC+jeyHgSTy6xz13wyIEhFOdMyjnz5kmAAIuKl4QVHQINKH2lDHclRlJ/t2zD9s+qEg2k3
Fp94uGYPR+y/aFZ3IIxq/ew3yPkDuAh9XywvZCjPw79ATkKemODcv8jIFpnO6Eehm5zury2wJA+u
6CRmaPlO0ekeTMGq4X2o04ZuzE7SLVuGGbhdIYgGardYe8EwlrHD8xIrHBJjVn+X61Wgw9l04pde
y/JFlCUNDCdWD5zfx1r1a0vmcgpin7kHa3LpE+lr0K1itk/I/SLHmuTzIixDOQq1jY0+o4CrfSA2
orqzLjlEz77V+ToRHPVcHb/OkdwuAGV5TekngN2Z+5t+9c+Q26MwTqANFdRm9bg01nEQHRzy1FIP
TdV0Um6CggQVuM0PUKBw0/aWp6BQwJlrcGbvUHYtCcC54oUTZp2PhtbDsOKU/N5uq+B2oYAQoSKD
5aWlZIdtQgvj8bJkGRTR/fDB6vxVTiHUz4kVawuaGwClb0TD+jh/U7GUWgSGNDDwfEjs4oCR5A66
BLs/L6+OpRNxNb2loROrWfdjmbHdwlhOloNFwtlRnYj1aTLK9n1Bct7wcAKrAYFWPVDD/l3vTnaM
Uv9UNyb0ZnHz+EL3xx3M1uswbvPcLN4OJ8NvT4Q5rrClK1wrZVOhFU+PEnpA0JJLW23mwiZ/wvMz
NOi+8Fh9gwA2/aY/gjNwO7p2TcTrcgZy/DHKFwldfPpE9rN+Pa4pAwitIJAmqct/7s617JJ7SDnu
qiCDyotGz5NVX8FqLXYx01wqdGwmsjiASnMvnvUVMLgce9Gp9qWNmi87T/fcp9TbJ5ccHflorrew
w7H8+qRnrIHuQlWvOFqFH+fH0ROfUbSlR+TesTU7F4I7TnCflSUvAMVjgxJOpZL8SSF8gEjysfXQ
cc3OzBa9LwtsIaaDH5oW85CRkHiT67TSp5m33OVVrJwKW0UGJ5ZOPv8vZihQpnwXJzeYdbShCMIx
3pJJdIvda1M+E5SP5sBabCb/By0irBCflxld+B/vzVvkSbd+nUGCFM781fKkRqP6rxD9QIRjM7q+
+SE3IjyoOMmN80gU8LXCCnd/6rmdRmF+lrlwGWKuRzFYP9Ji2JI226NI70eHqWd3qKnvNYQjj8Pf
Gawoapnb+WBkOw0ICJxQGd6gooZgvRrJzX7P1NESs8k4XpHICepIwRsUUpRY/uVXEHsjzUmkc/c3
ghnTM0Jw7cxW8M4yjzmR4PTn/O6Hih+pNdrVlDLwLsezOHa2CxRSat5O/jtw0oKvY+zLEY+Um+m/
tnAWej4Z6EAZJ7AzQXJ+I4eW96s94/rB6pnuIiXK6PIFRewpESh3CS5/d+JJ3yVUodf9psW2jqEV
+I7ZRGxJnQg7kDypuyVZnxOoRXSQZ9ZOeeuRbaF9jMz1jOy2ecjkNn0ZNgvg3nLarHJT+anwzJbO
mjthFOIQDAXgsx9DKFrd20yyQc7LtZwTOW0sKQsfALNKBoUUQvWPB6dKg/dHdwXZ9xkfIrX46qfa
V9h5CfE3+xtVWAmItNLg2rtUw2kyE+HgVdv+g5pL86wxbuTW679/JejgrhSPADBrQyCZUsj3fFFG
pxOsT35B3S2NkCYF58lpik0Bzk0w1ihFNG9bHHNd8JIvfUr96Zv1bpCubFOTdQCFVYE2PpvikyYq
y7CPalgDR2TPXJXIJc1yEscnfsRi/5MJyifGlqixD1n0DQI7WhtVaZD+J6kdk1ZqS1E1s/W17pvh
NujxtChqlmNxVosADZk4K2xn49+mwVJ06iUZo89NsxgSprGFL2OqVuC8Kg8Js5Zz/djQT2b/M8Su
cWKLeUfmRUAzhF2ylYREB9H3ByfxJBGtvuGXqyWXO1UtxYROjJkVtxyq1vBiUCt05ZEz9+taPS5v
6He0Xm8GXFBit2zUec+MaxiSYfBU20xlqSrh+4kxWWf7Eoy5VZ3T4FziI7dR+E3S1UJfS5Dv1knA
QWQEfY3u6yv/DOgSkaf8SlyrbS3g5VD84LrojVcWL3QNkUs0EMztY4KEZWHHJTA/Pwai6DXQsetC
BdMtaXQ9cUotlK1/HT82oojAYw0N4bheGKuu4Zi3kR52eo3ctmlcW+4mqgZFHo6/BxcW780OYi62
47qBh6SpseQ4xjEvAxW64aw7K8DjGfqRkvc+IOM5VSvOik1uV1af0rKWjpnKCyO0bQf5T/pCa0jz
467rDTEZfGvw6MWyYLU7Hvwkt5C3HOuyGY8F9Z5mcljI/QJwSgiDHD82z8HTmdm2X/jCdcSE0aK/
sMMZxCZpkd1P4R+RSUNdd3pIq8UZJoMXxUcGajp1lbYHfFKMHfTIc7s86sU5oZyzmidc+nF+BHmQ
Z3IUcxoGWFAiL/s2EqPcwt6dwsYxoOY2JazvbJJITgS6usUrT1JKWuoPqo+L90oJMvR7h4+ttnLr
0V3gTkzKqQ5FqKrMx+zFC78FOJM0f0ceO29Y9z3VB3sOhplSRoBSo+IAcsudtBuzMvX1yL3Fd4U0
V8fiyI9NdaigsYbUdqewuqp63mr56Po6HYDMQTmNBIq9KcIxekrz+BNh4r8pcBw6GTyqlRPa6ZqE
aRH+eoPRQ2wc67JYMk54jiI/vdWVESuUzaHBGgy1x/E2HL+I8hv+s0TNjrVcuLVN6hUCjzS3NjKQ
b80UBpbUipuxIoMUZjD7tLJ+moKACG3+gWgBrWpLo53GvhvCiBt2mFmpCBm/7icCbK89E1cv9OAQ
WQuodOofsAHUCtrj0lnenQ7MAR7rOC8HsF/pLgmPYMw7Pk8psEGBPAHBHgSdzQPYfpYDz96/NevA
AWbY7Z+s/Zojr7IoRX5ToS5Oxtk2GqhmZStSrebIzejuujfdIkEFc8dQts3s1RsyuoYDQioJrL03
qjP22rPq1wM3rk0wSyRB/dvN/qL/6gwLoUegYKDgOu9fClKpItQFba1ufCRNegacvVuCcZXeRofg
JCwuiPWoUAxy7yg9Z7G1pyvoQHBmaUOwdQZYRTLhPBrGn0HTFQ1AEhsCVVDspU/8GSymXK0y3a6e
s0U9RhyWVrbOLEtCHOvshl8N7U7d8aoiDTbZCduGbBA/1M4n73moXDPxMxXjEO2MFQuUJ9iXDy4u
C9jRz52BFJQmkJ/gGmA+Ou1KX9StZ6S/GBGehcDqXodfV9Jt2CSAjBdw0mSmnGwccsTb+yAR5LdU
/kVMW34Qp2N9ejXjIu989crz3ddVjXvy5GwYOKrO3n8cq0KW45WdTrd3FPrqB1YplSlhgg5D40X9
k+AlcLeNJVZVAV2k4mVIdNz+PeUQlhn650fXSPzsfj5y5fihEC7JEimS0Uqgu/pW1CH1LK0sLL59
tuAZOfUVznJz6p2rBT3C4sR0fswiM6nEtQsIIgYiozOiCVLBjK7mONFKxZwTBOnXKca12WnfzyPA
rv+yE6T5zihcknBVl7XNQolIUOiX+hw8IxK+WPWVh2JVGfNdEqPzSurYbt6IdDgoVKZvJBqPz72p
yycCYOyrp79YJ0tKpQVuf4vXSaWcb5VSAlUaymJuAAYVwzM7LBN93UP9uwoQYIVS1lrJ3P3Stj6X
aNgU1KY7aDV0zNcjqOIBMVHaSLAXBaRFTDDuiHbPs5r4xJ5tzPen2UhS5/wZxcDhze3XDLH+cfl3
kOhC0Ld6A0gDkjq5YDT1fBXueasiDTCsNYiOYvT07xsbOUT5+jQkXFsYcafu+tWpSIAfH4H8h+mR
y38Efijq8eP51Czc7DbEmi9mbX7mQFbm+53qvEpjXjOtQYkT1zYtiAQG7R5mfGLJWAWYLxiQtgFI
4qgWj5hQ19XZYlkpX/X8RsIbBVJpOs/MoW4U7Jm+Zy7gjgUw8mI/T1KsVqCvK4LiO02E3SDgDGas
aKPLx108SCjOSpBG4Xa8zzzXiijwn3pjO+FXi+OCcbUUdH1b22+1XO4DB6eKiuDXc9AhjH2/ved8
9ekLS2xQef52JCz0ZlrP+QyOlYIDBPPSYz5Ib7v/VSHbL7eUcaYDls0s+tp2FSiL4ISZqAu84XXK
zqUtDz3F+sZoFGlwHbxaw5GQVTan3mN9HDSYvvtspyjnQiw4X6UaLnq9fHhvEli7OkhPJ1mMJxFE
lxwndI8nudeuJQU/i7wqFJMRJBLGmiRRm72JK9kHWm0AULDI2cQg8UyUNYNTcwr2nySX8nltxGww
a8/YtUaNPm47tQsUdI3jAnxKp1Q7E2+Gjme5VRTnNDM6W3t3ecX/9OWT+2pCAmpmAfzd45Bjqj8B
MfTfxVgaJjuoLB/V501T29REPhMPq2TOYTQToz4EiWO743DwmLKik+sp0SeXvKQd5skd5kiOSUOp
HuLcfpqIdDIyrisKOjKkxUFTfWtKXRkT/liVr7YP7LvNtAtL2DMnAlUrg5uAnV4RJznsgb5FAcxJ
GPyMLqKiwq1ENGI98JzQXZ4G/s159uiQEGRE6LF3zgB9E0eXtxvf03Vw7EtJPj9KYVGw7UU79MAe
oFuwI7sBUEwrBNh+aqaub89ckQietjQ1STiAFYF6ZkHY3X5vfSGtu7NcO/cECUJbXFAp8F+Ptub7
wSfRSSPF1BeNQghLWLHxjZs+LL0ArHzml6HyVNJU679Ib2fLIxlVRycA9wb6Eyy6D+lwDwVcAzk3
yW4cxUp4O+rjP/Ln66N1OXaskpn4Dh0TcWBi1JKJtoTba4OzWtNralq2QlhREX42Yp/y75iLoCM8
9hghmO1b6c/S0TCshOYxx5hh+JCMujTmE24ACvkwI9y0tCtYVYRtBkpA/U2phff1q4u/ewOfckD0
QyAzcayxJMQRgyaFlNXZQA5690jqZmehImGAfxTnPEKCVsMmt6mDRVyP8IQu1aVZBSJbdIh43Dly
bRohZGU+f00N6WetPQjCAE5msbiGtMckptHjZ+CZ/4SauIZPNx9O4T59J7Pmm7LDle60pQYDRDAF
MGqyeDJJEpcNOl8OZ0vTZY5wQx7VFJ3nKJS0XsEkMJbqrL5g04Iea+0kc7WK29T3jSv7ftDoBa2n
5wTKYDGSqKizRc9jj1+BO6CnfyCly7He5CXsutQlSwOUiFR/zzytbKOy6wOyNmhECBLWwgWUMUiE
C7iTI0/gFGhiwQnveVAWaKqRamqamzSieIPWfcyOcZXnjzGjteyXUSMwoTY5F1zcVZ6xclpBR3mM
XVyrGVsmmqCGm74tjbCaqmfTcC6RpIG/MJuoOBBIX6eMhzo+JK8oBUZYDjeGgrcBX/mWIo59mhGE
gvMYVARDJL/CEsxJw0b5iJ/1F6vSGkbxJbI+GTBz7pTfMIb6GJF7LugsWAV1XgdYleMD5Pzdq5VA
0mphoeT10ovDbWCpu9LC4bo78ZuJUigpSn0SyS48XJUZ4moriWT/WTkZDUJzttWpEMO95KsIyZeq
9HvqcKBwHs0xJH9n+Sjp3YU1uaE0vY9jiF6+xeGuYk0J+TiApozQAmDrFNp2tQTXEd2oIEW7xu/v
05mO4PYTABIBt462Zp1hbmyx6mA00bFmjNaYIafbyf34Y6Qm9rzx+RG2SsMjLdH7PoCT6ps9Tz67
zmlnf17jpgiDDEhLZan0ggxT+ERF6JCJMnlj4Jukh3VmT1BBfG9rQ14PVqrnpQ5GW1W4xbFL+KYy
1ToMnN1rYPJv4stWaW8ECbhY/CKWnLSE61g08i5KB/Hq+b21qB85cHSYoqLfUolAHobDic5QApXq
Yt0mZIL+eS5bKzwdaPPjBctYgs5bPPpeqzrfXarXjyF9BIGJs6+IEUQXNv7FL+wuLANnLOz4y0ga
pMiXEHv9ExQUBdjGU7MId09nn74AjBay/MB6+A/j8uTewYyC0IeZjQ0nyw9euI1sWNEwb+iGJurp
X8IuqgbVUJveJCMg/9zsbjvXynTtcE2U/uWZi4aFHNPN5YG1A/NxNGnv05uyRDlsV81s8e7zwRb0
KnfZ8M99rihmFCZjCKmP+vc0KXIZVCNXkoOvN5p4YXbPhHrFdAsGIYG8dNwcoj2fqec1OXa6AdvQ
unB7X6U4ihOfzxLdzLexFyC3z0Xg5klyjVT0sMYUmQ0XK2qXmj8gcBrYBuktFefjnSc2jd0/BeyI
dO0S1yDOYYCyZLardt77oCAxtQd3/ji+AwqWlW1JO+KqTyZ6NrQ1vugoDh4Jx/3i6z1mACrq9OqC
JrUgBytXkFF+VIa+iTx/axc6UMryjnErxV4CMj/DaUwvdSeLF5SizZj1a4+oV1DdrKu5ABFF8leh
QT/hhxxG3Z3LwkLtdXkslM2aVJ6Mtwayv1P7KHCwn1z4Sjooja8yNfSPPwZNGMzPhzU+T5ExZYSU
RjCkDGeOLzN5Y2c5CWQacc/REf7afPIM26rAj9rLDDuVZymAyjCnKBgzHNK9pkkanDFNNEgrjmmG
bUhPqmN/QaTKCub2zD9+ufuxnKhQKNVXN3sevutWQsj0kO3VobWYYGi1EWznzWw689v41TZngOXS
1dfkr80Al8jLUiQAmeXWPtSu4u2mOw7o3Or6/kslDBMQ7/G3un7bL891JyTewXC9cevwEqRhT7x4
DTAismXF0Rh+hcr6XDG7MCESwwA9YFjI8UXkZfwLmjjUHFzUGw5neSArUSlsuuvRyXv2C53sce2c
XJOGWfbM8SRkooSzj3w8vqszuineWstci+Ktb5x+3qf0S8lWPt5gYzSaEDqzFDtKoV99re/VTAYB
lfnjEzz31bv5eci23PSR5MTp4j5y8/q/OejAL8xQYdUJwjr+OlixLtVF8fe/v8k8Og8wVOtb4Thr
V8+oNqcDW0gv/pzGtS81+ravkhJqDn9+TsLRQFGTeQdD4Nlg+hol6eDd1LnoGWhLTU0Wr3z7jSZA
5Z5gNrbhB8GGWFjNUiAaHR+/83uVokENE4pIjL9JNOIAIeqQmGlVzUC9uwN6mtjRfsbBsXCprRVd
WdVzsfXDXQ4cWGwS9IqlYgZW1LeJ6teNEWXSN2m0St3bouQNtT6tA9TVQ+Fi+JWpzz04vwlAE3py
eHUEr9vBBXnPzFVsrhBdSOKGNxNQRM10f/yNpNslTrLYN9VWIIDqdAfFygj0OAfRIIM3TULD3um5
yfQBGLgO2zvxp87PdJ5SeeZNEihmtmKL2Q/H6FbH19ze/ouI7RjYcTWgRxmbO4nmGDii04E55ECK
YxDDkc8yy5s+to9J3Me020Yg4WkaK8H0I2nV0ZLyOfIL9+xAlBAnju92uEd1kkO9UamVe4i38tk+
/a8LfWpatGbDciMZetcERxH5WXZQ+IpByi7LsOsglUlsepnqsNme124os1L7KtoeRVwf2hhd/4p4
P5GKrHd0I7LSZOa0uyQRVegwF69OY9BT4k5V3MPrUeFjXIeYHvCa8AnzoflNMzBo+nwtwkBv8rmt
YX2bE74dw8Kv7gi1zfW+cJC28l8FlA1HLn7vVZ4JYdBYfvxl9UWOCyNVIjNTafWDXIe+EmyCnI+R
Yw1Y6QY0ppd1Zmg9XAnnTh1un8wzboecrVNMJaDzUE3MkagYCaC0hvSVvHva24QPUk3fhw5PFOhj
ZpBY1VZRuQLZsrEson8FLRU0LG6zh169wu50Vr+2nYdpgkssZ9n3kaunv/VMPcsooyS95mArBIca
cRHRN2hEXDhLn9nM+51AGjBltNjgtRKjjXofUrcuSx4YzpoF8zkNK2CVIunjjStTHSmsuzVBoVt7
PBi1IBaWtpVFoUEBuSGRiUjThluJ8RhmgB8NSRCJKvedUgLb8l3RWVRXZTlhdDVxFNOJPvJeLpwn
/RlRMz5mV7EcrexwkeuoPtgsl1KbamsaXp4WNtjMJwcUxnl/29MdLJ5Qtp1AGdjkiRO5LUr2FcKq
zChHjQPB2pIlX1ZYZYiEFI2m6NVUC+/MDhsJKL1pLWU6QkxpGTr4v1BNp6XGnm+vnngX5lwYuXF5
SbdWV6CX0fI55VKjtHlwPHVmzQ3U7gj0pQk6/VaB4EMrFIQROd/7D1xR/vAglH0pY5VTgBS3UmIo
qr2685rIq0t3st8SmijXDwlui3ePav9MRKigrgr/AsJGv++OLg0VX3VDNiGbA8qUmLmMqI1BgWf3
A/DqsdjG+ti071GIITxafmK3RcX9oEisEEbqO05RsvVHR5osmOCkQ8SbecUFsAVJDDdjRI7QBPz8
jZ1iatBI/7BU1DlimXhAJSShfGJJjbEoOuR738uKHDI8+hI2uEX08A+fBTnYGKS//yLT8HN7Aj/3
3gSuBnPRGEvprv6EckRTRlmmASP61KI5hwV4+aMQgTU2n5uwQ3xF+kTQIhkqAA+k31olEMqUMy3b
RNr7cl3w4376Uhvny9D0fZbUk6UJ/debCTohCK6F0nfBCeRxMRqcJbwu4MwROg18xPTc5asyRU0c
JwpOR+mr21Jv3Yi8ZnapzWSMnTilMzvkB+DicF3uKmRQbKn97Puex9XABkcFmPsmykDxSkPVVjWb
P4p6DsiuewOkEsrNtJRYwYZlNvykjRZ8SeKR5H6l+TUf5bKGhAQ8Ju6hdFSbist/B8pcXgXu/s7r
3/rdYtalrbzEpjCXf2ANav8nxM8ITnRuzeQsLuQCAOy1aifU7hCNNXyrjd4XRIvVEuloiq4R5QJL
aAyenxSCuSBteWBE+xzS4PKPgazf9dB4c7bbuPe2+0xeBkZkZD2a9Bbj951yiZ7/UVci01RfuLho
0O6d0cwB9RaUPdAKILYFRe59SRGbItspGL5PSntOcIqZ/XCcPKGzb9Bni6YGnPgkAb+2qWk/tob3
jQ3e9gtLskUkowKHyvVeWh9WQtjnN44OuGzWHSVMviAzXdFTaAGc0kXmGUqFJ3y2w57e9Ha8ExKa
eGfTFolHf1TfAhJyJJ68zIpEgPQi5D9F68rGQgWn2KtXFp37ZytPjEIq3V/mnW1TolQVb7KBP196
ON9tWCh9Qwscrc+G5X5u+/DU0gX+58675ah5bAU5JuuIuKlxWWzHnaxkIYGWBhrGFmMFZGXUg54y
NLbHIb4JxFlvelqBDR3ZW4wsRkuC0TBATwK2egnuQ9OUcMGua3TMKGjyz2mruHhF+OSK1cUxU0+x
yrtXsMmWe+R4j9Ubwo0lQO6UwzU1LoxzBcVMjoHMWFhVhmbHSffBfgWCFHX+OaDXtrcKO67Y5v6/
T6AUtW4/dTxcEw+/BqGC3ur6mbcnbOf0sRTB8dzIqqPckB7IuPJSDDL+16iZ8tLwp35Yp0EkDZGc
pPmlFITcb2DJzHcp5QnxMCU7ahXAJgQY6nrLroDiy8s3mJex5X70EXp2zaP/EUtRr6pFNDPgTcY5
60sgyjMcw5e1lv+bVUJWvdMIGxVxwXvT2AJgfg+SqN+NzKBsGsIgSntXfzA5SPXbzO8ed6Q3dcVY
DPiWe9ajxiUig0Ai1wD1EM1tHqOMjzJcsbmv1Y0drYHPghYLo0U8zM7PB6+PKH/gROs6atSf59AP
1gX0wH4jVPPZJ9neMeDcfB75B8pwwPUapMJj2X3ZOdbB8Th6q9JB4ZviI1M0gsFMJAXVmwJB+t5X
+tpqnAsSrHD4bHRI3W1SExB466eTILqAwyFF/rrvO0biZ+3E10sCbN/Y31VDJm+vKNbBsowPtatb
/LYWJRaSp1KJYA1xlcpNs44iXObge8JkCkR2j1r3E6JStq97StV93JqnK58NaeV/+UNLWXv3uCWt
FwDphl0jTr6LmNl9gk0Ujpmf+S399nn9mhNW8AuxS+gLUe2hxtE0IFKGy2GcNpIVpYRQYXkkeAQO
zcq2LFVQ43yuwo2j96lQbr6WtRfVmceK+eSAtZ+zWQMmePeNOq//Z2L8IMqUtEChoj7pJrjOwCxB
I17nYrEHTGxicZNKVhB2Rze/EG0jAX6N4iB8E/lxJpt86fG8u7BsQhemG8KELBvMot3i4rzhiCxq
PAbMlQqUUqifA4ZR2usWuz1quzrmGq3STMfVt7x8IK4sOzLDuxfckHtXM5E25Xs/9Q/zP2t8W2PH
uIm1QJL9QGo9YPMHVJKbHp1TX2TBdRfs0oPWYolq9WdWPpNdAV7fVsi4YrSl30QRVWh6yvcPMGyP
jAVGCpb0q6JkOHOXjUrlWXuY8oxMLOXkHbicrSnAFZ8YxqY4Kx18MfKSbVmzX6y+FmF1MXuaAAYZ
9F5XjKWR3ncLOg7Zf4LSwUQfg9qjEt31P5iKsHHs+7dFahN5j4EVjv+5ZzldAMkSj9vzY5yJhPi1
/mdo/pxp9jpKNbecz5yPFLe3W4WuB4s6GhNorF4jcEkWk8I3GnpZw2Xb+lFTdYV2slVoFbhfyIoL
8JZ9AXxkbp6iptf5jiE5NIPkA6ZLASBHeoF+msKkC2RKuX8N5of40YRAXFJJHNlY0BpJh9WC7cW3
dNlwDFjZye5oq12QP/T+lgCdFRF5vAo8gT84VG8k9DXH7lBjxNC9D5hg2T+vMd7oXICPEFjqy0Gv
lwj5n6t80mE6v/Ebxd4VMiEZvUfxdXW8AT1NT49A3S+XmJuaVAcfxl17c4m5xsEWyY3yUb/+F8fK
/MWTfcSPNsMf22Ni7C+mFZbmMhBh5LglTO2YxYCx6aLZIwhqfsx54l2jHeRMbN+/9Ia6DGfOUCPo
nqA0Gc/Mh1/hW8zLrgsycEjWFO+2bgVWySNcNPeH4fnp/FFNbwtf1gyrg1Ccwt8n9GwaCO7Agagt
j4RPOMR26j+MzaXly920EPu44OxehNjskhi6nl3IeUp6XlETv/K0ZkZOA/OXyjsHeZZc+k5Hz58I
vVb5JStYhvLkTwOLsxsnqMxxc9xYwvySVumfLKWXyGbPjrBdb0dYQJCk8DwhmG748SRlq7vQNtzB
qoZFXsdcJb3Y2mA4nNt3IlNXqc1ahFcSWof3q1Xl/pX9xL2GE7BX5P/17SEewABNkx6O7ZAQH+H9
npDDTftKFaH9AdmJV2V88MrPQZLJ5ILoHl9XWNTHpJnNZLuETtb2PqUN/15nelPEql8/sk9zQsw3
0CuMFme8ZqvHHIgTX/nJ56e7gOVcXP4dFBf57FITHIymu9fdTXMVlqRED4mid3zdsopBvHYapOFL
GEhGE53Igx5T1DRHCxGYSoKMaZP+Uyr7i/ExxANq41AErYKWWdgfyuRts6ibESFqiqR/NalhT/jn
J51fEst6AEcPwSLXqTrWmR9xqmlx+BhQlJrV4Adj8D/51GhGVo1ihfTL/XTkCJPWhdvCvjt7rBvU
ybZjdPXMMhaMWOmGr9V+wugX/jG9XfuJ0qTH8Ty92UvSWDOHxkcNon4bqNBQi69AkyEwyc8k2wP6
SxFftyqBCzOV54HxRev1lFrJ2DJd3P5MidB4BmB6o3wG8OQpPikEsKpHruFQNUgApeULvcQNLkhj
ozB7SJ7qGITXF1LpSJ7336yRvuAlFY8NHDGWLNC7/z7B3S/VFyPV/6AoTZI82Gi44ibL2VWjCSU4
gIVA7X3853BiKUZv25SBUeLIyuz92AZD3xi7OKxNX2gh3XHdtoYunwKDA8V6fAh7A9vO+2DriXvH
OzsmnxTOvSaJwqwRR7m4CUFbiL1qAp5KVzGlqr+hS6lJ2JucO/5u8UXQupOG6SDs28N+JUe71RmV
UGPDB7BQ3hHZJ59KUNd7fdyWsb++0QuCEczjcstnU9yA+uGyjnPkpAJ+1GiCCcelDT5n1QcTEOp1
aaPvKGssZvwluA43nIgR+/P/5vcZWUsBGJBq36o856nS63aaGOWpbgPNRIvQT1csU41OPWMaR2fm
GibJBI3D3tathS5sOMuu7DZoaiG2M8KoXbnAQN7bo1u3OXzlcXP2wHE8W1fA3HDxVKhP42UELpSw
gzh5vIQ6/KNZsjEabQdGjzvmAQfjdLuxkoU8WJ46u67veGAAkQwYHzKxt10HgxWnYAaAo2WANQ1h
io3Arz9IAIlBk9jlxKhuB8Cj43SRjnEmWn0u6S4i/BjJAEfNUweBiKHMwHc4j9jNuBeWYsLlmOZW
ohyFKP/f10E82vU6UIhJ62IqpTYJ84HrZ1pgG9BLtGgCCVzdoGafLJD9vmtc2GGfEKV4PV4Azbu7
jcuCe3of/3sWX3Y7b0OhPnA2zTWZtWyvWiQ4k5Tt6fqSEE/VLrPLWezF1HI7hcpNpea8QYtv3A6d
7YYr4xHfUnpF52VfG4zOyIcZDZPbV9u+URlYuSl+Wo0ulZEepD+d1yvQMCK2LOPRTOFBqPMzLe0p
Iy3YlMrtqmVNB3yUVvX8fthlJHLVw/Ck0/g/0S12gidRL9CGvyq02YU/T1vuFxoPgiHzmQmTqcVL
ASgMp59yEuVqNZA2WudbANGMPv1k4gEBsNgTkWaRaMWaby8nscWKXENaUTxXqiqAu5xvQ15rGay7
1tFmem053kFcDbiCXaxhLcbXm3zFIrXUV851f0mbSbQFEcHDej8y0hQhwzOtR5ujEcDcizsB8z6P
ERd1WEszvG97PpzAbqLt/Ksgw8xKKD9cUbmwlNMEPSvm96KM9XUjdcv6Dv8vqjgozONK9ulzrz7v
UUShE0ZCs5+Lb7g3bA38nIf6w3JDdJnF3sODmjXE+RUV0IJedpwcwUDXfjPXwN0++BM085VvLQX6
gJG1+3KMtFrpwKbn+QiB+FB66Dye9QQAZTMMHNM5j7DyanMeIXYddKh3MUy2BbFoDH2cV/cBiL9v
tgfqLwQpuKo2dBbN7Mndz9ezp9B64mb9VaAEGRN9jKwKTth5vtGvm7micelAnMkThFVDvK6qE2Ip
gbg312+/VR/VBzPuopJ3ZoHI0SFllyJNrbOjRX8l8Nbc8yud7HVQE3Dz+HZLYGU8C7x53CtiILhd
FQcLQcEzId5Ir2X7piHdHyIYh5Qww8mLvByBSBbAL2bBM2RQ7sp44jj8QO1mfYIFRFcnZwCsryCd
uWuFtuS2WNyZzCpJ6rbR6Xm2XbFm/7gBkoThbhRbjWQcImNCbW0L8GCQ9KiTrp6OlLTsKchlj9eh
wJu6eGXSm7NUKKrWyS2/vbvgfCssciWOxxDUflw0TTUV3hrRHTfZyvau0V46ziSpA5Nc9SkhiYLS
Wkn4YxvNJ2pf5lWCO+qZMdmpKcBUsWAv7JAuqpnGeoV4YdOW1Jes8ZTyEs+MKV6RU4moJTl6EteH
p/MCIY4gxJRXQHoO8+J9Y91qkx956HNOBn/QkaBeIkAwqpAb0iQpXzHWd/fRqdahqj39SXtjt/mH
wk7e3qyMhG5IUNLAOPTuTUOF+/SNSz+gpxfpcuFpj9+furht8JkqVzD7JHGSYbzM2fC9mmU/ShYF
Z5krywfQVujzTRhtARU05e6Tp5yLLB0WNzEJjNXKhsBrdx2SqnpYa0uERBOprgexZVSRjjsW+jpl
x649/tHA83ZJC4pzT/+yrwJLztO0leqcxhmEhkKsQmQ7PY3e4kI38qTmtvdTjKQwP58937gc/Aqh
NM3Jr+xkaH3jGr99RWvwJqd0FJJQ/f+yv2Li11OWVvQGO+pysc51Z3GFvH13JuR9HM9/NqIA5rkg
Kc3uBdstMAcRAGBA1Z4C5PTCW65urTiuK1LX1ogjZioWJhq0/H8VwdAfYls4s+uuQ4liA1zRy6U+
g7i/Rh7FoLWRhut82/rt2NQSTHD44WGkjL1gOIxm6zi9Z/n3OsBjAMl/GFjk/4j/yZIZleqHQQy3
OGxOVfwCTw5uk53+n7gnYeJ590ijqC+qhb8gkf74+ZSm/q2CLd9f+UJ0TlKhJ6sWQyqAZT8qy3G/
bcB2Da65IHrEl2RS/cY/ZwaiPi6iIOADTwCjbGo0SnIHNzGv/6dF8UEDrVrPX7GQXTr7G+veE8ZE
LsC+q3Xvm9L99NozDwVie5WrUMiunT+zKLZrSmg1rwktw/VypWqAIS9gg5Vyy0NCNrhvfQAF3u9v
rDYNt6zjqOGaJpny28TF6zylM9BPGDLNPfD3jsEAtIf22SnHyAnpmi/OSANkKk3KfSi47HpH2yvn
oUwMLr3zL7hSeRixpAlNJTvILx3gPx1u9Zcxyf82Eb11nuEZcDFu0rBGZGpN7Wfdh0qgG4CA72nZ
kMIwCSC1QvALGnKT/NVSviSs/deQiJq3S7BmgbBvrVKTLmB5LwpRnK2H+RydZS8WDkMNeRvWehQa
qeDt18SUIlDmc9AeAJ2tC+tL7K9rGtVvii/sJ/EYqXWcaiEesc2QsGRScdA9nSR9zH+ipBRea4me
zT4P5po3yeVYkjcDwnSwgKVjc87aBFBLf+ItWMcqBNVj0SVTZ701U8U6kaxSmgx9foJlWZlAPRtX
GhK0OXkLwI4X9NLJvbO7hDwZajhY2e3FAe5Mg2t6LXkg5FuFZPpfTB11ya/WK/jXNzq2VecIgIyd
E+z7S40y9GvXzKW4+WRcql4e4SW9HAX1nS++dqLrS5cu6E7blq2oCdTeytbR0KQIyHy3yRMvhgTM
2MCyzRwGDlvAfIJAzV8bprdQ9Q0G8b/Jr6ff3oTrbYCz4JWGexJ2WWsEKGMdZg2XNBHv8rMCGFFp
XI1jf0UaeiBcd+4ormpL/fLhjnftDIyCvcMQEWJg7o3qrMTyoEuCoZWuA9/BEXwVvKIvxQwdYa99
kca8dZKNCv+322rJSFRWgqDx2SF9IHQcFGCpMKXog3Vds7opJwhUkLd6ZMrYFM1Z7TIoQU4+y93l
AOuFN13QQewWSnhhcGk4SEIa8UmOWuHJ2vX/3ZUAe97pipw1c2rRPn4vfgQR94ZmA3ltn1adp2jp
x9vM8HGwF4djH0piyk75Gz5dYbBU07njWnl8Zvhr8bGzMr3EsuqoFgQZJ0NW+fgutDHqRvPV5lnh
zr4RSirOt1FdSGaJsbMCfgBZCU2oLGxeyDPJZR0pIx4dyJN2vMyR7ljRoEkiGrRpaFdftD5yM+3u
7yDb5aqNx045dmNzsQduAnctW0P0FlVcAlSUIKP2vGQ1PoRICgBu1FSCJjbOeVpY0NZkCC7KUHMy
wLRMa/zbiEoSShf8u+btSN4eg7f0Z05QHgwTi8EOtBg3Y75wkLqRIOIW0WW0mCdBMf6bCAV0o4fs
MAd0c+5pQiVZiHYLqJHOuyuu9pYwXz61mbCn9ztR8dNrB3IMKqOUi7l2+BVF4OEfTVlQVpNi8sSI
FM6MOa9bQY5ZLFEpLUNtm1cFE5CH9Llf8xGZWJmm7r+hW/WyV7tx3Jt/0thjcJR/zMEloa9v6oY/
K0/YBMoomYfz6lj5NBW5vZYFMHNZp+4qY5kO96OQV0UsuM78oIixjUSsGB7vuC3M4c2g9Y+TEzqE
S85SlaBe2Z9aPqBcZRskIyLqkNNlwfAFWd/niXw3EyVgJWVF5rb1U5uTgwrBZAUNaEiSgX7FY4Vp
0Q2v2vZi1YWeP2Gt5lfHXciI4QkRrq3pFHziQ8BVZpPjNP7/0cCYLcBuDBatV8LAK7dk5nwU/2wN
vPzOK5LmrvW+lMwxlIUhqJXuyXpkzvouQn8spZNIuXcXtQm0eIF0Q1W0r0qbK8zNZbCG+2acB9jm
OjfG51er0bx1cN4Ru90UWqWC6WOHXpES55ZCpzbHj113wmqcxHbaYIAJeG8VtIl/jQjWvGXjD3UO
tIy9BIRDstNrp6r4zUlZcJToKNOUDduTTZDIoC3+iq52tFfOfExTk25x01CXQpWv7YLztTDet9NX
enX4tD/fbW3JFbm0vMiBcHM7ftVu1Vkq0xkT4hp4Z2eX2SZRdhvdHE977j3EsnBs3+y/4xAheLGq
gSPgBSA05Ed+wUd4e3IvfRMIrYhcC8Ylv8xAVLVmy6GhKEtapE6pxY6UfTGrVOwhHIBgHq18mkvo
emRcQ3BbsQoo9IheJWeRpNeO8++KnOHxJVvG3sPw+bQN+x9TBY1WMFq5nSFfqkp9PfvVgJBHS0xg
nzhKa798FCsxSND68Bu+SWrRi7G5y+/Wtig7b/+lS33o0vbntyi0eBqd0zrDePHu8epqahLYWsF/
he56sWxdfg9MWEPHTcLjRvtkriuD+l5LSeoxQpJ8XYq2nBON+ynfoYac8uka3HZkAOz32nqHdtRk
GVRe7SZct/yQiJI6TNnL9yc+FXzsoI4rfQsvLyJo1ZK2/nFM1AZJCxpLQ1+tZ9DP12NYhQ8sa+Qn
xnZDTFrJrRQORpzKpplDn3Ynvy7PKj6IDHdtJ5sgCxJt6ZvwHNHvUozZcNn0/tuXOEHvYJSvxCI0
74DzrNw+cEJoEf7G77njgxPpBAVlk3kRnPk8lVwSKy7oGMlquz8OxQgJwuk86j0fD1oCa3PVWES4
dnUCRI/RD/mQS7NNxE9T/4X4vIAhyIsUfKdP05MWab5AwaMMOlNLquSLhQOhOoPmlfYZ64yJ9oyg
DiN2LvzB7Y2o2AkeH++Hm8UNtLMseO1fllsDfBoVZSEoER5wdCvRFf+PKCoNppb/7ISG7hiBgdBD
oGZoyayw2oq8GQg6LIlqC0s5CyRBNLh/15zr4a/EohWc4pQtcryw4Ni0Dp3wTXgaMXaAIhxE8oK5
os1DXIt52rSyhLOu1UaOdhH3R7u7yrQdHR33Cg5/I06GdG2KKZN6RuPhfwj4bFO/LFWuGxPkca7+
Y1bGxIA2skbd62btgtq27+hIXgbJl0CmVAwB3muFBILfyoNiZpAJwMvRN866gXZS28ApzUuweBNE
XBh3H5ZPEUpJ8EI4pro93tQtKPRHWslA5zM86mXihF0mfIVpRGchq+ysqyZ8xQCRyHZUT28jmPA7
dB2wMEIdkyiNuViG9fzVXNSYe6Yn97gPk5vPtOxSVhnUnoVZ6ukpXzU9H2nDSpp5lvm0G2zU04y5
rG6P5OhaFZ8Klplv9B/jqOBR3AhYlGwdK3P4iGBXNZqQDHWOdPnbuKTAIOpgBHijE9tZBej/vtiO
GZVjvnZNhu70NbdDCC9fSgVY7RvisReW8wvn5EuviX3ksjq6MAX3VllBnIQbw7SZmjCyE9959X5c
BzGM2rCnBPZAwaDdgY538VPWkPSSM95pzjq+kes4y2K2gQp6dNPCuI75qmtO+LMJNb+Pm2zfzWhN
d0A/vuQYwwj7AgqSfFSr/TO6869ia/CohQ9fpc0bPjG0njIotq2EdLCxI0eXc1LTMQXhZBYFjPgO
+wOvce2zecmkq8woS5oKoU3AiwWtipfjIOGVeB8eV19jbhf/ObFP6KabDsHW+TH8+1UAIatZ4UsW
Xmvqu64lRi+rh8wt5nEv+XlU1W9ZsETRT21oCWdtyLcQtu7R9yFgy4/nzkGuAV8lN6OkrFBe+WWL
4escieccLZUL+BtRnzWbF7Ftlfok46kJAsoMB4kOR9PO3yksNhFbuoPe4Se/AI8T0SMFyizUnaIK
24UNQ0l7cYIlw6BBdCKQQGBju6VVBTPSyk5N8oKKlbIeegH7DpQxI6g9P4ULnxEab9YNeFLk2XyU
t6jUi6QZP06xkeWWlhEa5oo3nAryg+3i90xEi9uJAyha2FWLkUPz5eg7CPkksmIgmJLJ7ma8fV6g
NKOiPCyDN1TzV5S2xhWYPBwVtvs/3qFOuvWcmRNs9q58KE2Xk5aUChfRzJgjDuQyDhYO8whWg/VN
45KObLeRbFmOi0mBvKrSG5FeKrl/MoHVhe6NpIKPc7aPz7sCP9iD5k6VWLgRrDva69jb2w5Sm86N
n2iPWyvMfAPik2tWsuMP7icOjMDo00ynHY2qXTP2rnuG7vKTOJ8NbUz8v6CX52Em27XxpUX+dJcN
1Nw8/fBiXLF/IyxbOtlCvW4ULfADsNn8SVetsj0bZ8AuYyMNnLPYr1aRfaVFGxHi6V5+Liyvnavm
DlGK0gRSPKe+FCtZojBAPgEd5VwNHvucfmijv9J0ylbaEhVFHpR7armjCuWH8eq1beIidw0Rj/tT
1tV4p+iySWMCngKtDLtPfhuip3MzjA8hM1l169d2AEnbBEkljTtRdYh50dW35HGjdEwefc9xijnf
Zg7YH8pa05Z4AEi94k0jWVL8+DvC2+a6Tv/et8j9h3XF5iUblu1AJC3mbYHGuE3tRzooRbRrSiSg
1M8g/H0V42SDORnwoVAgk3KV5pU7f90Ma6oBZNq65jVvK/VeuE3wmQiIssEYdHqFrpnfsMLlb7gH
MRnNSOCxORA/7JztWL8O6PszrwfXCfNkGzSz0rkqpCvyLNaPH9u0yXApgUHkGrGQOM2L3AAw+plj
PJihB+0t9u5cTApLZ5ITMnUKW95juEdcKQNEGzG8MJmku9aS3nyxjmjzmQikUwbLrSV/LA1Dtin+
fehRQHAshJY6RVUWe6YbZPjCTcZ+8ddDfx/wrXJPnQhL/QrQCc0nnfCayGFV2MUMuA+Vbv9Wgfd1
Yr9ijSxA4J7lqC76q4a3ZeFh5eIxLPgvoZ4Y+odjRFX6NnWDT6M11UqHYBOBb4QxGj4yejjI9Adm
7OMq8vclDuDcwjIH0sRb06zyAfKqXwvvpP2KYshOyci0eRgIxL9E1zMOynnLxhN63pT5T5lFF33L
pRNRqr9FCr2Kf6e5coDILTCKIZGhyoDXbe7UP37eS+vH00JAQbsF8BAgXA1INq7Dv6/eueWAcLsl
xv/Pcdeg3xbFFJBL3DqWtoIy2pOTyVchZac705SBNOzzBy3of+YzAQBpZ0uuDNU9jdc9k/JLN0t9
4Zjil++bb6X9I+oR1y64PIzFEOln3NT5i6OpiWm6sly1waJxQhyb61LJ4/A23Vb8/T3SqGyVw4gM
EB00cp6fb9jxvTtAjdI7bmSrOHpD33xHXb6QeBh/VgoYSwN8u+6+qDylQc3o2IaM8z1PENMZLfjW
JnugN6fasK1ONB67ihkofrHPXmxoI4qgANCySOjZQow44JrMbtdYS1Rv35K4rvDvC7nMl5P842b4
K/te2gvkdHBnLUsmxqsXOg7lOS0Zcd/A+Pa61Ykq6ZUL2EWgvjEfUA848CDbN8Z2iqajjkDR+u7Y
PCouTvUEUe25FAvcVmSxG0RoZN5B/nw/UcN5ehpIHRwOra2kmXxOwtwAVB57ycYabu08vLP+aphT
GDhXuyhCJrHrn+u1Y6I3il0tSFLTEBdK/hI6maHJHEsbFBapNeKtkqZF2yjgHvzuGOartR/A/0Bj
q5jcYZ2MzbevsYOGCIeMjYyH0E96opMC8C7ZhTroeLCM8PxasxjbShGmlhE8Rr5hnckkFQkF8gQs
cwt1T+l+Du1Y6NE3OP0wuxErtcu7mb0voQlCikIZ/W7AC5hCVihl1fANEv+DZxbzYeI/oFzXhedJ
2PSQ6gkMVD4fo2xl2L+3d/tSv2kkCIzE0S/Myd6gwgbJRq+PB5DDEs+1t/nI5MkYYjhhoBvGDg1B
QYrO7mPLzMor7IocqXZQaIDYS3OLnW6ASUQi6LmiZZjifVATz/BguO/A3TlcbOEBevWUMSLkSENY
2LBKPlYps8XxNUvt0cmMmSGtKVEKEg8kb+768IuNibggyiMU3k1Zf3MfkCK2rA9W5+wfZEDuOdDD
VNm5x+MtWKDSPrBFOGYxCsVERfWGwAZbRX2HOAqt3pSf7ptf0lnmD48bwEl9pVvYI0bmhIbqOz2Z
jW+HpD1KGihA5fbuZpmo3/DZeCI4SVS65dSodxP1/moT0AXyh33AlEH6DKVJXc4owO1KrBmr7BIn
ZAxJpJzuHAgRfth41PmtBlSgdCCGFn3Z9o7QOy/p+SZpo+kCuxAhVzL2lhb5TQ1gt3DBxbb18vb9
AkW5s5Bk3LtuplFpyHnX3bpHEcCsFrc7497HnUkPlUt1hhFQhz3iYFrI6oB2z+1lrfuTTyjYbb+7
J5dRe7MK3HMLlTgxa6aWEGaNsSp4b8BA4xGe38Lub9Bx2MjL+p4nIL4rKyrVtw5TVaSu7JQUjQ9j
q9PF3+TOMJI3sjY7sdi2RN5tm90urSOaQb24yAPf9xPBE5RasA6b7Ml56SadagqoiUK4tuknbb+H
bL6XWPIIipuzzn/xJUN185n65Q/pNIWx/UbhOCR4ljb7RMvjNNJsI++4D3wM+czfXm4J//D2DSoB
n+Ln6bICUmQE8oVSYfS4+EDr+GWajxcchWucUXdvmQnvn6yPBoj2mvUfbH01TEYPwVuGiJ4sB48c
5aLKRiYeANy97gsTolxopLIBaUiFR/q3tHWPCeynoV/ee5CNyDMmLkLP4cBdjnSpAHZ/XT/6nnSE
LaU6NYlkHwHkIbOk1S3gfxgfjhVyijHL9JPqD3gLJjvYNNRZLSNLsX6rVH70rp44UE6Y8KK4c2C+
Cn4ZRm1oqm/ZG4/Q1RABGDAbMJakY98qC0cU2OWLpLJc75rAdJ3KS1V/k2614+77OttbFpXdEvfT
Ux2omPNWWRaiAcxc/vGDx4Q0ibjUqmTBdtqJsrYPtGEdjIIjAgVwxCoC2GIig9/BcZ1xAuiNtm1/
CcPDhchkDnlePnqHU13MjR8aQgMJZtTCCLqNIQXqUi1ElznwrRWZAuveu3Ade7XWAH48PaYrgBIr
U/VAJpmoYYYy8B0KxU2mcCdevoZBC+mz14KHabpO6LrJJTy0mqAa9FGztbRWgAcm1B9vHQpGf3d4
0f1E3srABdoPpaiBmGQGUgnT82s38WuClQEikxfpkx13TBZAWijscFAa+yhaxZrn3QpZN4VJVvRb
/k+9YpFJCkFRUeRbsddRiTPUYWNGObRwn+uy1xzDsdw0dlXVcY9t4sKd+3B3Js/aJc4iSjz2Ol60
oazk+54Kn8g0A33DKMhYLAVxpIp3ClatN0PkWZLihHdn4klS3eySSDnuhUI1TTiLlBADs8N/Xkqk
Q24itLG05EKfccQLH4zKgDA3ollijC27qwexkMtyTN6YZNDbHkUybgUOQLx3qbTxShfpotN8CLoB
OPnkzWQZ4tkzJFh+zrk/njp0TfKOgpW+6bcOkTmpOnGdiERwpafHT1lqZICpvNst8GNw4rKpastj
5HLafJOe132YXbe8Hg+71UiSZ0JPs3mygQD14Ot1xmEtvVY7QUg6bmZgLv/C1KV1M4UaJotIY+zr
rvGBTc2H2CQgp8UTvavFZHi8cdkdb0gO0ERBTMt77K/wpEr2X14jMYC8NlKJyjTBuPsdo/qBAhjd
HblnrPunLVFlnT+9NMeQ22PPOdpnNlxV5vTQo3hgJm/GqpFzNynaSxo1a7BpgP93wGiecwOafeQN
cngZZEtq8wgh1G9ANn+8wOTnIj77W6XbzOl/lqHWjfwuQo7jz6WR2qWILawXy6z6TCADWjCooeHI
ZYqUA8Qbtn2tnexZfeeo6re8N2KP1v3yvFS0EBYHDigPdX+dQu0RJvICUW+JTDugsp1VwbZruQ1r
f2ksmHkiMxaQVolHh+q/yKPyRUD/6WD4XY/y4l1vZU3dmnxaUbRgVUfPRzYrLRiDRdpWLmZFNoSE
zRCzb7BMXKYs/snCBNsPnTUCwU5ejJm0UVci3EczJxx9QUC8JVrm/3iU3SRORt2UDwmPY9cDTF+T
s4vdVhcnS8tux7FlnVRPXeOHNMibPXuw/2NU2vYIGjBIIj225RyPOofqkwbWKxt4qz8YlfGuZ5Mr
Mkb3Qt+ou9T22xgh4LmNNLHNakQ+eRD053gIHIZ4vRjovsCXge5Fb6dJfq3D505HRWx/TpvanAee
tbeB4NkniG5KTYtmYx1eXzs0u6wQmCCPSNzOq8y0LZkev5/y3wkJlhj8Rmw8F8+flVT1gv1Rqj5n
tQqD5v72vOt2zzhy5+UZkInEbTQ4DbCm2hIy8vK4trx21/G1XiCR0vmkWOLqnhGXx6PUsOu0qqID
+O4KFsueyROAKx8/OJM8SEkYy6FDo8MNYAPQ7K9R+ACu+XnjDlP8fwls+f6yunaUoOd6ogc4B8WC
CllWwndb95zLfMB8Qqk67IgVWWrlapWmYxb28VRHdT26UUAbKtJrncDe4LwMiaj+heYRmWufK+is
6JaXm4SsMF09o+1XEOGeXTQAcC+6M8xhgDTk5hOY5EuyutfaRrfMMK64EseqM0TOqACcMuRW8rqs
UFCEyvw+45ZF6Yumth7YfMmZRktpASieePYgFMv0wmxF0x7rhrw8EWQvzJ2pWfuzrhK8s80le2Bg
jpWBZ3HMuHbPDQJKY3blKYj8KHKIj5sHKsDfOzCWnCXXfhNBhLqqufkDGniN7RKoBnUszTu75NAD
Imt7GCdsx2FqdYP4WqokYUGIQUj8yD6llFX8hsAAgQhh2jq4zHwaVi0NbaGiyq2MVPzPuWhHmnHo
KyQKR5JeFPAj8hnpOMozmBcQp/UTgAJ7JwF5Rl+V8tUToasm5o72hJ+jxjseJNKAOZTpo8Fm0oOf
YTY74vlqmvxd06GKJyMTSZvgwaMqyMH82I2347p/vATGlZLb/VFcJXk9zR0lR0PEErVG5zWl4QpO
peXBqFiHXAj6ud/GrSwS/EwD5Lg6zwWud/GDARXM4/40YYQn55KJcEafvbByaf3ZPPniZdTVvKb5
y6kEpx6bg6NM1Ec5GEToJQhDFYdViyA+Y66WqFZe88mlFlZc4zjOP6adtD2s+UOrfapqnbFvrFFI
zwsYaWtvI3Ii/A8WoaJepYLpy6ZqYs7wxepgHgJny+gA3Teuov+qNN21fmxvQ37RrTL02OEzcliQ
jEOVSrg0PxurxUCpRNntG8apX2Bi2bydjwyJ+lc5DE3gOKXDWK6ZyEnJCG3M0ZFWmjmu7o+DEdoW
hhiAX5ME4czULmNlxg+ckNp6Zb7BNRugPMZZVscLqwmu3b/kclZQS2wCq83UOia9hofohq+6wZZU
kHI0uJn6Q6AHxv+LW8L3hI9FA87AapIGlXrEmnTma9RWvQ1qA7yzAfYK+ESxJTBn0jdeed+5wCDo
CaDsAdpHA88hjcIfZY8X7M151986xIfr9K/15BKL4775MIfNa4PLvqtsE24foqmFvSxlcZMllO+n
znkcTHrOXx0a0zBph9VA1ksJOM3P6ZOw355E3GvXNWeKoV+BGu9Vw7M95LXhpQ4DI5OCpV/0IiUg
i3F+Qxfer6RF4ZTUWEUe3ABcGBVjt24580o6ef4pw5c6kEd+xJ5nAp9knR7GFJZhM1NDlzqfP3vO
ABkyYu9809JOELLCJbzu3rgae0QNCk9oRwAaoEepegmcZ0JXGwaTjr93BnFonJFTGdoxl+2eyxDY
DkLuOwr01Z3hZSUnpDP51b8jjTuWZNgqOEMiNx+HsEuWv41C2mpr1LH5R08T6mG7c7np3Wh/ad+g
t6vodXas9rVQtvl6nFPyZDIDscs533i1n8EbhBO/HbPmJnoaG1Egk/JEZG+p2nbBdYZsGU9b7Aqg
Ju0uwDMDdYLy9ak2FYVNL1yWUyYB222Tp0N8gPG2Ei48FFiuIrz4FCMeVbqgvw6w1Hrmy0y/2FQ/
sm2U38D3MOeh4uiefSxkv1+2A6sFyKeLYOi8JtxzggizpjOwkCq59BKbKxiBvSRhSC3aosXg2JF4
+Wp5bvpGdrCCPdBd9h9OarkLt4ADoIvENtheJUMtc8fwaaY3R6AitT6Wx1/duv0S/+VWnAFLQXdU
7iTcnB0oO7YS5EY9BjIen0cNvuVRJrOGQiG8SVM8//pFAjuVUyk7WJzjGE8mM8lJ7gZpxm30esah
8CWHamSxDvr+l/kRNbNaCz4oGYB/gAt2/sBr4WSLc1D6vys5U7Q0II4nxARCJ6jUwmWSj68fmKvI
CfKbztsIAJ5cIcUbxLw7VOAPwJoSxXvfSu3eugPyzJ3d8ZJHpHSvN0YkJkWbwPckdKdjRTIAyt54
iIWsOg4iQ2SsHt/ZB9rDPOoF5KmLeA+BTDzJqDTpcv0pkBbTWLJsVi5yX0fqEH1NoGMsptvnGJ6Z
T9hYqn/qgzn2Y8ldSTtbD80LSDbWDyR1gbgLqcXFFCRh5wuQP+W5m6tOzGF+XbpUpJg6Bycf6zyg
DuhG2SKNzOWHUrFyvamLaOduQXMtYklaWTsMFMYPKmSlMfv/v5QC8Md/CWq03UJxgR8smIcn7XcK
ttiWND0m1ypJb5zHKPgTh5xbg8i3h+9XPlriZJrQqmrpKdedvusBe+q0l5+N10crmywB/+xGPFCB
CiG1R6MpRBpBlu0+ZnTA7Loii7ra8qAWWtnZxTkfPX9B2/NaLaRadr5bUmMt03lqXzxR22bBZCEJ
GBjdQlZuSp/y22ElGeTzCHdi/BdlFOSNqyDYYPlTYtZMFIVtIleMNyj9mb4zdOA5uqgdmLEANoJm
r18uWr9XbmkQ2UP2sgdxSc27qvbhobaYZHJaifUuZ26dPVfGVu9xrOQPlFv2BHSHn2OxmZpu86vi
weoOfwVub3kzoXkkh8aqzD2yYnZEWI7oxoKbw+CfYWeOzgqWUPaOa5xND/rdpMjHQkWJyncK8XYW
jzGPSK5xljfTfqDI8knbSyVWx7QkoGlTeqr+R+89kN4ZyAM3CkgbkX8PUJd3icbieCHvvpsVrSAl
rBYTIJ8qdODiIdaFEvdEZVxErqbnBlUjhVXHIgAjOECAlVkkl2XqLQGBCD4awfe8kr72iSR6FgN/
BYfPADGoFN8S5QsP4IuSz93R7MBwgbWsZQyF+2Uvep1xa7cc99VEhgMTCKmcOWgHf8PxN9dxwPWx
7qmaigk/XKcdrANZimqOZdldjw56nfW1NODZQe1j+OKso2OzjY3ETYxM8V+LmBWMwPXqoZ7LDbvC
CPYM7puA+xR2uL+4ysdQ93VZ07STE72mGqklW6CC8oz7diKiioZI7K385i3Gx7mJ3d7H6lhExnXG
l0bZ4d4eg/b2+V5vgF14I10hRGWXgUfvv0EJAzLBRg2CYHp9IhuOwwaBtILXQA25e1OxmPNENI0B
4yahSSkQQMQsYUas6APQUUF6De8lXLfqhTZ6QUn+UtWwyKKDA33DdYLtSIamNneHiW07UA5y2e56
QzHnCWe3cgbzfja0mTaLEJpcja5yado64XLUGezNzCvoKv4wjpjUDrxTw+8ZMvkLcXvyQN/DNDPc
Ew274Mrf9hiAOflZTTqJG74wD/Jlf7nAhHcrTl2i0fzIZSCDqOmQ/iC4+a6j9InGXaW9Ce79f9mU
DgqtfzHUu1Cd8u6gvPdbHRMqqhmrno3Vihp4MIEM7ByRPa+BaxD+33haQJY8bG9avpQsUjd+MXAn
jlhKLwXzp1FteJVnkZ572NcafE/deYhFIbGZ54i2qIlIEwfAVGwy/LfZxMk2klk8uaXTA15bAnEC
dNIQeTL18bvPf5NHW671JdauiuiG1W3o+jJT5l+kv7OWk6sWZqFc/QxQWxGU6yuXWSedZ+2RirAB
dd2iflzJWo+HOvHZt1gkNPjO/LRrDR3ys3zNdsytIQTlaXMpRzHU9NI0J5DcGpKJ9wK+K+/HwzeR
kNkZY80IHR2aBgNwbd3kVvEoLh7nER+DAUdprMiCD7b1waqym6/Oj66S4wG3nNKTI8ZKyQ1dpzXF
GrNOgIUjSlm72DPDrkmuk2zazFVSQHZJkCty4NepclM+l+krANF6nFrPQauJFF/4NA7XXpBzhxjS
U8AZNuKiSxHypCoCZTCkoXs+0CesUJPQzZziYaNoYBpPYjfiFPdZ3UU82oQsDhAwEem8hIvURNNH
NtN7K5voSLLXuotVFAOGFFibq/aOvaJ3KmWgarjmb5MyYtXz+SmLpxhVQX7NWnqumg/C7GVSItCr
OmRRx6TtVzz59G/eBGlxn5A2ofC7W5dt5z9sC3buFRJyDaGO5XYH3RhPUh9kBpaUCAihedF99IjH
jRVseRbx+elRI6DPkgIQHKLkWwCKXXBLB+1PVJEYQos37Nr/0rofMpOU1zl9po+jpkyBeHRTuiiO
X0d3biAyU4gT2SjNLQnTO2iJpYixSnkJi9sWcMDxv9myr8sfq9IhKr69+Wqe+VpVSrokkH1cz6AD
K+HTP6Y6UM0NreBuGDIoyAp3o6JPJjqkIpqHGQ7b1aty7Hb2i6+v/6rxrlXbw4NLNzPIln0kzHjJ
a0ILd+7Du1/i45emXA5zR/REm5Uj/kca3oFoQ5dVzZwvLkZThFhzwsmVS9n1kHGVpTOsByjSPJ3A
O73Z7qsQ1tNmQIniemhOZnI1yNyLgyHF+kWMvsLYQtOl4elC+ymIiOC8W4G+Lk78w9o+3HnGYjYx
7djRwGzLtQJGFwCqzXEKRqHswXbKV79p4OtXKD/3JdIH6+24YPsOgnWvLsGdAEnY75tiCH8YAApG
SUwOWg66gi2ETYdGuDCP239w++XgmXHGY2e8HgRFd1i6H/93/X75ptBgJFw9yKFRjoggmycZQ/nY
ub3uTIAnfaW7fRmpaEY9jeeBczvCj9b8h79bh/wD+R6b2gCqKEDDd/zIzpAqtWFau9OQpWv8Lkwr
CYZyw+SwJsXQgqtNM7HSVeiGTGnxwCB+Kbg0c5GGDmmkGr8sddXS3g1X6T+P9CVOVHDl3dzsPKzq
BKPAaQKxt5vvg8qBlezkYuPIknj2R3u/theztl/T8Zkt7Zg4udk60cCJRAfbNWOKf6gcHtwKzBga
Dv+TGiz3UOF/NY6U/gzFSusAFUsThCPTW0ezQY2CWb38sXzJ3nieBkViqWOXPg7MVh1UFV8w0RQ6
iaP2AusEbjdJ8cNaEOh8gqmKDHNkIE9dC7hmtoEGgdmmGNXP6tYt77yhHMhS3FqYsmj++tw8Rvqm
efj8iLd/HoPgLzbAZae3KVJ+iCX3+jm0P8UTVsXtkybd4pLrth7aUm93gwQeEaO7D9NSpmLoq3ze
SoghxJ8V+mnq+ToKUNkku/WraLtKLZek7JXPGPZCrcle+DxP3lhi22z2KaaTK9YaRks7gjJjsF/Z
a+jsUJtWKG5JJ0OYhYH2BrL4U9rZsmJn0U9OGMQ/ONWlVjALftyS3Dhj4m0JMd76YlVSBiM2D6XJ
l8QnmWIjodznDcW5NlB8j0fhWLvN/3R/kwelbzda6PfQjq2sQT7vZ3Wmb/H5ZhERVKqZi7Gwx9vr
H/E1Asd6rVXu/qrR9GycYpG9QdM0EQ2OjoD3P/fj0dO6xhRZmH7YJpntgA4Rf/PP8XadlwEEBhHE
em1dpPZc4zZEEF3FrpghYKXw4po90ewYTslrsZTCsP4WLiKdiODjBUVqDqCeyevajPJPpf6/UJyF
8Z+ZzPSEmhRetPnm0sEiJpLrkRktfSLRGIZNuSk+gkCCy89nUotQI0cU8cDzzRyO/2uij42Yzloj
voeGTFPCMUXFjNxVlQmCi9wHBCRdGBtBqBgBw4LiUyTWL3XmtynPGLgKVQdXNDY3bpdGAOaZpDWA
8I1xbrouVcmNjBk/zDGgRtPUlKv9QFvjeSFjtcAr93ArjGupVPWrcVB8B1R0tKA1BLX+SGQLMxme
+oQwbviCQgos4ArjxixYeZFlo5jagzk9MZ94sf+MTO0uazxCGpUwLVo4V5YNaTcoV17DWJRiMZ1L
mD9irjYh5srK7pZYGscvb8UBMyqwxcnBv3ttL4AtF/WyAyHn+YcK38vfWEajma3pdzngPQlKrtzo
DHClXFjPY5Gv1tyMExYkQh5sU/TgQ5EZ4aw/u01WvockKN/N+mkALdS28IB6bPrszKvYgak7KUuX
mgPBlBADh0m8kfHcPDYERb5iTAY76wAs3WrSk2baew9TWrHL0y7+vsItKOB3vqYhyb351n5m2dEd
OIthaWaQMBbPJkXcv0NxP6PBDCx6jo0h8CkuYinHUXkq1INlDCzciKkuTtqMNiydwt19CJZU6VvW
UJuPwXVQmTDTKfJNCP271d2DH5eAJOIRlwjWuT1oxeh53ScZ44hnW0pPfPlvHl+7LgNbcnqYS7Yw
ZkzSHfEk8nUcTWTd1BNwA8lyyUO7wwkAAFQYlJV37VgBbMD6/lLhfy1QwWULt0VrnFNyyCv3+azG
1zBH3zl2JnTeTCTu+KkhOCvPRlSDKxS93Qw5XI8hmOzzFhX2f1bFYpsD4zIHmb0KMdCOFtUm5Bb9
mUBaBAZoRW8S4oBRe40SG4Y9NpsfbbnpvH1ZrjzpTumHXg/A7Jzcjeh6G8OswYvDdzc9cXJ0NIzK
YO22mKOMi+iFzAwQYIa4TjN3Z9C4LJGdAOkssUHRq3LUKY4fGALTMT/AWnS97IxpwlSyfXMI+9i3
NLdINyghTmCCjTqS7q+6iMDem2Gi6j2nbod59Jmw0gR3+n9E/MuuBfcxdA5SHNBvh4Jg+4yJN184
s20c54mt5F1FF1LFmTpwuP4g/t7qliVqSekcvowzv8zUiF/gahymItIIzqIAqGrFk+TzJwrOrtLJ
BIE9xgi5n/KewtOMixrFPRCQYWrN6N8Yp6EV2pD0oZCMMcM/rD2gabCO+wrxQYvJqkywRzvATv+E
yfJbSqDjzEMy18aDvs3usvrlJm9D0buzu/UcvkNn3QUbJdwufcMUb8pV7gqdrgkf/HkeZU8tAH4S
YgV6/3t3Dvw+TRbVAA/aIXWyfg4AP6re7Gn/vfcSfqhqRFkTLWy34+DOcGcpk4e7U45tZsztTcEX
gWeFJA3vCF+1Iw3tERsx4HBFwFUgSnZ/mDG2iQkrojCy582mnO7FPJYF4JXIISGXj5NMk432O98F
vLks0ze5b2zZKDzHry0CCY9c7faZz8ITq1nrwt6BsZjkYVMKfOcDhEpOaLgdP9I3ggU8w9cINjDU
DaeDMC3+HXbQpPEKWMQ/dspeUB9hBM5/ldaXY1EpmROHcDE7sRyh4f8YEz5TxCif5LXz1sFYKoQA
n4PsGk5g9dh9KAuf7OvZmj5/PHTSKPByEG28sAzsUpAqlr/28K3zJWVmZZrztELVs4LoGkCCKEXa
QtLVQHn8iXxKB5jZTla633G2TdLPC1preVtXCyeDxvECz0TSwon12U2uuHHmoiWSbL0haijHh6/A
g/Zrbq+LAWsafRK9jam9jx+D2cYnLop8IInfqnheqAYCWtduyBN1hVXn9p6qvb4Rvpcj3sb9/3up
EficeQA0mAYIPXljmI9qHl8VMRpwbtIgSGyAtKt8SaXymago2/MqQmv1Yc96DL6wZXCkb783S1D8
jhy+hrGkpY8gt57FqOHZvzRyZ0CgZGfB//tW6x/azm186L6E5jaOB8kWzBMi7jm9pT1ShoDAKH2g
N/90MSnScpr2RC6/NeH9h9xZJE5ssPaOWeaB6fTRgdPnWupQ7UTfG4rkliZ23Xh8GGqvtA3j4imN
ugHvW0jddDrLMHtF4fiXDLD/9inBTKhA4cbwqt73kPSMJcVXtHw0e7eF0pQyevW96SRTxnsI0isx
3nBppds2NFiwwvG0UPLgJnFInwLnFZ+o+HCNKfZg3WZeBGeWaFwmrKFXBkZBJZ6Qq/trz6RtM74R
qSaulqciSgRMpUAhqmrEr8dRGs4MlzHTGb2Uep+L/r5dr3keBjfkLkbn2XBS/D2Bnu+ZajJ4Y8JR
+mzQkjRBrud8mDZ62HtG9cMU91B3WBInCBrv9892x0e6lMMRuc3ER4AlwwsPYJsmR5rc4VRms/xB
uczBOABR2Pd/ywMEqa3z3BzS7TNtAiiblJEgNHvBYua9BZx/heEatw/uo75ZpKR5iEVMdYDuhcb+
AQwWUYZQhiJQOThS2cbqX5HC5Ur3NvXMNjXXiYMvzVU/CMK0CbVk0x2vQ5HPptDY6QhncdwFAx6f
bi6yQbDJj2g16j6Mz8oYNFDFpEzaEiC7dfx6CDhtn9hYOzN45NYT0iWQAQXO7+vVKHLIeU8j9MML
qvgSyfdmBAKsl9nXwepnro9Yl7GrbbAX+9YtnbEtgo8OOa76OIrhuXyX9icxgHqqsd4imGPrUVFQ
qA8RaBRXhl+JALCG5ILhuYxztBNCql9X6AFSeUo9QF4zhwBW4Jq7u7lcV3iP+lO2PfqNTKSJ/Uha
8DqE5BajdNEtgStV49f7iz1T0s6qWnQdkzWP/183boQ4hNHvhbGaY8CNRwDjtgz2lnCBLO4z8bOm
yerkQ/OGTnbVjmc20Hkk6D7KVQqD03oBYvD0bADoZC+UCYQ/hO7eqmK602GfuH7rsKr4uy//ETVM
A478HU2T4IsQDWn4qJKvNAOGDnH880E0SFve5s1CCYcddAfSZxMN5DFPzlTPgFwStkR99TeXzh58
XZCWXKmgVfI0NeKhQLoPVi1UZNqQ3l9PkO96P4a9K8Y/au8H0a4q2/A3VLLGk4AXe9Jjlp5Lfw34
cEkSPHynjIHBSc2Qkz2sbf3pUjMKhW+zfM5ZB89XZ0BElmficKy8eG0DBAFx/VjfoJ5eeq1FDqgh
sQDCCnId4lZUosNJSgn7utO7UTmOwG8ecHQ3Vouvo91PWSh7r45hZXSnrwe25qJU9ZYE452rcb5T
k+7zFAw3u0d9ozZAQE9gQM6/5u9xJeoIYIoM2YynZRldGD4m922IGjAMCVMqhvviOX1mdrrZXhla
c4zFQ98RtZs3v5VjSqBftqTIYXfOlOvLA6U2Zt1Y+gg+07AOQlaHfAwiocsu/nK5e7njT1xznPDJ
V57BIL4L58OlHfbEQa257OYEEYgH6KNkNw/QjAy4DRh2RKjXsNa8Jqt1r8d8sb9YT+nblUS89pSR
36MqrhPPTT1dAFZleQJtt56sLIv9SAGZ3NXaUmjPAAuhhO3ReKJDsH1/HePZwQP3hKHnpYjcUjCz
sDezt3pENHqmN3xyrgsXFaCADw+dwdObFfsq+UGoJONDzx73mpII8Nd10XiQW1AY+RJNWqvpEJK1
4p4HTUjCF6D6iFlbCu1+XQQ+CiBt9wDvrS14Yee2NFRH26f2ASus9Ya15xMAntKHV7AYkNTnfsmz
msD8G9OW2l0i71S9dNaKVgvPtSi4Gk9EfYc8A7DLxCGoy9u6KfoFrRS+JOsaTF0yCahX2dfYNdI9
g8gG2CVLEC/wDUIEjWizHMzuqcqEwKnAK25rbFUqjZ8b9cOuSypI0mq92gPOS+CT5G+kfVhshmWS
lVaY/W0forgBzYm/O8/81lcryBwWZCd7wKaFhejliIy/Huoarc86rjvJ4MOl6Vg8YpVfKbRdzA4c
WNmcwevC5Si+TNxNXfH3teJ6EsmcpIOgaZiHKtC+XGrQflxXVZc9f3D+2i2vmCloehR6zpjkKe65
ztWnjQmv+FjCJyfZx3iEPw0stuA5me4dKlz/PWeZE2jFyL7DjekCmqYzqoL6PDhOd2CaSS1LQMZ3
lGJcYc20ILSqdVNCADwNOXKadhebyZg1gKJ4Vl127o77+vsWFIIpdGjlTVLW9Zld3fipCK8Sj7tb
GQUNcEKY1C3H6fbaDptLAq0i4NSzhbJuvyBhmA35HUE8E9ypFfDKEzZrTK58o6SPKxUVlLFk+Wjt
8Vliyzn6ICOKsUh3vVLjWCZO+OApCrGDH6km1XWlkVM3Go1l0A41m146wR0vRqKwQPmM5FTVD4bk
TKdPAzEAtLfCmj4/eU2u/NDFXdic72K/qFfDVX5QSqEkaK2Nb3MkDfti9GZNfyQCoCgYOjI4iHno
mQZeBMFFORG1Q6qkTXvmQFpArKnw4uVtdj7rOU+MktR84rXWq7tUU61yvbkpdrUlyJl0X78oBoBB
RXaiWSrzZLxzvuPrP3wLdT/5jkYwtMauWp/GI4oKfXSSMY9U/b32LVhPOKGEtr0rj34KOnN8/8wM
p6kMUK0er8OzhXDpsjw7VJELBaxy1XE5GQQuB1qiNGaWQ5eOj1M4JIf2wShB8tF0rd9vJZhL8cUy
prirL7dUgahHC2ghhgE7PL0W+aadTXRUsrwhgFKbYlWY3ILiHQrBdsjNCuWAZr05ErOtcp7UFhAR
TLT4Hs4dvPNrDC+r5gOE5mO9Dy++qivK1wDEaQy2TXHXxWXQvU5Uvw2TarEp5/TH9uFthD/zNB2S
skNukBZOJj0mlHukD8F+ffuMhS9PcMyZTgxh1Q3EOQVMlt1Ftm1TLlXnJF2vyieNm5au3I5ydrco
B2TNEwEoYH7Z8b7qHspGLyVHi/+wfMayNX5YXhB8PUMBCAmIjUJaGB36oViLkpvJnWHakHK2/EIJ
t+ODBNhAZmsa0hJUafflnmxmCESeCAcjkiYYc4Go6ZGWq706jwVIv7QTPeTlHz4Y7XELoCwhzcfJ
2YSCBxfuwngkJc/hswVL8GJSmPokAwxRiSHOa9oGLfLA8919IV3LJblcq1A74YX9nnRXsQyBbX/F
rEKfxJEeG2ASpmRYrysarAFTk5OZpL7/WPUNpQnKf3mz8XpblbLQkwVfkMBj09s4kDQ+fCSkfMvS
uYXiA4HfLsbESDQnzYJ/7ITxZnVp5v49zB+t6hj1XW1YswfhAmlBqvY8FkpcZ9iq3k0iKbRqzgl6
Z3Nb0V94TXGioPg8iaUc1RGUHwuBnziOWbSB4r0iab08TZFpFZklct0eaBv2dDCqocYGUjhH0tFJ
WPoUYrhco8qAHMM8yAWZkr2LLWjbF0cIGQjkQQtlbmYHd8PxtrP0EcWtQL36fHuoUhWdyuLThTat
UWDjpI0kY975Q1uUKhHPQnYqmNiOXiMTC49Tfoomr/eMXJ2bUt6H232KOBfNHck+hpp/Jxz7I2bk
iZDVi8PqMn/eJCb04gnWZqW8nE0g4eFyEBlGRZoj7Jvga2ScgDViQtV/wPY2zXa79LgkE0/s3yCS
dqK+pUR2aDSGTZ8xgK/gPboF6hkRYKFQxJMOYQ08LfOwPYR2cotsxe2vfCpPAzf+ELc+tOFBB54M
WzvxisGOalhaOlGm8/dtURwL2AAoA7g8CKd8JthGsUgHXTQQ+ANu2bD4pqO+ODA1Ju2IijOFh0gF
sxbH3P+U7SLCwcL3s7k6QCQBWcg8mJMz0Cv7xU1/6zFtsuEBNCqn9n8jxd+kH88GS4hlEYl2OEZS
4mVwCOtXga0FHiOu8T2V7qbSHxj6J1H5WAO+B984tK3LFdsD1fxdndUc7QaSpk1y2aiCmylbxTxm
kOhyyZHUTMABbH9xEEJUQ8jfOWfjY6N5ytPAyejQ8NqucKCrr2t6f0PpXkIfYDKYPolpJenEies7
+bBRrcwxC7tLgSLmvIBLMXiyS6uSQV/WZFfPMFFZfZvomlM7oo1Cnw4PEC3UaCPbdtRYRUQLiOro
09qvcpXngODGuBWpA4Ye+kHFk56PvNz1sOX/TuZphX9ACunNxLt2/TBXpA3wHKJW/esBzDUZfCjO
cokx3jlOxsrJs5PQF/EvBniTAlpShmbkBhzRC/kOjttbdvT2rpyGoMObT+ZOz7I1TOiYFsJI3dJ+
4ua70qq3ekSDRptviWZ4ZrjJlNGYYzW/Zq+tN/enp8ZeYk37ux5ZQhGwVm5vS585Alqc3I0C16OY
mKweLLALIAZW1eLkQi0N+mzz6AMuioBIs3k2e8kmeXSCqKt9bX6exbHrJJK1QdbU3CoDawMUkhlq
XsP+7vAHOkOzaI123tUUiKBjX47wdkY+Z8e4WcsyilEx+mFyeZ9J7xxv7q94L2n9ofBbOJl0KbNx
MHpmZq1AodV9FPccYW40aY9xq5ciVWbxKBkKdcJx/qxSpHQkCAhGJpxypqoyz0DdJMDkiMknqJNf
pEQcAAgT4XAUohMYcz+9gyltW8F2i3FQPttkNkfNqRY1L5C0bZefrcd4wSSHxDkd2kbWMrIY0jgP
3lwNT4nWM+3yfjVJ+B09OgluqUvaoIQQnYiinrjEHGJrmQAa1ZLqX9OnfxdNpyzSGv1j7ktK3lKR
cM63bHugV9s+5PimZdw9qNx7ZqYs+LyK+PN2LN2DgGrnc+nPvZEYfyVTvMqSkvgffZp4mTXk203f
U9Dbbwj6rBagkCcwZF8Br/o+UnBl2J2iJu98WVuNyXPB5MZ49nZuFlCwBc3q16Oioe3zN9CB5Wha
Esr51FHPU1UM/gnxeDLmpov66t3up1bMHBuQHeRsBBVZRQgbyBCUjweBjl13duVPQqmtWSv0WetG
Fr1YmA0Y7m8cFgQGowev6xvo4sDclQnAZ/QcaN+MbM8BgsZNinrl/6nNelcPzuk+0WiX2GX5AC2i
78iwqixIWyrBTkFMVJExiaigaIv/I2NhOol+yCL8GIZ6oPc/+hBe7xcBzlRr/ry/DSSTgsuLibL2
KeSJsCSYyGubRcPYvnj2H5z3t40VtNgduGkNM1UhfEW/1fXIFPhOTSouRr2ldNd4WqTMCigcBEX7
Ws9yQDfjEbnZCYXwWGOdOuvOW2AALMFfj5fNcqgsk+cH7BHx7WHimwdi2FczuefFGQ7Spsocl9Ph
M+m2BYqci8NtBpwV3M7rymbsSmYSzQlA2XvyP5GZKMK7bOUy1/ScTFA+Ehh7KJwY1LItRFW4XVF9
I6H7KQZdpOkL3/CXABB/uoV/UDhqtLLK0956QTRrPxUwYi2y7aKBGIaDXBL//9lrxP45GEwI014Z
FM8GeGmbpXr2SlZVNRuOTsVoi302BIt/ehzoFP+WoZ7SgBGVKKhOhqX4NEN3qikGXVD76+EoJx9R
q+GTK+uGRcECx1rIPBHX1ztF9KigbB+MHbup5o9jDy3eo3tFXIBHNtGP2In1xMDY8ivxPkIlM+eN
xacsD2kCEMiSs/Uo0PEx6tyl5RvBJN9z7Q0chNIDjPY0xOALB25YvJN8VSRQ7YHpasTGRt9amkbq
HBvl+zG/5IEP21XroLN0Low2g2YisZf0WgPQ0gFO+YHBqjOzIhU0xAb2mJ1s+NXs8vUHBe15AeWl
Rg0IdNFQ9mbggEJtCNIv+kr+gHi1OAP1tnaeLHQ00eM3tErXSJq0uin2Co5G2EfUG+iu3HPgOhJA
ZbXnKrkvpy5qzp6K1cX38/3zAMLrLjHXuWt1rZZM4anztsrJESTKY8MMXWAa65oI1+91erSDcvVd
t4vK7Z0PoUr+j3oYNT89vYp37Wh6sxbFQX9GeKQyH8OmvADdtJvT+cu7GvVtArF7aLsg/w+ymRsX
4Tyefv5Oe05JhDtTTOHJ5refcqkVJVUTm93BOJh7DuctVC7MPigJrxTy7i584GiWGVPjrviegqRB
il5z65zyEd3PTEMABhFExsxNpxAujnHTZVmLyca4lHmg0m0+/I/0x/Ox+kNcctR0yl29WBWpGiji
cWKa3qJpIwUhsxi3ocBKnDCzY9/c2IVD2gUutBSQ/om0gFpbTThMw3fr+4QahvTpYohLq3k5zCCy
oxleaQt//2ehRDhQn6Wjd7UBLlXZFyRoNtAfWkgvV0y+hmytaLKfzzmV6TF3XNJFgfl6yrU2KMTb
oNWq8hvm2aJSu9137zLw5/s9P9lWoHboIW2XuPtkAKA62NlN05m11DY4n6UwEpH/Pq+tnLCs770+
3qMVwhfolUbBPxrgH6djfKvun1QSPI828aZc2l7TVS/IxHaLXG4hTsRjZhbtlRknwPxEIPCDPjko
SuypOiPqGRScLOakEV0z+Sx/IAWMu7S6C2KsTrAluN8QPHXonXqlUWHv2I+qK9XAYGRJq247TYYv
eKqqn9Kd3jQmsyVQ2v6Z1zN6ZjQOPqYDUlZRyZyz1PL6WLy9iWP0zWSaj19iFQ/9YdD7Ma9KJeL3
H79LqM4p80IX4I72JVydgp/bz3yYSC9BPVBWSEF6aoohFmZEqynfwv3zk/XEKiGcI/cfUzZnpeyP
XLVgcfgtOgWhsCLhSCdN8fLBG+XgaeMmc7m+RqCGFxZBj41LhrcLYJNMe0h5I3s1BFRB9g/Yvqbf
c/7GGzGwQ254rXsQMZLoa9+3uix/7laNlmPceV1qh1Kis9ZLL4JggQdYVFJAgVaobp3jSdhWBbOX
ulZGw1Gzz1kcvQBxiKPtFpK0AJmrQkw8rHIGWmA9dGnndHeyLca/mDu79tgJQuM0uwGi6kUw3ppr
49c/Z5LpYtiFSL9k3qPa504djrXFCMUpqEMJp6fIUPq1MChLQ7RNUsN7OkHMRiv+IXWG8fgwrC9X
9is/M1kzhZPsOafmOXlqObyAVCb0remMlalo2As0echoAV0oIpmsJGPkhQaDIGrH/VAg2zEmupUM
I381aTh9vc3rQ1XBjubKfumkz8sib7RKMklKN+mf0oucfrf7eCZ4aukyNF144xZvrLhgPIVMCFyP
9FPVrmxT0Ltg/zxpgrHCgKglof9+VQPUrZmZmUBvvpLiuLRrLr2uFM5wAKjhmVnifnNrH7wl9uNw
Edx96fvehIJeoty7+dSt5bbjy4EamJis69nnm+u+KwxwSS0/wojXeQ31yqKakZVftUB1Fs0PNSrz
BPTVGs7BTjTRV/+Y8GGFbfjmkOgbaJSC8t50HIXuWLFAXt4/b6DcqYpfvzqtI+CKa7/21ke046sf
TggStKt0vtzBgKUQk1E1PM9Og8haRXXXx2W2XdexIh0E1p6NzAxYqHaPLIKD2xs8eXzcFFvrXXOG
o9w7dHRoNInWYzbI6C6r1EX3hKeiIcBe1RXGGXToPbrjdj3ojmTT3PCeKpFQa0bbSF+qx7FUI6Uw
4pjtN1EaGfF4SIZUbJWlexZvjcjjMHliwSHa8w4ZomCwDIh0ZzZDt3fqUhTHe2Lj3zU+gth/4e0u
dmn5+zjdmsHCFxXPl7s9x1/wdsrZfR/dPHUcQuFEHH0j29DGpdKGMNvuOHg2PXCc9lD7wnbMheYf
5g1bZCrCIzuKERcpNXPJ8XLpnHpbU8qB/DoIjzlGSqVTZg+bO+TAzqD7/8X9MslgAXCDSsNd7eFr
VCgCqGDdjNk8k5r3qg+e99RMShZZT5MXX6jSXKBTqH0NU0AZh9UvZVokSILjLL718QXOIIm1EZbn
WSrNuHUzwNglMucDtWFxfLxsVR+q5CupTq4/fAiAuxs/uUt3o7rIdzdiDEMGJcdgwETWJOt0XuHs
eY4rE9PLwcU5Bt7ofRcq+IpNFbhKJy8Zy8JtmJzHJbWP0g/U9kdNXd3noz+y2voDs6SulBvMwokU
0vN2Ajtc8cLOBF+5cZcBE2HrxvaoMGO844jgP6Olm0psSJqf6r1hFxh7wAgHYlrgC3H1jJzFpFoF
LeHuJtnmi0MkVpsRPF86C8mVm/wVuoh6/DlhNNrVx12y7yuJu0I4ZbwBeEiBTe+m3RC24jIupzEP
d4Q2qmbD99kRKefnMXNhwA1SWua53CgL92yAn2QUv/5gKp6zRcwB8PUU1jCHQn5hPICRuTL6jQ/u
L1r3JXneF24j6b0VFl0HDSCzYm3bvmmslwJNj/wR3IkJ7V2zQLfXDzv2c06A+sEHl7o+a0pt00xh
+zj3xYatFAz16NA4vkPxkuPb6Lji2aYxktfPrYm6I+MPALtnsl+D2GrpjtcHmQTM74q3qn2Qd25w
zvu7y4I95g0aez2yZEg/sYwZCEIWy+ZP/MJUXOXpVdffE7LeRKeEkzMfMiPP7zkbUGxXTpMUn8jZ
RQE4BiGUxJZGwjuT3VaTHLk9ww8/ARKa9Yyi7NIpe4nC6g5+F57WageHpTZ+irxjUxB06rEPe/9e
RQZjy5Fs0P9OZWgP4+WDHSmJpwCKt5iKvUmMX3g6hD+K6yTCcfrA+5EBjJwtx8htA8ftIi6pzcIu
HTNNGeCkW4youdBsC/HIRut8g8T5saah0k8wL/PO4Q4uoOBTOA67jndhh7EEMU+Dfi/4GM7bTlXr
yCh3IzCgb/x4plz0gI0xgQvzwtAow5Xpy4fFYzwQG+ARTg8PpUA7jI1fpufOAZ+2Ien4nyg8/IDh
trmrZPWnuvjdlfRvpBWdcD2oXb+H7tD37Ar7DZfSvgfvz/mIhcWHFBvDYK2itguXO9BEMCtaZsNE
tlIFFXcAivA8QN/jBX2Gj7yVpPS4h3cLBRAWnvEfypSAKD6faLJZ/31TyPZZ+WUIGdsbc7M+oB+/
tNeE9ZN8QzuwDw4S1wpI6Ae0u4tCJOf6hV3n+4kINwC0S6TjgLMdmpQqbsIgqRMGMFNkCC9HUJJ5
Ks94FnUdf7kloGwCwpiVHUxw99G3ro0NPz3WFUvsGugnTis7jFL4JojxrCC19o65HCbTPXP3FdWm
5rjBzfs94yLwVm5sj3nzOlNq0UhaCaO6KQI3SB2x6Zt1yX+mDDRp4nXxYa7KxU0s2Q/sqSYi9vMk
hm/jIZSQuAQvqBNHDlXS+5RojLw88M7cukPGT9UB0tZgwkey1BmGwxVnu3ZTHL33JJ8LzL1vqzMU
mSEd5EK2aOFufY65YB4JDpNuH909ThJ+MUvX2apDU0PunT8MuR96JfcJIydt+AYjddUfR7/HnKU0
/3hHMGJ15FIa5O2hMYXRRDOp1Zw7WpnwtDlq1oHvA91G+p4jOV616nQQAgtIVZRNE9AAK6o5nD2Y
hmo2UejwLEIuANDYBNmQMIGUDA/et+do3qazpcj8vVVqPEyMO3Kn3C0URDl6O7AJ3+RT6oYp8/GF
7aMMlJQqfIYA4F5I8zTev8HZZSQK2FDlBb2EeYkiDuelP4muSaoyK1JYLnnjNZDm6Y3IGgJtkk3D
zS1zcKOyutbURdFjq2jh1XPkGp+VjYrsxJvxSQNOtzeBlXc3LSpcakBnFKVA4SzrxyI++zJG8jCt
h8S2tm3wYDS5DLsxtoz55XuE0qO277MFHpz47+gR3+/pHjHFNKR8G7HVNVufSeb8GGaNLAFwh6Nk
oHGoa13FPf6SDpOeK1sXpKRhnn2aCobejNKAMiEE59zxM1bdmPC1/4bYG4uCALtoFDL1mxIXa6KH
UFFdoQOxfyV+7pEO5clqJamztrBNNVGDTg79Sm71TPSbS6BrSQCCNvJtAoe1cwc/iv7ak98v3k0n
Ddx7JJDF9qIUAbY0hYswJJHuL3B+K8dBrOzVdzlwPlUbT1frtzBJLF2sNBLzqOl1FfRHo71QL/gU
R8eyfEcSsg/2TG85EjjybfGX+Nvg/2bMBrASkhUqQ0jgBD890VclEX78gvG8q7HG987KkWkkG4xa
nsArsBQxJCW9r63syc/zs+uQWM+O0ImWPb1XlVCywIKX7+AFjoT5eTRGUgCRWxqmcCH7QbEyetbI
J7uQeqflNWVdbd2xztLZMJ2zUX0/orU6Ub5tbhXHeoA/BvaiKufq1gTNVi//2Kbx9QJnWEztGL30
94fpPOmHMAtIFHuQ39yFcQ5lKLXya7ebI2HWIhCLB5+7uMheEgcnInxRjQOfqiebrzSK8m0Ac+7+
HBpz93ji07btiCJLdy7TLwgmBI4jxN7a1KFQLq9uhKmnN98c4XnIuHb3KnhjkoJUIf2hpkoPeTX9
zJRdROu7NcHpHmqQyEO44zafOh05W+SeCMopbX+ycnoLoqTggcT0IwA5Yfz1xIFBfCr+S09U6e0q
2dpFp3sN3UhjJKvkfQrvMTL/VwPA2prHkXgBR2kUdV9P274AaFeJ6vuAjQKP1P89yGiig8fHEykh
2K74Zdg8MCnTr6ycIIOlFnzKH651CmxEyH/SlcQRHYi5Wh3bWlZOw0n34uH/zHTotuEfbf0MIErx
tqWb6yMwll1Lvf03XCkgbpkX24RKf/QVNPyRZ2wpl39y+hJ3Yuu0xt/LSeDEbnMM8IEjtZ6RZ9Ng
/pE82fzdAy4LPkxiuZCBcGoplrL89iAQ5OFvhlzmXiYsuaLAPlALEjK4EmtPRGP9cqqYeYkV3Z0n
M1jHCmLV/OdsFhx8CEATZNHjAj/2R6pJKcg26cDh+nKQEMvgJtMwmm0l1ZmOizv8jW1rVOot6VLM
4NnAnzeufHhok/j7igmQaoOh1wnwC7p4WfRnBfJu5Q+uILVbiWisQBVIN52kBUV6IbjaHCPoO0Pz
72SItWo8A3OZmE8ywNME4dt3yHLJ+gjQIoxzVBUYjLurWy32n+kuY8YfIQaCBT+OS3RmeCEDfKG5
/hWCUNDQwwfEJltGjDry9jMAZEhC9DjObc3jggkAJgDaC7k1oKIf66kXCuTeRpzHezpZAvz/bW4G
yXxXneenrpsLJZP5x/lhyAoalgq5c1TMOMXcrQlwS4B1LDmVEyn/fuEuXyKNxyc69z9XnCHDSUED
mSBzBQoR8Xc5RLg/9luQsJhdrXPdvs1dV9zPHh1x4yyCaJu4Ik+T7ze39defnZiZWQXaJO6vtGin
FLPXnUlIY1KnHzPM/CvibRp64Wz+qy7Q8eyO2VMt7FdTojk6h2MluKtaLs1ftOtsWnZyWyk5hv0L
BDL0+fIkPh3ps4KprTVLM9z9AIy5n+WKd9KecyKmwEHLIgDwPa9IOfqxdvrCJtFUPs+9sAsd2TTo
iN3/2rUwG/m4WIax8dvN617Ob3NCFZvqArr+yWkGgYjXztfRkgEfeEieWsLGO0GcFJOEklIKjI/w
bMD/2mZDvrwCmIwLve13UQ28tAHTUqnqdU4bGcSQ7C4p/r1SgJ3FbfFnAvoIo+yBDvsVle598be0
KUoTF5FusFPZxEdrDqXiOMuXNoCH9QagcM5j59sLr81ofeko+FgVlYPvZP2y+JN10AWOFx3VSdkj
H0KSZi1q9W2klpJirw5MecsZKgB+BKHRsSft5gBtsPmGPG5G8NBP/SpLnuj3YSkkMLGlkoXkcfiU
ZZ61tqknYW0f3qqAK1dc4H8tXftmhnsyS+jHRry5HyxN1HDJH4G94ORSu4U+yo2+Eka+GPC9aRV8
FBIEGUGrHWpBKij2Bm061x3UgM8NfyKPVTF4gSRVaX6Jxm5IftUlIfLlhwJEpDJ9dWqU0VlABwyq
l9oyo4hi2pcyTWDSxX9P2sUmB/cM1rARLTdnn00bC4jsJXfOBSpFYoZ772qXNtTZoNZFDO8HMmFH
1elpTsmgu770JHq7MS79YAnzTWoUdKhgworglSrBy+1RKkxFruFHKSqeJ+o0tVeEO8dd8+M9M/4z
7pwtzm4/imYeAcUvFRCA4sGtz8Cze5xUfX2Xpd7ZMlbXhxqTjEsJl/e6VwgDZlHMIrijBcg8fs2g
Tts/ahQQQhAacWQbG4X29enAVjvzHsvhz6VWK7n4Mt117THa9koECDDkdjSjT7eZ7uzyCvMf1Vs+
wvLxzzybfop8Nob8dcb9EdVmknVia+toAwGLK8dwM+2g9fbLd8YOk3dm3ylSgCYm9qPfAKw+Qp94
rE8/t9cGilt1NiLNhZKRNM+WukpiFnC3p+J1EeBKUJRyHbFYZ+8oqd+BoBxmJKr0Uw46RJayFgmr
+j8i4GkaRJ1oo1Vr2XyqTS4r7vpjO7ShseUvAdteVdQWnEUZTlxiSAiFUhMdddxHjIMskNMTawEh
/ri7lARm5TQeKSMeSzOOI/3l4Y7I6wf6IKYhlwEdy41hGuozC/3NOgv5VXgFzOEZzE3g3q7WR9dc
EfcGLZxa580dqs5VneehJeUMXQhu0L3Dxbqq+HWtpDlh2aYx8ujFnPmqwaSPpnXfU8tk+XKPGAbu
pAFDG+mUXy8RtTcPKF7kx/0weYAG1u24yE2ll++pxcgWNlqoS0dv9/buJIBvUQIhdXyy8t3n5mwj
MJD6u21BP7kT9ubf4Ad04qqMqFHSExRb/bvRCSUtwkmtb6/EYYH3/nSjNK1P1swJLLk71coerPVP
JrDXWOFgPlRYoZ1wgMPQApgu2RkAWAWgaxLmf73/iVJiKrJK4hX9vIPMunQrRHYCqOntj5bCn0e5
m3IIRQhO47ltheaftZ84Ak+yKTAyyzGn7NxccosTGpGSgOpORCoZGznnt1VdWBM3pj7X1tZ9xZ13
NfTRy2FtKz6Ve5W3wdaf3mnBkTUrzQC9qhNPqYm9h0EDxVwZkExx3EB1KFmW2KY2bWcCVBYanXbv
A7YPP7Ekt6FnP8gEpV5+kIkUSlf72HQ8gtl+6FgrqDVOultiBA5+cl4iVsLAfzpM/iQAYXW3lAqJ
83WFXUjHHUxzOuu8U0HNWJkCklwmZDYWGMokRI5y38gEUQd8Ww0OFjXUK/D0y5HHry2SkuPvkmW9
r9RzwHqweO9E96pu1OYRiYsQ1k6BMJdSga3sBR6UmOTSxxEm0To4iY5TLoTubH+hrrH4OEo5cIQU
Uf4vvb1rm89a43pbSYJsZqVKsUHIwsmwoYKgWKK8h1UORRJo1sdQQ2FTM1l+DtF4Cko03EVPNel4
rFJsx5WHLKs6Tl75fyKPOTtaoqGwbdpF9DJV10y7ysEBR0dEUDwccsd/i9YA2crA4rLEy7xw0E90
2wX+2WNa6vFQr805MjYHA5nrrM3fHni1JqEutzGFpock3HKkw6wX57YY4c8r6DIedq/vZd+gUjoy
O4uBPo2PG0f3cB1MvA0Zap1h+/NwDCON6yXONKwLvMpzDFr0uuop17z7pWNMclSeQ5fGVfDdiPKW
Gwp2U6jMkhIqgooGgQVGysY5ACE4Je7G9GgWB1DOkDYWDD8VZQigb5mmSBy5GwMKkmE95z7svRkA
UUlI7KTf2X9Zcv6hAgZrjon/2Lrg1G5UFBkT7K+31Brx6LnI8086e9Z/Okhg/OB7MLmexbOmJDhy
6IlZokeHKOd1gWF5YAIephjJEJP6/IStV8MmjDPHFs0a9luLSmvtHm67wohHIlwbmv4M1kMyIMRL
ToTr/IhLs9MPdFYU/uzHPYvkf8T+fxG6oU/jJtKzWuEIFoSTkpvBDAgZmyC6qTeqFj31CPOi+SII
fpuRj5mtTo9lIK8Jf0DwXWBYfRhb5bjKQrKx/4YWB6TpI1t5hI5pMpOws3u82MAkiKQ78NsilQjk
AX6D4Hwf4MVBD3ddK/5EYI2UITziABTsN+3s+jRFFdmh6/By7//HfIYHMBeKbyvvKQb116l72Ej2
aAAqSTAoj6LQByM9LHTuoiFr2XmJXm7ZSEZBoz+aE/+zyf68EpqxQRoOg7rHhwbU+Dq9QHFfZyTz
rVIZk2KhN4XWCeOkXHq3x8Uz58/Iuq24l5twjvlcP+TbmDmTpMDoM50+Lnnho/B8rt0HznKcnByz
n4Qvlo4vOeMo4jtBc78d8W6iun3jjMEvZ+aZKPrXGNl2E2CEbL4KSCwUqcv2/71Ut2u0SjdZjx48
HlGAb+CxtVtzB3GAcU/DxzPwSt7/0I6+u4ODx556CuFVFnlZPfB9qbuL46MJlINE2gyvNtr54DdW
cg/ysIjGYzxM/2fbmYyyn7OOyKDTkBev3s+K8RvZW1Qj2FQmvghhfvHbPgLOEAZxSI1oTAEr05av
o2wqpBP2Injnn3eL+Tz8wI6hRIcJ+/XVuvLXKO0+LV9euHln2EyKooxlpUFgI7crusB26aslEs40
T+OTZ3G3MqZxGEr33xyqoAQw1pRhAJ3wzCnqXy1wD8BKW8MabITVbO9y09L27AAeaWN8VaG8Vf9C
2NIyGswt7ACpzeR1LicBw3Wm5NTwD0kyVzsaS2n3wDCOfOSOkiGIkUWdFy2Hq4cm+tqJf6SXeAqI
V7E2PWRIdASi45tP/hF56zgYeTPs26fAPLUGo7YDDJR0ojhGjd4efWZY0fKTFtv0VADFZPfU6RM9
+tkh26xrkJyXNRXsSUuNntwK8YAVy37I3pK/lfNdXeNoZ68K/xC7wawjpQACbi0pIAzlqskwmA9+
zEcoG84+bghEN6PLSIBdI5iqClFmbtPZ+6+SXlOJO027lmEGk+atoXO36vDE4/sNKHLRCiLZtxTo
jskaIITTYFh3hDc7zUKiZBp2yqxKLUtvm8Zqqb3MfnxycIwGcFDLQq2rUBbDBTb7kh9osHhYxz02
vW3Gf0beZbhN2i4BWmmk9ZFLtXLI0KewIusmQ7Cl1YYBiAY7TpOCYKUMkCSxC6x7rcUifiUomucj
sj9VDuxsKFPocOuDt07kLuc5AsJQnVUPypBbynt+xa8+2ispi9ppeiWoqBDhZ/oOg/0FMvgsx0us
GAnXJstHGkh8sm3GatTTD4B6buWOPbQP8lrMo8gkn7qzAIoKL7J6uwJzodeOKFmzfdy5lBfDrqHF
ogI+10Bq+/2cDaJRBPxB7k1z5jRIbiV0mlKZLKYIZADP4GhfiGGLZowSufHtD56iTGLuW+mz5zIz
X3d/RVgh0MUAqCBmRJZHb5Y/SdLOizxJnVHpVNRsqlrww3+mo2LAAwkPj8XkpwGaUQxQVaDd0uVc
VsRY4TaMZ0t1F4VkDWBdZvWEaO3M4z29xwqDUitnoh4hvxnq22rMdBE2rh9iubMHuvI94JV9Cd0h
kjflIfTdOBGEeplB99/QkOr38dDI8oNmj8vonRNaUCDdJsIN7WQw3Bz3Nn3Vq+lmFqpRFUkA17Tk
mtxmpDKTWPxODSxvERN3MBeRO3tnyxnT9i246sYEAhKRtKiYj30KKpblClweRSZssaX6DFXZrv4d
Lfc0bbb0lEynpBKOdyWDiNfaAA5ypgvQRLWBV75m4BfznnnaILpkOoGkrcYeTXN04/33cuuQuK/W
IC2MqMPFC4R5B/5milTNt9buOhhHrcF0whdP6bRXtF97PqBJvo2RC8I/h9yu8pC2rHhPECZfupQG
EvQ3q1qfXSYGFLK1eAI/qcLV0Cw+UKwfAEndM5ybDZVJgS9Yja+DBSkx4v7qaz6wnX3edoxCeFop
6c99zhtCs7nj6h0pPdE7c3XxBDC15B1M5jP+KS/eq9PLVaI0b2HmGAXWKHOieOP/v/zDBW3wIlbi
jrv76WVAo4ZMvp275QeWvNUv4gE3QduOfK0dVvQsLiAGnBbj5+3md3cFJEqs9mFrIs65mlrIKIxN
/AEcFfpoO7eswQVWM3zGak1NWVNMh/xh9HOPdI7oC515Sy/rV4sb02+rG2EjdAsCD2SEzpWajBw4
7EPAIyt+6WKQZZInJykF0VJ2zMpzMRsQH37JTzGuM3ZhvaOi8kCvKalx/oocWSzWZLt6pH+qID2F
i3yMa6rajYF6M9yw5/lDCUPGNV2QqVPBkaTX/zIoLQKPGCHXfmk4H1FP5aBzWaEFN+1PXHnqHbk9
AMcw1yAoPMV7H07vMpn+2Yq2EBFPRIvWSLYh8EVuuYjJxaBT6Dtx9lmshDoTbw7F2Uhr66dIg8Gl
bUh0WhIzAf+oWjDPOTUXiNv7qfLuvUOB3g163EshkYhX/TciaguqPJAI0TuATVz6UVakY8dPC8eh
mRL+vRK2gphRl9gpB4ZbSMCQuYQFQ2wQ2I6LsxmWSTcsYEYWD1ITgho3p5YxH9SNL6JrOsec2KvB
VXbiRK2Em9USITO7ZRBfACn3+hKzaRMuVwz+fTZH6ocAKGgUMT0/Hgj676QZCYqkd1bA0OXWBWb1
QoQV0ObGoQweT+B9/55VaTnhhXu0le0WibajqTfZ5GoiNxuaDsJ3DHIb3D18edtXI4ygslNMYOck
vwetcBddl4o0iic9B+PBgtHEu1MWRMg1rcg3drfKMPT0TMB5VAK3/VQwFl9m0pyeb/2FI0KnrzML
Db/89DRBPeLs5IZpnpX+peOccFpvnVRD3Ip6WyeEafoBdQbN64E0G5IkavrEIhvwaos9kIjI2Hfn
NfXm4aXWGDJW5/TfFYAVU3yvxpzhETg9zsyQ2wDDCacnNQTPO/13Jkx+7HKKR0jP07h/mxu8vHw1
Q+RXLe13lAaRRVplzsu36kCC24IH/a3jCUTbBnDfozIv6e2jSgMxZA8LgUeqKV9KMiaY+z9wKv4g
eBVnEyb+O0LaghqTp0RdtJLDKDIf4KkGzz2110oQkkTY1MuWJCK+rxiLRjZhppWNQ1IWdobEMmkA
Wg+vtPO3O3YCDi8h5fi+Lvuxi39nGA3itvpRN1bgPMajhfHxw2fLK54O3TdFIdzx1Zn9lZ/wvGt0
R8mqV0ByETouiyvO4I/AzcYTszMo4sUnb15qjPE+N7nCsaUC3mk5DVPvOdeoz6rOjdQZn8e8UmoF
Rk88P1Jd46HYZjuKIDw/cOf0F+Qw1ZxkxVvM9mPYfpoymrsyHcWu9j+xUSRLyMzwTezNF8NYPOQV
DhtcfIiQVDafNQGgPPveF6+GTCPcLwp+b6tu0T7NeKiabbjY5Y+rW8KqZ0jxeFWzyGqWNCC0KxFw
tjECvHjQSHEyAjM5SlQ1SmuDCpaVPK9KduMTg/T2c/apSOvb/gVpDBW+lBPaDHKrez8kNax2qyOu
jHemkinwwht8sZ/cea2VJZNOLV8Lx4v7K+m67cnddmU2iY8vhdsjEBsHQ2oiWoCcHnmq0qAeeHDH
rCBUGE/nBgY1N3LGMhJPRNL2hRRFiC7ZNeCvvZBgUzXQ2KgYwcxusUuSN3fOxT8CPjPY2a4XwwHe
lbL3A4HqK+UhgW0oQmcVWKT6iXBBJujM0zmZQdeewjXAKiMk6Ft43asT84i/PsbZ5dsI3pZrD3E+
J83Q5LokvqEp1ECv6eTnzZujrD6+MM6DPXVYTh5qRE0VLvWojiRAbnv+I7hfwMAubAQ1LZbOcl9r
nA7UfHEKWYHR4qNuNoMDEryjPHEF3e+9/ASX7FizqP3Xvz/OsHjMFvDmuIpgCdfRqvoXbaFSmdIq
lDgqfrF1Ng8nFSjFo8VG7j1tYG99xutKuyri/ZmIdHNdaeg2iZo/37x+rYm1png6xabBbOn6FqIS
nPG8PZygGM/54yEkJdILzCvhgOhrh1b/lW7uiEa4MCuXWLfME4rWIw3v7p/vXlW4sVS1rAR/x1iM
Ez7tlUyYaMSgsRz82TNqchBQsy6b2w1KwDRu32nfl15yyS+5thCeUDUXuWZaA20jRnAGBFhDZyLu
lOhxzPh3/kVfozxtA0aOQken+vz71vawn75aUIooIBjAddmk4q2MIvb9l5rHIhfGBoYDiQbj1c1e
rxuyIPaH4bGocZpIfiYtKcjoaVnnUCf5Oajo1cBUJWA9OablOBNn7BvjQF09GHeBO72OHRtJiEt1
JiL5AVgni9dG8izysIhtXaemvbcbgH5GcvqCpLMHTifF6qapV92StjIAU+Swck07NcUFVjzVIYDf
+TKhuTIUM22rC6D57RXyU9nObbRerMCDDqjuLH+IApEbr6vgfZ26G9giGsNSH0b05uM5NHhiFq5i
E/GUWf0thYkKAZdAF4U8KB2PW6QZfuG5rk+sswDeYRDXrmmymhWv17UpBUXeAoDszGpi4inBBOwO
ujoGKUqzN2UV8DOcV+1HLFK2U6ER01wsC8JiScvDKpbU470qPOcVKrQQlOPlozL8n10URQbweAQg
4uvHrTctNO+nefFNvAqbNs6XWptnRPr+NGvgIvPaKDAx2xHv8OMKQTHIGBRV8L8FJR027lXgFo2f
4wXD+X5rPWGl4zP1sKWIrFog/N6o1EmMObdBzhGR3P93BNzlkgimE1VyzeQsoZNw5ziOdUzqsabQ
pOKdQlAQj9Un3z6K484Xjx7F883vPQFqlWnmPx+Mkp+beiGkmp9InLPi3+nd2Y+ghpsm/+xcAjH3
3N8QsUTPiBiklDWCLj5mPhSY6fsLK55nezo5JW0vqSTVZM1IETyiBBlVuTg1rH3LhORjTdCGhQ5s
hQrUQUbVKhZotthaawfA1ySyYxP3EFQ1QUR9KfrtNlRoTm8WCdeO26sVwdNg7kmQDJwKbpVg9RXB
6yJ46tyiIys6jiI5IMxtp9gKyObFKdPr93+viAKbQiC3jUj+InbAnTz1mnYKLKx0wli4lX06sCvv
Gx5Q/kIlNzwR/ogu8kWgsU7qPZh5arMbDhtj0b87GZEkhgsXoPefkhlKu2iMkNy5InEFbhQee+A0
0Dve85AZMbXEuXv3dhXMXDxvxWqZBOBA3j8GY6iHCxEYEoa7ZhDrhPoupo94ZHW/tdJcRNas7OXU
7Qw5QGIS1Hribc21OMj3aTTNqE7EeeeTb02txq0VmcM1ACfKojBREN4rru4C/cHclFu8peRK7Igp
xdTofWrHZD1VSqe1ZGDSM2LT9erm5+xoR2jBZvtaimmPXdYygFPPnx+xUyDGB6DGMelZDoNREnJ/
VH6wU+KA5UFW6QmEAXD3BFw/j04OrGU7hg325GbDbkkMVYRXYHAefWznFiVZuQf1/PlqTGgDUUK0
msk1o719SWndEgL9QATpuk0xDpJLGtWUREOVYat4brkpdMjrom+yt0G1imMr3Glgf/VEoDN/TMlx
7/zuxmQgQsqX7ZM14hTvP5PmN9LhAv1qLsplyD0eg0/g0jyPbntJ3/jlmhYc3M4DQqLlRKItlZhb
bLIds8/82SDf/eFt+IHVavj/SMpZxFD2gh2ku92iXkfZk4yN6hpxuxi7aQWG14QlkcSjhDM2kvHV
0bamkePkUBI17Lnm9J4i0XGPdrVSfBZ5xK8Cyd2J+SmcOSK7d5O5pfbEi05AW4OLdbCif8LE82TN
DClsLh+mJhDNV18tCgVOxFUBZ1K24O8qGRuLCbc/RQmEMrMag4eAHi3ManSTecjigHOuw0JV0BeE
XVnHfaPzQEwnVfokTZtWZZEoP/kRzRWy2NGW0EQtJSpjScbaD7lth+0FFXw30ed7k0vqM9eJxoei
Lqqyg12Ua92lyHqmKIkwSgCI3D8ISnfo0S+burmLCsdk79PT9HBgM7pWI6gNTr5zwpJ913l8z8Iz
WJYGFOkoCXb1eGiltZ7IJArcqFlN4d/Ueo7+ILUFgwTwsckGXp79YVKcj3t3g9ZVOiU7QIYSvNTj
R2yQ7e66k1rDTUhPE/Db4TMV3/O+d804fGcXNfmM9FPMZjmtHO0zh11FykGWeSPsQAQLmd9zvyxz
kGkXMym8cSLaWc7kLzkf4Z2dWSlb+8FsEc55PxOyZ0US+24xcxYeDZiwOQYaf5TASVo+UDfZf7xu
UFg2f2two85ljgmAgE0MeLpN4J87uHg1QNcqEzXTI38jIG606EUhsXUxkoaAWW6r/LhZTr6IvnFc
vccvVMY1ISkFmfGqRDmWERa/av8WGCPs1lH7oafoDe5Btka3KKoP11dgdVfXHr4zvIgM9I1zbCH7
JptFVmlERp96dUhhejwC11WeL/z34lKRTilM5VqF1C6/Yb65Z/f5TA13JZeELuh9GdLB19eQ3r+4
2NLN3h5OEwiBiK9w9FWYpxHOBE2QI1RDEMMReq0/ArbaN+VZflG6UWSuBwhssWPugdZuJnCAN6Gb
ItgIx+XanQW2AC9LlWa+09qSWIYRnQK/Jl4gpc18fr7AmyrLaepaOAgt17Pjbla4brFfPinU/zhw
r2j/cvAJhKo+07PX3q6spRHumClrlfNKp4QcXuUTYgsFU6FnlwQL6fq2+lmE/JLdJgP3ZrkVNaXE
v6zWENHopsHTMWXub/agLnfZMxwea7rcZdVk5+yVLT4Swa+5mGUerc/q2xnjh9SV6uTeAL/BvcQi
4F9RU7h38FzY9OO8v1EzZJOGo7pyRGDOFg1mN8RJ+xEv/mpAb9sQZZWd1sPFShrSkZwXXZO3NIJB
z3MwNvhEjKgW9IEVchADqh0dtz6cgqW9YP3qC6RuYEy0PA9hV43qkEhnKlGepOypOHKakZHam1K7
4VOn5f4l/ZFqDWSle77uJl1Hm7ey4Rg92mQqDF5ksgQ9jwdjrT53a+zUFq//ELwWifoMULe0izx0
XaK5eEko1xpcC3+9i3kXC2HU1scDKh1hXGrui5fwO/wcuFZYb9HPFqDRsX2wqwqUGyoMlqBf3gzR
9xvXkJpjq/ow/WEqiQB0zVRQ9mfraLNqmoExPkCYlg7JVzP1tXeUooUuwniEjEat8qfrfYocoO0t
2ydHX7xI3BoL4tXRRN5mmHZIRXHBWPTdQKERRC3IOYbitGODS/vfPMvcBtILFZX/CdLttfIvSj/A
7RctLoIh79yiulZk34LyhO3CcbI/GnWTJtG2XcF7EmmyOiUO3mPJWkSC5wXGkYWd+CgO+a/2ZI05
3u1xbXw/fsseNB0crif+LxlsIYRUnbEoD0DQqnyvvRuxxBXvI572N4nTi3Mc297JKeQ5uASNcL2f
kgKwiHW/eNtDpPZ+EOtoPsxky2BC4IME22nCqBrjNuT34Km4mCqpwBfG0UTtFyoHo4TjwTEPK1TG
QcIKwd1BuhaAMd7ZzEgk3RC0L99pV8hJO0+qmPYVJdanWi4eq5o+uEdywdPrQm0GQHL74YEhBhVO
yccE4HX6ul8TnfMDdp+NBxUSNGfwbipSuBS8KCR4frJ8p8vBETNVfrAbuDR1egBa/XwCqwUCQc4Y
YZIXrh4HC8F7cDnaM80qPJ2XHu1ZV5/fik5hM4kxl47fk+acqq8E8tffKCDGe7nhk5+BOBEaIgaF
mhRxnpwa4d0hOvT1WXV52DXBR8uhEWCNQnlkX2z3N+CClK5HBwO8ZzJRgK28h4XqUn5R2JefU0xb
OF68NrGo5ZTldGeVlhgt5Z6L0VUcpWvs4M4iFgBA+sde2XVrkIP4oof0jvqH6gq6IB/CDp5vKOUm
6Pf+J0+egMZCb9sVnEVFZ+JBpbwb5Hn5GrYxLZTsRxNlVFmnQl2YSiy+i+YTVomoSrPioE6hTPbS
6LhRWXLT1E+g0cppQ8CrwmazUHsutjYlULRRv0QCL457ofIm7gYuiO/2iRPu/wvABdQCpPw/+o5S
ObpCEtko5ed5deYxFVrb0IZLUDonzbpk62Qh7L+baSP4IvIPENNtOzRBjrvR7bRSuFTAzldXl9BK
rsETLemKYvyZp4Fsh0EQkSFvFqLf08aRRyes5ncWGvErvzsdKnJ7uwv5yBOPhCG8IxYezzXSRPdy
V7TBGvdkNBHkEZtYjeDrM+gvuRPZ5yxqpiQogfENZv6cqDwYA4R3W/nMNSpYVUQ4MJSC+ry9CPi0
rIlFM9a/2K0Om0LvjGe89rt/QxCBThdtTiSsNg88CRiTOKGEMQQmnHHmPb/GEfDxorSk7ickY0JK
P8ugjcbK3S39l93ddvMLH+04iqO8BDHrCzj6jc1UW0XLMsMzoeEGYd+3Fh1mEtvYqQHiriv9EyWe
2uBPnoCe+d6VvhXw+x37kurHyTyfkdWQJjFjQRPmmFfx8bGcen9MFhm0L8SL8nHcll7/wl0HPGWP
Q7e9ntSXTZu+O+i34oL7JKZQLaId09OqqFLLNJ4vEduOwCer05K/FepNHnSMUndxlAJLeDmYli1T
0oQ+8Mr3R8rFhG4D2Xfn4XsV5aC+ILGeFQo996u0NAvTY6/RvFwrluAoJBwYRaa5vqoIjMQsV5sr
2rbYGJzkNqEU0fS8x98EW7N3g6oYR6qfA3dv5dw87OWsVWOIqIyJ5ANfnpHEfJ0E6jzhKUzGLNt1
tvgwuKIOp3UKIf1Sp+4kMJxX8dksBuNkTVksvM4V41lIXY1NnelLBRuU4sRwgijs8w6YClR5jc/8
xjzSeVo+GYnA88WCAst9jnWg14Md4LxBT0wcQ/eLhFbz8XQ1Xo/minYHKpkxodlfe0VBPUftkd3T
AsBvfPd0uWczAFOO4uPHO58JoYcJ0PsZFkHn6bzOSZm7uYQ7+ZBuEGm+73NA/nWY+rSY0/4iz3gd
DEHl1SqOhqLzobsljOVbPChAaBze4VBxme527HGzwmWnWMXYaNEj6lTi0ESZsB1u/q9h0FdBQ8PA
mCunk8fTYt7BUbPDyLvc3parECYym8cndp3XqmPdugX5GdzdXiOohhiuKdb6Y8WLH9yuBibzJDGE
xqG+Al2YlT7l5xbHgKMyXuj1k7ehT6IGUAPFm1Kv2m/EXiDQ8bqkgnrt5CL/4R9Zxbi3qDaz4zK1
NslBYWRFpG/2phkPKPHhqVpnyGSOrx4GIIMMSE/udLFRlnlZfjQG9c+tVrLWfJYGSx2woe2wYm3U
0km3Q8uht72g3zaVknkY8H/CFwTi98NEv5Y+In1qOU2DPtK0ioHTZoWEPLYe9iqUw+QRaE4MpbVG
tm5+2tV9blSvBpK2rVR5yrEbmYz/36XUY+XixYks7ih1HsE6QTe7CA5NGaYK1/4pVqnfCd6uyNxP
JRPhR0Q/l0kd5DR+aH54tnldEktS2vADl5bgqNZ1i1bFoywZwX0dGckAeRFU5Dn0Cnh8/V4OvMEa
2Nt6Wyfv5sPNCBT4odKE/0ZdB5lRANkcAf1SjwRapPxqfI7fn2xJJGGpNV1AOya7CqTEvdWprtlb
xQ2p9hQsxgttUbh0nhOWSBZwocV2C2JRmky4Y0C6Ctyo3N2tuI5a6jBKBFTas6Az70QlAGAoS5b2
S9SvDYkDyt7O/pzGYcjjEdKkArDcRbIUGl1VZ6ZvRozx0azH97NHCkGfPZbaJtNKV6JCbsXznBxx
s95cAHF0Wu1VZrCLy0ilD1GWN0z5xa/qRJ2++mWAti1G3M5IhxNVKer2tQbXyd+0U6IwrPr7kpTh
kbKzQeWoZT0v5u0IXlQimlA9UHzRZi5+58SI8KrE7g3Uy3PkZg5h+mrEGs/xGNh5Kil90jU1GLgS
xRZX5aPOJ1z6CsSHVHGx6vDzArnOAVnfAQ48ni+PDJs0FledwcJQRv3yJE4Vfc1rFX9IhrblI/DS
UVedPFXpOhh6sx849/mRrXCuBYU96RlQIcGpW/hbLRtSd4I32UGavPUwxv+kh0c1mdk0NmxHT8Qz
H8gMnINnSboU+0egd88IUx/NTbq62k0hWCmSRW08mjmlThZeo/KUiuoki6OYtV/23O4kaJq8mSfE
MTXBfZqAdlslc90WDK/vBx41LFc3mPP/jcuLzTCozrxcZUggpGYiRCMwDuQ9FAoxEYmZSZmxmGqR
U6QBfsk70igI4hJ1VC6Ae9ksaheitZVvEJeZ01fAr2IswcIP7NSzhX9eAGNS1gUb255JRsby/ALF
njeNCMDsZSwuNld3ORcCIeSUuI/mwBXDKJV8LPN3lDwQubaxeCPahDDTVURv/P7M/pEkE6m0K1h7
DXJJA3yesp7tCTYW6xGnxta3sjvHWHq2p4qJyR1XvVKg2+gTFR3cPhXd9qwZEY23mEzqgRYvgi0k
jb+5qYZRRIP+SOpKSoN4fMwneK4+JMoh8hbG9KnNv+tGpA896ir5mmpxu806wNIWAOfKCD5C8bV8
9KtBhLM0ErAGvYhelSo/9PyGtSHdsmnxzLtIzUZYcHD8M+RovteXitj+Ohd3ECi7W+bkCFQvhIUi
f/VDnUzwIQH77xc3/teiyisLhHtWVNDqcqI7UAn/HUbs3HoMksf4PDyJV2yqq3/Dmt03NBEH2Tz1
jj3zGUss43mHWKenSF9pgOJNRln3drcUOHhT+Pygn4UHSAfCqGOeDzFxlsXNeCN1TXDCDeD5Cm2G
bvxun+kGZgCl6fdOpCbWFzmIwUDjDAJ+2FKxVdG/hNtUYLrjgc8KKRHwbdEsztJFABrVXbEj64nJ
Pk225EohATgu/9BZfuDHTDGJkA5hoqKuRkppYXC3XrEsa3MQVduCptdLQlkFS31MtHyc7WUDVbPI
E19BRp4742nCfWlhD4aCFZcC2JOl4WkxOUKFnYC6T2+eAnVxJfQA0H/pXJQLXONuZLNA94IB0iL5
cy+9n/KfsGe6VMK5lMJkjVz4kVhrhyOnVq33fHDO7157OerBh0fMgsn+9YMgJE39X+72qXUGMIyr
fYDQ8HZ4u2oRkAHWU8IV7zQm5XF2/1uBccLI/OhW4LYecGNcFwTCLpPM+8HuaVaKKFNmMxawNR7Z
gxJKJUkQkBiRengsfJN1fIs7TvWPMAEtYt+zGZdNxKrsrPMn39/SyIDePEUDQejWbTpZTpW06RVA
2Pe7nxo5h2M9FtDqI3nDqKgkaauvsNObmsICUa2VcWTCywLpY+q7OpzAMOD3eTIaVfkf9iwAmOYt
twtZrnLmUFkgh5hzSAZcHIVkrm03ECJ40BeYZRNZAhJZxPLE51RgDR5MOpRqOnwjS2a3ht/cD28d
WpKZCcL/hLYNz8x3pK9GlEYXfKIzrKcj1fK38A6UqOrTNDBIS4mO9yydYKEfRq0tzDv/a42x7FLr
2H7q2DuQgsfjOPl1UEql5KDpcMrYarlzp4QeA9gG/GyfUjg2etkyjGOkZRM4H9iBkyhCSCVwrrW5
RxP6YsdSB5anwxX1gWKmNsyE/1tHYjYbQ08cXlfBW+kFq7uOlpbPAe3gumD44Q58l+Xnmvazv+XI
nZgxTAh63kwPsMOt8rjkidyiVq7msfC+f04DZi3l1NhlahS2jczA4erP0kofq2cgKw111Z3Qdoyg
r1V67Uuh087bpo+WkKhPAbp54xm73wRqDLPAULobklXQkmxWVnuTBAXaV/S5knZYUgPdANMLG1A6
jCbJS1A0rbz62/5pNwC8pu9fT1Vn6bkSW2J07ml5/9lXO+pVV7hrceBCBTmfa5j9VBx+3UqG2tzN
/r955kJvFb1AD4Su3uKZuMn4ZPgzjpZaKSJ8oUfOsV4EuUFzL8wxqq8j1Iq0oXTsCBxKDNkPCqHs
HYMUp7h7J0eq6fYCB5TFVdla3v0aToulPOn4wGGvXJsWWTtyUxfzh+vgSsv7WAKsY/p5+iAQPfet
p/zfJxrEoCu8XOjrYgodKfUIs6cry197CHYrnL/iIN6gZ+6lZQf8I5QS6Gwxj5a0cE1qBEn35Nms
D6vMYaHQrMyElKfqwdgNO4KbltI7zsoSwrwRofUegSYyW0/h5v0AFuTi+AJ0auDG1lBFUMjnIUUb
xAHmfX/khEMf7l+lWKF0zU3aVk3ZRk9SC6xSgyk0aR9V/O21jWlkOyc9bpmZcDNO9smqNSHvUDpB
vv/zCfgcPe7Ik+Fxaa+43KZyTnWfpKU9kjzWH1gGyqLiDc0N5KOaoAUjaxOH/BZTQOKOHWKsB8yB
nbaTnrnxKSdXbzpXIu3qFUK8RMNc+3PR5NyF68lsc77RSJccWL3nsGTOj50sJFVd7T3a/GhgiRds
WqCXoiEGhtknDQw0wmLysLiXd2+Wf4ByEV0cyNOzizSd/Mb1ISUCp0ujsyNnuX+eUUK/Ez+Hxfyf
O32mCGAkJTt7dcroYbKtG32NMz8pQsVej8S3OLCqW+heo/IRDOH5vh4LqRUFLawhaxU2dDbgckRq
/lce/WBCcz5i+tMhvNr2wS8DMBlI+t9myFmXNtD2qnAwq1P3JeCQLX30IC1SMF8khddiHygfB/B3
htMb52apbiPFJMfUMpcPk9VFoA/yOvfjVxcTPMJwaM9xrRTi9hP7B+bGGgOELsA+rjnPoyYvcCuC
WkDukqsDAlzkBBIe+WNvPqMMASr1qcMpQuIXBxlwVAzo2x8gakyTC4qcYFOj3aDVBHbCBQ3tVvg0
W7vZNAfn66XE3+UuZhFdn8lE9m1uBj9pEPu0ylhuhb/QTMzvo8+T5NoO07/gy5d0X1UEb0WOZHvX
ObzylyJ9Thb/L6NtmvQ6GmzzAsc7lSMfk2YxpND9DRbVDFPLiHwztDT+epU3K+9uTbV+1ul7bAul
3pgLRbLCPKfMyBa9x2KX5ed3lZhCbC/iLBzF1F544zql68Gz97OhQNrajGGDQ6CATdrgiB62pr8K
CgQTgAd7ls2IcxSi9Ig6mqr8CknMJSP+XyJDktSH2GEK2UIXSs9Ac+9bp1UcU3Bf6k4zCAeb3P6C
H79e3CDpQdy/dtr+ybirSo1wHeGm60qR5mzcUS7RLGBp1LiRNmfV0o8ePGeiCFwyRtPMg73ZR9ac
i46Sf1RQo6jReO2kx4lh7XCT0r6eVbt0NRG2kKKXPvY2gmIN3ZMFKQu+I2vIAMbS0tVsYXjonCTW
a9LftypObtENCWaDa6lDOLer/5iKojeZHAWfH3xjl8h/ChcxfCOV9/VR8C37HZCXquwd+9+PP1Fh
nrRsYsAR6B4cTKU88TMvHWKB32hwwwFvlHYm/UWBmwBnNIDXU/vxm61rdmky54nBot/aIwkJcIJb
62FrdUbgZHI7J3YzvSm7g/9thAnRLKCHihBtRyAV2X1fTLEUFzvMecGLM3JjLUSj7JPDYzqrt3mt
t3xV8oW3QDGS9O262zg94BEKUvqwzL1uahvX3e8xPRzcIlKQz6f8qS1TT8f0xw/fooTAjJeygKLk
YYNBCvWdnmLadGd5v2yOYrwM1BLRcOb+4Ye4Cfj6xTsd7wvU4OPgn3MkeyOjyMSBH9x6EzqKhfh4
KZhyGSIr3dt6qVbPOMRaI6IJwAMSivJ33l0/OB8eCFpHJjq8um0muNCtqbphpoOy0Q+osdHqjsK3
AsBD/6L0rvczH9l6a7RyWWBcoBYb9SUNn4Ch/tvUzJEfA+5DUceN7IDIG9ITOUU5jT2sxu3T+rOp
3PSmOJJCJazb4TlwFMIOIXnH+/axDOC7MGLjlHcWoALAD6Wft9IdGu0YOzhzztbdl7+8eHE7aJzr
XcGmJVgY/UmHAkWto0HkUTKrCcpQkG5uHLK0Pwdj4zX6S8+qRXE2ERVfsgqPy+K91rBuF5Dnivm/
MtOaIxdPJSwz1xsNvDFGxm169q4WBLV07nIeFt8J0R0JZ2CEqKjexseuTtT2QUpGMNRjBg/YmsQK
9oE3fKNPCLmff8BG3+CezZmJgNTN2/Do8QJdA5MfB7EktRrGiorGVfE3kJ+bZATOxyIcZ51rFMNp
OdeCZkF9QXnrCjZOBF2qQVZF1uPE/K1e2qoARKP60bth0M3PBrAzMyCu7HlwbUocPAkSj41iAxZr
MIDSyfxA8d8nVmCP52w3crPJ0mIKzZz/6WtYdlZmmManqG26QwfK+YHPfMs+b0yNf/5hqZ6xj4tf
Wi+6y2ujqsxQbyrYZ69X0vw/yzQ7S7EISgdYwJs9Juv6C5iA+T2v8EIjf7Fro8ee1/+a9IESU4bv
sKgFI+0GFFO77NUqMw5fTptW2gASRCOyt7atUzBT3Gqut4QZqjPJ0yuYYjJ+O7JoMIOiDWbXx2R1
aKZ8fJILZLd0c07vQ/KNaMcJba5bRvV2ICwjGhhdKXzXV/9my/4qtW7T2eoBeF2pr5mVBoyfDtEb
f56JZcErrIh6+xVKhQaRjodxkjSkGMF84y6YcMlq0uM6I0PjkxCOly20Utp1H6lBDWPqwdznOucV
Vmsv5sSSH7zShLnFytz+SAv8c/cXItswyvEXVVN6PwrUoiIDIwb8y+vJ/HAP/DXK3SZWWn3bR9vI
iHIx6lR3FQmhCnJKZxTOlFc29adGKpX7/Vkj3wGBPAFRlPfHwBBhQq4dJal03gmIY6MesYHVJSPw
yQXYFzokpnNoeiJce1qfq9I7Q7acjG4BjjqRws7ezlEtED5fVKqwj7VOw2QC/+BjAe1LTp+wcZnA
xaYqwDdEQr2sBUa7DRBY+PXktBAXgFPK/4H+Rp0JRCK0gltLSZPZE0fiDLi//MpAElnWFXPDxuke
AcKPwg/TUXgcCR4PQECZJYiVTNnJXPeG2Uq9ObEMUf/7Kl/DCa+Ai/NdkKUXIIZBV8ECrvwP12fJ
zF1J1kBjvyIbe4TK6EcuDFkcNutooP6AeBvFIEzrVZk8Y77IsvISdLJiafh03ZYDTQXsc0vwb/u1
8hK7lmxdALHKjxPJFWU54gWfXjfMe1zIoJ6/HByOY0Y2Spn/0Xq35Fd5QX6Y87/sqZ2vEL8+mdao
ihNxQLag7GehiUd36NmB8GaNmAdfsJEWNMaYeYjYl141ExEgrpXv4LagVhQldksOQwIKYq4rmVpj
tLQePX5iMwbhDnAela7ifVP8Y8KbVg5kd4eqn3KQo1/sverhGMgPZIV52qxeqCQ8/km2eT/kVelL
0kRQw/uSljD4oRWJw9zBMSaAakxhkGAwyX7Z92ON8qgSvgNZHoSLYoQE5cUKrkTaWzyZUCoQD/Jo
blVN9KcELVxonrwRV26tPr6bZzbXWw/otCM/g0FPTTxcScO5wghUrruy0Fyz6cFFunDi+jeSdMsQ
grfUg9PKrlVRTi5KNtfUXTOMaggmqfLjlVcUNnKKvOxVCscI8bgVCd9/dpVqHgXBm9+xtRV8Zn/c
qexQmaNJQKdV6lx5/xGkCLmWx2VYHQCFNBtFMopO2rdUZkAN8mSuJe+MJQVc5ojGahx6OsDtkzzL
FK5gW4nW00PekKBi9eTbLkLV+6A6wWz2HCiAIkZ+y1DtNSvTs3tY/YkzZfqCdQcDpLn9rfSB86DB
wD2Bn5g4Vj3rqPtODKfoDZO8E4ekib2JtzycmbV34n4zS4KUhbelOBycWTEd235TE8JMmHCuaFIW
LJ9KenggzUauErD1peIzPfPRCSo9If9tH5iWownDAwgTDkRDuHvh4joejX+K3pqZ8ORqBXYKSA+7
Yvt+svtv6cJ4h2GWqwW6ngZ5NXBH957FZr14WKWQb6PiMAyzDgwwPjqO9QjvcsEHs/TZ5Hu7n5ml
52JwmSMtfDcsw1a+d0dmoHYhJaXWq4PdFewTl/9YSnKHY8wMh2tS1Vn+NZIS6W5yk51cBNkeHTbr
0zaJ+2QlrWakMFyfPJh8ZSNxz4TKi7GuyaA5pW20L6JXXz3aX8vcbJF2MkLGcIud45MMUHWIXjYu
agezRAvYwH7ylHEuNgv/0ll9kH7xmkEPEL3uuL1EVWqJSgNE83z4eG8mc6pz0iBuVwQLojlJZGLa
JmzDG6Mk1qFD2HK7uMfVJXBxrbJT1ptksmcKj9nMrZJMvnwiCIKYe+impjlkW7xDyj9pRM93y0hZ
YqasxylT4DBtgUGF2YH4wlqynypHa1H/wuT7BaJoV42FnXjLyFHsI0YdTTvqkbxkqeuep0zN7yHM
uSeH4qlmhRd2xeKBS9/FoMZAgmfgXV0/5C8DgXp8ENSy9QFmRBQTi0/mXZenkZpRl4g7/k9D8WR5
awzBqqNhCamqNrSmMc7IPuYf2OozjtJ5uaHkUakd6+drJGJFq8F2oB5fbDRIBvqf758kdjIdhgfo
yb1KBkvNDeG3IKPSEaIEpwKZ0nEoww8beCMHarPrx/3dJd95BvZ9B1b2khEjyVo+OXvvqTYWZrFi
hRqTLJcFllMbH8wh0rlvPIYWOaBV61Wz8KBSyJC7bI13a/4/l6uP6pODSBpSz0fwGqsElfTS/8Sh
J33Yhgj+cZdE0Nzz/Hq8Hk3yhw+PUYklOSts0LJU58AT1haYYRF6Q6erfYBvJ9WVSmAMeGnsDAM9
EcBLvow4zRBA2xXq97uRpAIfWEcJew81Z9J6b85MqujpugLeVmBdj5vgOLQ7mxdVjtU6u4TfSfl2
Vsa8c0JjSkN1HyYBRTejvEhl5kmScyzkzs8OofkEO7v8V5q9PmEMHiqVqPgBAIJgMq1eNEtkAaQF
sYJmaWdf7CxP1qXPtbtcNhjJcIsLn30vqSQBJ6NlkEJC3AIJzfbnfihQomFJy6jvXsaZgD7kVog/
08+gF647DSPATjbP9YBZBCMWMVIug8CnT0fEtUTo0LVkS742ZXipsOA850NnHAOX3UZbc8dxphVr
9wRgXYPDvvqjqn3Mof004PfudBvQRxTHPCMicNDn68wlHPJD2ucVxXk3hgouBVCLxueNBLSXJ3oN
brfUr8H2W8raiuBaqPhMBVhmB7X95kkZNuztMazRKFVbxAU3tRlB7jfBXW0WtmamqV0DdKPPWM2o
j2Wm+eET+6pevaXH8zfSLeu0bt3g64nJPkZ4oMPuaxuJn+6USkwLbFvEKzzRtBfvcoTnxuAS8Q4t
WVrOajK6EyBrDnSse7iSuawoS/thWL1/ivCK/dExqdChA1k9sb6rzwfTKMg8oaSPEnREsstLal3Q
IvMGsZSQ7uXxFYu5wh8WPKv46P7pXsV1hjU/O+/ZVEbNAeC2dm5fzexB+Z3cfW0r3bEWhyIqj8Ma
6r8r5SCSEXaq1zijiLcmCQ04hqSTzfxGak8dRxfYLbbx0JmX6YHG2h46aGXhO7hraX6tVLbY3abx
a6ouJ0qG1G0cNHBVv3kSMmTZL/9j2Rj7LjV1yOQllfJ54Q5O8ynnDl4YtGWeh4GZUmVmOJCNiZbk
QkEoxLeXbmAiuQC9zUxSK4jvO74+DkhBFJgJvSwBDAUKlkU+iK3sDPJ8WiRrG7ck0Rr2YVbbboGi
26QQeoyUYwsTfbHQBCu717yBZ+jG0lzLn1c/kzhDHgL1IysUioqyVYLc5bRK1+OfcIqQdnRQaKjJ
Cc7n+0OgCrkDcv96oAV8fwC6kpKukziO7AZ+Ll5CjIt9OzZLz8rTf9X9Z3Ap5/t3SBq2h3TYNHB/
6vapKyFQ+wviE1YBby2Kev600C/B7hq1jNHEkR4qxGYrGmdYCDf7HpOkYTjsbLsLYOpK7o2F/kCX
93is7/C4xAkt9ZrJsFXgxMk1hV0uNw6YGi/8TUn9rKNuBDCBC3bJCTRSqc2rOuY5EkR06SIgVlCq
2aOBZPaUCU6bM7XG6Ugs3AyWOIuFs8CgrTHJ8vyv9UOx2mbMjXACGfEqCvQHjYCdrT7F47EgwHk4
iV0ogPnsJVM55DOLJeTjWSTe05Yz++LJU/nwk1tcmOdGafSkep4+7Ybnan6xxxlC9iH8anSMq+NM
XYFNewAV/iI8FbLsFXCt8IW59sHKchHyhn2KOnDJYbHtAM3yOPcsSaUi9KgvRI3Xe03ITbXFbCbF
VsSJR7QUd6pJb/bCpOqn3iGcRRwGpY4PrwB4eQFgyMgdWXIsGZ8ld72hDrf3OImyotUbZOYF5qaU
rchTLwGABbh88XpeMKrIFnYxFGdt4ejWFLG5gro6djWBwyMylCM/mQ9sJfhBUXMTBSLrVan7TfQx
YDgVaTqxfRO+7ZB5cu4fRdUeD8IMJSr0DMzhTOqXEvvwysJaCnMhXEt4KEL5egtIlqj3OojK0aIl
4dCRKB0m4ULpKFsYppuIv0ypMlGJx0mikQQApDas1iXqmlnWKAXQWfod8ma14L2q0XS4SimWzggF
l8SAcVVMrexewp16zEwNJCEJh/gm4nVa8M8P1kyVGb19dlaPUFTRzDyH+3d43bOJTFrOqbowiK7c
Ci8S0VwTqWFmbGIriYsm5Pg9dpej7tWqyv+tY9Y4BR94w9oQ3b8zAxYtq9C3Ci8pGeUw1A6bKdTc
kS9DMNToQzHCrelH+2XrZBq8VCEHaJ2V69sRGOtCo25GcHiQSfpA/42nIaFdF2FiFNzWyCpjelD7
+rTfLoCovMI72IF0ZQ4YBFRLL+UHcMx+FkpDDNShd6dr3H0+do4XKs3edXkbv/hvVf/0R1qhzuFY
JL2bctWBZC+8edU51/KqhNQ7wHzoIHGb1Vg5FKteKFg0230pTa+fi/6Lg8dxJbbXdGd4jx1mtMdQ
9LDahucXvjVpGpVISYlUWYZuUijM0wXI1/eYF/GuGIXN1oPBBJzAJ/hPN9PJ4Po57MOxojFsLBvZ
wdk4D1EpvBtisX8vDcyXhJ5Wipk0ErzUKMM9pZKIVLn/RZ4WkTA54GWONSIxyOXxEaLya+pm6KOT
bUGOhNOUXCI40Lr3+mippCfqtXLZ2tAFjXaL6MzRvuPoMaDcNdNHSTOluElw1La979wvyhWPlMsf
ckXnEko76jsYlwKC/wjdp4OqNc/de9JuvwYI6AMdzuOwIoDxWWr3tqNbzbEUb12C51dohP17XgDC
Ou7bkmeUqTBW7Aa2WwcOAiAWLqMvoIVOsOiUB4qYphblOB4x0LUE0rg/3lCMamSv/Zq2bsT+kll/
v0fAfAcjS/uuq9FIcjagukPjiNOaBxCImCrFDe1B5No7yOHyKekxYEJe2XmU3+CilwqGLCWynLg3
jFuor4k/AJzjXd64AS6ps8roO8VMopsrTcoSoI9XYs8+pKTr0R1L63lCBXx0vv5fcIHladIhi2hH
ecMvOIGyWQnVQe9pTrSjJR1C377oDS683nqKGRFtxM3V/WwjfHGeCG7qC8uDBISzuhV/VX+0D2BC
vdgwM0sQaBdarpLPwOCyUzSi/+bUzZx6SVL2Wym/lSLKo6eOhzsIjVUoWokTzE+MCHoIOhI8nIwa
bZHp7tP8pNfmq6u4bXyzxZZniAQaZ9ZblSyt2zSNhp8yekYPykddZgHqWJSS66C1MT2oysZs8dZJ
iH/+XY4daRhfDUKumEOv7xduH8YM3dWv6jfv/ee50T0A9jNOoUJbDtuE37Hrtpo76NBR792qD6EB
Hzko99PpkNbb0H6VTApz/1iNKxl31fStCAkq0OX+4jEJegASRBHl2WUkzJFb3jsYMW8GR7VcQWb2
qlw7CdNHO8RiWISfxeYeXYcklWl0KC7LVPmPxKT7TWHvk0vbrWCisLSRv8C2CxKX+UAaQ3SG6fSi
RJQcJHYfK5tRvIh2lYp/Nd7rhWSmf6ek1QRHVgtb79kmhI1ea6X8gqOdSLCjaC0gqJXF8FcA52LZ
TytHXYepNHeKCkGbw2XefQOXXS++JJ70wiQnMcvz/r1MKNbQcKyE07LwjK6d2flZxYH1SL8IeFFT
FNybg0+xr3jP2tgSm4g7ierXHpHRQOJj5iDh/K5TwPZKFswn7d/5NWU9fNzQv0WZByF1S0VtpVgt
RjAC1IEQQfZDNmA+R0ezQsEDcinzvBu1o7SdNasUpj1+8sV16FniYstsOYc9Qu4GYV/+CrIVpjj5
811joRC5UkbM5ogmduepaHm8D36zKJL9Kd8rJb5WHzXNYhC2yZin7qZWcZottXBzvIgXyOFp+t/S
iSjxJF6hJdMSmsxIfivejaeA8SF6Ug/ajZCgnJs7u3JkKRAFYVz/qgzGGIUWq716/HeG6sPJO4lw
mo+RrY79SQ44B0H0MJElrqjsFT+5Wq2hvm4iPet6IlwAEeYkXr5KcvA93Slz7hwUffvOupfRaRdg
YtMX5DQiQ5uitTmYeo4WzO39F+mPU1N8cx0+eW/llURnCrepj6S4lsjLiJe/z/njYtWU4yHUl4br
VxkuqDNLW5SglTC2/CfF8kK1WUC8O10lAMARj2dZ23lVyNwqzq5ooWZi4EMARUs1tQbAABD4r6P9
l8o30Ir7io0eVLzCwRzABz6CYlOUXBjl+oc0YLc0yIml9RQBikzBCkkH9XigaXPMnTolaIjp0S4B
YXLo1AxG0mDi/njRQ6YQ5RaVrX44vnhu29eVMiIGu40oBgEkbCxCYsmjaO5SiYEABSCWNsrouc6C
YD0+zKtXLe3oNrFYfK4PA3N5JTyBK+IiK9hA1N3je+DPz6HvZdd1lxJt3szHeT5ozuglSbM0W+5o
90tyVqBnxGH0ETDekQuXFa099Jvz+cZcSOKkF9R6F+ge4fY33iNpZ1fTz6o/oPd058R/VGML+P1+
bXK0KrJg6LBlhmnS9vxVahDCoTLw0D4VkLGdR2hKw04A8Bgp+sfKDk9vEPM7A6s1MoDZvMrMXQc7
jXEqDt6gm3dE42BheAJHpeTYxj1lkfXt/vRLBtiUWbsyL+jc2ITcFX5BMoaGu0hQ/RDHLOevZJNP
BQ4LiOcJCGQKXMMG9kXpMtpw1qEbSqBERLVYJlzWv0wUp+j/8gHhk4GRRjZHLXerLf32cKq35PlZ
gm0ILT4ufPFBIECSMW76ERvVfHKd2x/RJ2wShoNxy5ls300cbggwRFUNLd6/npV7SrKqvlO6CNJx
SPZ20hftkgW3Q1ONLGNbFUEN/OgRBMaFuh9v803LteK2EWkqIZNDxgOAjXvSHtt09OnDqCdX0kMt
5l7X8vtusIeMa5ECNEoERtO2LvbrL3RdhhhC6IxfWFpCSu2xiw9003/NO3P5eZ83CAvroypfQt2f
nYqmXK2qcXnfo/G6a6sLByJXYmAyHU10KcU+nuEyR3CgEVTjJBoB60dDtOaPyaR6P4rVTSXeWI2h
OiNqB5RXMNiDYvXFrplJUKeJbTGKzJes/Yao6vdqhpodi6dgmd8OsqlWlMT3eDBz8oKp3vGA2DQ9
DL1OlwA9IM4VOCygEW54xcNj7kjJz9hRW0EFZ0MDHmHStOx0XpCMqqLgQwxrV5ybd4/yWiSglwly
zV24VVfPKqc8qmPF6pa9CUnhmtUZBGcW1jfvAdfukaN8sVRqKwjTPX21rGQkpMOQQxnT+xKizlJR
c+xVIk1movAb76GVAs7GbIPtHNjJt477MyqTElCNKPuDj8wIQi10gmKJYMJWzjMJ3TOaAfhPK9Qs
g9Z0h7SyRqTrCR5JGMGdKa6QZSYb9ZI7Qk0ZEPJbP/6n5hFuzTE5726nTMBlvYSeuJzf23ckFxC+
2bKdZVsBT1hLuvFzsCTOppTAq7mUGH0VXNkWA2R/bvZkoYzONqRUBdpjzQaeqvtUN9B+GasRkV7P
S1o4eoiNVCny8X075GJ03NDMmIzEvCFFNVs398nXAFto8s1Kr9jsPV7EaFHvgnv/GpYvN0lwVlBp
WhXFNQoTYZmoFOti+XN/hA+pg7MxDC6NFl4XVITTDMIb/aKXYAXPm7/ONwDiWpdlENQ3XiWNuk8k
jnGCHFb+mDYSkZVBFuseWQVyAqP0483tBasMQtHQLNwWHo3fDO2awwsEHXnyoU0LnWAN+7nhtbua
ZghKT7UF4LytcURjxsedoqMWi5Btf1AJYlz52saWA8T2/qiFOdG/4oxXfk/fUjhcNVjQKwclO/Sq
ZnEzfpwwoO0rchaRiG+IarOCnD277HGj/B0qgK6zIvDWZtNRNg6lpAUc7U0XWCx8m2fbTZiuWBuE
U2GqooVjbhig9617lQ+UZ45NQcb40c/Y9g3mu4ljHofP9L9WZXzmqOqtFobWP0SGh0FHuDgb34g/
qnVTP9MXmMcfEO01ZDCEhksCN5nL4JKSw01Eiv1oHjqY2cbCU2Q7uLal4vjC3TSJno1Ao/6tAB/a
wytRIUNuMF1oJ6DoSixntkncV2QRM7xgAYRKb4FnCmdzbQRmHp+Ow82OPJnQ31jNRnNnIwzw6GKS
CI8z+S+wZgMyCzXe6fQM9f+JRa9EPWiKOb864swaCQZ5s+2g/F82vupxpnmKwcs75wwvIk9JRey/
W1bYNKa1Steg9iZBbuVE1Po/U1pd9QHZYk6t+OknVeozUQBP68VMLopt1Sjrq3M6bUnrIWCgrAa1
6VEeHQl3jcPDzwJs6im0122TSrGWZYjNPLZK0i3kwMG7Gq3HDe0JyaV/QMkQM+xRaO8NU8DBbobI
m4+3P+elA0DVrF9AWr1P/2CtpC3BqjMPOGq4+tcZrD/rGFMzoeT42n6fDRd7/8lzDk3T2ZWCIhQF
W9tk/McJhFLhx1HuPwz+2cE+juoXGvmwQvUTumRW07xCuvpUZx192vlLhlC3BD6x5QF53vMzdc6d
BArFrLl5UqdFhaTkqcDopbKd4D9BJOqMCecFBudj4JT2hlHQ6roCTOnv/YgaIJ7i6ASVSyTT4UYt
ZBesv31kHqAMfAYHjLd3UQn3RJyTr629PMDGIMCiER/RJfta+Y3GKzNXjyQ53GrR6V1GExKvbMuf
6o/bie7nfkQiNoargoWcixnM72Ecg1kf3FEOJ/oL1QcionpvMICZH79bYjxmImPl6pdeD0JNqCXv
GnCuRbP9Nn7+W1ILTlyYWzi4WPri0sIKoIAUtryd1UQwsR5nqPnXqLcgoBTheJLROkaq6OJfvlQ/
lXO/a3wgIxfna5PcCqnZhcgim1PVdMWKSADZHt1c8zb5ixPElqJDbIYbBzfJTWfxstC55FnpeWKv
yaea/+Ggd48q1ypvgv17dyEDLQtvSjTHn0e6BYIUGmxmf7R10bxTU/klpnJ273jQ2pDsAyWzSNFL
5ITlDzCrwNAA7pNj73RdYttkz3M9UMChYtv5495OdLbqt3HDGqgy0T2IHijE5tNKuw8eb7vfUH48
r3oLMbBnCqIq4vc0uPANeAlaP1H+iJjxOv2goD3IhSjCLLYPqtoCtCNVmfefcDq1TubuWgvPqRhn
GWWz91xbY5unQ1VXeUF9stzh/lVXvXhyPstrxb8SkBiwdI95f7OE6xeNkB3HOmUGE1dyiKCFK1sN
IY217KVjPuJJt03lvXHGg6RjkS9RKYXVBMsPK1YtTID0NghnQ3rCOVhzeA0XtbNyxoL8WldK8M+g
6w3IDxJpCB3D20Mp2yC1lokXkm2gork/7+HDXh+01pfyZrS2PIim4Z+0VQG6Z3CV1SihOdZIwafv
yEM28H+U1iL56tviKLXnrwp9cTJ5JSLNiSunAR7SYOuktOAE5OfKKXgJbDz6j8Cd9aLIjR7xd8jr
r4bGChAJfWq7SB3a6Jpd4L6Za5EoXDSE5aSZzzahv3WWpXOPaCtq5mkohVAFh0JXN8Ah/Tox7tEG
xZqqoSICJwqd68xrud2OLpJBuHFC2DNcKVSjQHSugNIhJKlJ0T8CpG5+InWhLIf3lJK5bAEt76ej
ozPdRPqMGY/UOLAMvajwfeffDNfhjWZNAaBsjFS2Leq2RKQLI9TWTx2vyjAfMxXl+t4f3WaXG7jz
QavsBYTDrmHuMgy3klK/oV3C/ZELXDMnNSvIvA6pHQLgMjAH7OwUhTzaQGDVoAhCOHtt2LH68on1
KjvmEpT0H9pa2Kd4qv8y2JzRUpqVsDRJZneh3wPasM38Obt7o+ksJyDx0sLIRVYEQU4Z/+9luCux
B91mspOnq+KcW2NAKAEb71wlXWCk5JEIzqftPe7da8xMkzTrxNeu/uvd4DHOBtHlYejX0Q0TlhAT
ApwzwPa1chJ+W1vGWELlC2KOM/7DAwMcUd88sGkPkdoKzZ4CEEGf5Wi/4do27OrwtgxE4AOZ5Acu
0mpMU46VHiNNTKlwh3/Dj4VP33DJg1w9cDKZdaH9dtBuogLQOilddiN8e4cPzsQpb6kR2O0Hc6YZ
i3kss7oMlyZYqqq+xnqojF0wlOPkK6Hnmm1LYBDUOnXvyUyK4nZ4X64i3WlkZuEHaw9LcPyq+0nK
5IMGSIWvXJZFs21UR+foT5jz+Iat6bUVEMSvRSe0mdD6uxDqnviihSq31RtRA4WTGVWmh3q6xxXa
6n+E0gOabB/m81wjwnP7g65k0GFS0P2CrWZyN7z0LQ1X6bixkcQj0mZLiPeB7a+BqNhiVPae18rd
xevebGYna9042+ldwv5Nk2rYNA6E8Iqv8OO2F/wrAuvTbaqWkAQqnxJcWikirvgmn2oDDyf/JEU1
W/q2nv3A7ytYDNyZuBq/JaT4UeIouh5hSN1JDbQKNM917wlXq8ZZz60MOMx8FwxKp4uf4f7+/RPB
uuoLx++B6J9tdVxDMihLqbtDPvAfGuJo19rJuzGRebwDgjG5b9EHcXjeCkOJlyWXsZa0TbVdU+FW
ctor0E/yV/dHCNBrE+fv5h6aBuOwnTsfUJUygXW/wy6+HCgRouf6MIKVUyjKjk/HbD86PTts2yCe
+EylEInOy50jAzkx6PR3efhPo1RV5b/etjWyRUXvusDdDsFd7ybBb4CROB9aB2RasnX6SDvl5THz
C/UeCLj6dXHiru/FbwZxTkdx2NuRT17QuuOLngAfy08UdygUyUcKIAVLRT48vsLeZyr36hAycnU6
yF/Ijf0A37Hk+OH/UQQRrojCD8pqwYrhwXOkMi4uDEj4L7GAZKJ8JUs4Uw/IZ7MXqn1iMTs6TsNO
PE4Je9IVRXvRJx8WXXlsE0YXyqYnFDRvM12XOcAxkSKY7c1bMWLpNLwS3SnifWoumVVviwFMVssT
Z4l+yrsH82t2VfpGmWXQ5CMB3caogVO7jOWQS3bpASoxF/g9KnTCcTdPUlzwICb1T2u0ABU43ykQ
d4yWgaeAfO6nHTwBbvrwm4JfDadck8/xIg9N+45LUkStZ/lQZ0+rSfHvr4QVA1W3xEOb1aXBbqxd
bu8ExSkJgCiKzlDlHC8B1Bn5lteGQI19TcB5+WP+a1gZkYYKQbaTj3XcHkRZgvtDK7Yc9gnFKQVN
wqxmsb5v9cIFWNDjfWSEmq7yfp1wtdsFsSBrAPUFNLZZsuyOSrzpXY2Ug0O6LX09bgHdayVZydBi
/v6OZYm7uQ8jgnOs48t3zhGq8LbRYG09xmajQIB0CVGJECJGzbbFuUG7no+Kg3EwcYFoUlk1PR1X
G6WAEqyzXBmlhEitRDJxDASCne/1cNkHwWYISIhs9iCo8yUEcAk08BbzmHtnUPuqIFrPFkDHPLjA
svYr/4171vOxXgrkiK7YthbdV4S/VZM86P5ncg4WVW8oU4MPE+jfdeWU3cU/F3gF6ZDU/jgR1UXq
wkjhTMHVHR1x+70UaxhiYzKzVsi5NUDdC24DQoeanx3O1So3k9nYEK4NRAQAhOC6iW08ov+ta/Cw
blXlcx7kD4UNF6MatVqVTwHnNWcPQTCFVTBQOYtSNNfOO4uoiWFfxhrM58oqsNYhQbN9uzBBRtj4
+Gd4z8FeZQZBi+vqLA9HsVxuob2Sq2q3lvKdS4GR7OhW4MTABbnWHMDhyuiGb0VDkd0bIVy8KAG0
6AHZdnaWPT1lWWEOvi0LbGFBxfdXwmEGVjoY3otFtwjrDOXzSWMb57xRKcvnR+/rqv5so5/DD3cf
QC/72+GI83GiJIpC1CdUd8dQbsy2sYmo8DRFAn+GjChVd30Gou3YE3+oI+XCW66Fng2DSdLd2QEO
rfIV7vgj5wyObjR2TVxj43RUYJSEuzPfx5MGw3e5F5pvccFyNeNrggvePeXxaPb9TPLFt7TUlQUv
25rF/S/RjnOMci5dI99audbLI3+ob/XKhgfpXtTw0iwoCuuT/rF6XngLuoIHr8HIq7w/OD+Trpj5
v1sToZH31YnO9N4N4+M3xhhqgJfHdO7Um8VUmKdayR9HJtDAA7ns6S2Jfp4LReBFHXcr4ddLfO8x
BTqHXqJfcDgrKdNelVyWHrj5ofkoveuY1bdbcWZfBZVP7j0Jgc5AyoJ7XJSZii5uj+8es6jhRv1H
iuOOLXhesTQj6ggjVExSqoVEKmxjwUf/X0Gme488A686rUumg/y8GzdljixeUAr4quuRP0mUktQQ
3qyy4yIiHVq+Kl85x9mvDdrNpYeG0h8YezZa2bJQHlTrXZqDX4q6Vp/3tAaUFXSSzzZJkCjBiCKj
Bw5zOMbuFVDeAWatGqUF+rYqbYpFcsZFW+Lf27EQG9HnbdSg1OwIc2VtWLVwL8sTE6eYgXsbCxWN
bHiJeaDXgGyZlrA2NJxKbDPlfyg6E72sBaecvciI6tkXq8jka3bXfjkbq8VMwUG9bLSbNrmYrWSH
BIIQyiRHORzkpt1C7lzFI6XmxATvEGB8JqyFZlUQsSucfSsiQvKt/mpTA4uwiiaVW/cnaEyDAc9/
Fyj6NaE4u/jfzrgp9C63Ful5XV38+br8rTNmbgDkadqDfKLAZPIL+LgwxGqFUOKsyUHkQDYXdUvv
vcNkG4sQ54ctRLiKynvd4+iG+jrnsGD3WauOwrP2aK7KutgtBcEO4c//bKhzNZ5PPvVFHgYByb1n
/fm7twftP1l635pU3x8eoV/19AbDaSKAe/wyt6vrEDwQCGWvIn1ogV6ap3FJqeyl0x3WNOqSdgoo
grcV1Tja5aWg2eg+lzIbRLsXctQzOoWwMA1s0svPEerH6I2YnYY64HTcR4sf0JD7LH+ddEPPJObQ
dtlI22Qsyj0ZldM2G4Cb0GN5dcubGAmFsE/kHuEi2ImuZmc36lBkk/DkWdantjwpQeGTkynyIEnx
v28Hvxr4t8yrYqi/TOH0T2RyL++3Cv49bu0TmFpGDCjfLi/p7FrM0uBYjeu7yHV2RmyteBB8yJCd
ueBS0Ph9hSKEbjMKPGjQ+RGiw5o7VuF0CXnzXxPHXdMqquzxIRIo9hMuQdTkWrIeBpvdThH6XRLl
SAheS/x7JLzqXgd9aMj3wahFpg4YQaioJGop9+uEMDak4LwODLfsRJTdRxTAJgxOEzPactUuhqog
JD/tMwrdVg/HauH1tx697ASyagbI6sBp6IKVSJfqvPtigbC64pZ+e7wUYx6/ZCXN8vOt3dBD2iRe
Yg7ajGppY2Hm5K017/RbyRSJIGMWc9mQELzls//cWWjY13HhGqlNB0ByAflBBzoU2p1cWNZV0z8H
/KYVfWt5obQY6PTCbOtUVY+uN86sdfbo0ThLYifYNXhU41hBycgiocob0y0thxWT/+RXdQe3ILU4
0258WoCzOz0X99z+sa81h9rcsgJNWhNXVYe1reB4GxzrN2QIo0YrDKHynZyyXOEIu/wk5qeT4DwD
Yh7+2kwJNhAUIT4E0P/980naiDoW8641rBY7pMnnl3UPoNcL7k0h4XguRP320eewhs3e6R/zE0/S
ucZhIRwrG5ZluYJZK/bzsJFtD4CCdX3JjgL6kYq/yKAesR3+6uZn3RzM0uLY0iaw3KrbWWpwTMLc
ZuktZkb1hFNHgzZRyym7sDKqoSbwYoWM0fWkabe7lBlFSL2aRLyoL2qQnbJrpk856qkBz9M4y4uA
jj+dbC4POuM0/c1Z4moGpGyaBbKY99+eizmMYwco+93GYAN8XNdu+e6fhkLSy4C4RltZSLSC6kNw
alQWCvQbEQuijVdsMtxAFfB5HQzOxo0I8I9NfGe4yhEySPWkBPH/A1xnCeIcgCC6yzOMyCQextG3
o/xfGllY2T/TJ25caQiLDFeWxKRF24rV3oUG2TkbYx3wn3h4zgJFF8AngkgC6u7aQ3GNyk2C0h+x
UW+XabNbnicT6aeCKpgrXEws+6ZCrrL9MqP3Bo4sNMi5xUxOungFbOjvdOeK7yzENsSCqJpQOzRy
bD8g08aKd7CwOnLMbDzOs7LBwMeAG8D4VvysQX5xfGqGGzcakPEcjgLc0pTvd2lvrIZWHCyoFePw
EtfGHg00b2CHbnQneFwv0rVxDlxEos+e5OOLfMc+qMLVgQl6MikY1wQMYWTDVus4rRbSjtRoNOjk
Hq/6PZBDjHKj2hG1T/AlUbl6hBLsEGlEtHXIRIOSpvB3CdD78AYTqohDe/zox8tlU5x2d0zkMb+L
pZ8fpHsA/l9rxxXVdI8fCuSlUeE1qMZLB5YvAYHuyLhi6KkKq9k0lAHw22j51CgfODc4L0YG8Ir9
E8MHK1u2pb+a2pnjPjLLQEI+T/iJn8C4U4ik6Tfp4uo+BmZc0V6AWhiCTDEgXMV5x97wwVHPbXyU
SiIv6qUnfuavtRZ+NG2QQu6faTnAR6jz89it9h+k4ANjXKB+zffKPdJMu54UJ9vxxxLfbT02F6j9
KiU9rF/4Rhouy0sgMQCcDtuhvV3++8Z+KdzZrzNJ59dmEWLqXZdTDD5ZwLdAIBdf9hzRSckzzZOp
afTilErsfxfUs2MLjnc10hbPtTl9Lt+E11Wef6Mfx6tpAu6mkFj4LSQ/cHiW+J8ne9zefVGzHdgu
dA84jdVc0iV4L+DWrQ0Rn2k/ZI2TYdhKdYKsAQetKD8p1KVbI5/t3xpOs0cJIg1z/pdNQdFFd1R2
uWqzoacyn7X3wT1lArIWXVflDvkegDabuMGrLfySKZFtwsX5hbPdO5418NPx0oMVuBWVOmqmCfXp
8oojq8k1Spp9gbVoXSCtbwu+oLdMxoEsAxMlqQq5OsEiKbdLg0qy5v9WoIiFlcC3id22vI95PQX8
cU1rjsXZP94078SUtoG9t9nAkt0Ib73aLVvVOY1U9/POu/iB14ab3GjjWMby21ZyB5wjvVJ8hm7G
TaEZTspdnsjDakGm9yS1v2PeVGYwm+0J0ioEL7l9uxITXjw7JlhxM8wR37cGhMjpqBoBPnE7OOxg
+QfsmeiKWg2sjYIfidyIWiktTFrPi5in8oC5O05Jf1B7j3KEuRG4GwVNSdYsysd0/ibYgjk8ncb0
QgLuYj4+y2jh8Lbkdz1pPYXOrVbg2eD/fE9AuYbOn+2Hij2Lh5kU+u1sgnLbvApX/jCABYSoRXOJ
x9f9dv0L7eo50PVWO5Zt8+mC4lNBWOSPqFM7+5O4IdE0Abb/NHNs0cpNCz07CNX3YrG3uUx7BKQi
hQC69HzgcY+s+uIbNuLzDkooeW04tpmsM0WiLD7OCjmr5q7cVk1bkyruKgO5HtLM5cj8VvlAeiqg
0dOLsdzTAtVtUUnOmcoetaVNg24wdwKlS+5UOAHV8GvlISnBxHHrBSL0g6nBVcJYa51LsOHCXyqP
0PmIS46ljjdWIWsZkLA7dhUezWstUVbjcBjD9sMhCEAuNpri8n7bMtSaE1RVVKvkjrYTbjcr4ZaQ
7XsUpGzRcGAq7YbaodDQ5LfVHy+65fPeyOQAjKf0oI/qTCFiRnWTuzAptJiQiT6X+UvIGhdKhq0z
0DzRQkHLfpimePOI8EjJ58861L8wNMOF/FF6bCd97mQ2YrxRjnzOwEzCTBdlkTwEgmMg4UM+0S0N
GYIlDjmGUqwmapnFbqQVQBUu0W30E4K9L4vJQLNkt/EwD/lN278/BotI06s9vsMhQneCN8aGmoTv
CvQE6C1+twg4lm5qZ0zfiCjqSZ7sCY9Z+aoNJBLwRjcEXU2nO7PDLHJu7dQKosYNNGZ+LtToxyqY
WGpJmvR9UMCSlIebB1lSsNkH14LU9Kxdp/66/oVoxc0hc/8to4e1aodAyQasAMy87Lwj7vf1mZUw
2LIK2fK1fTg2h/T/sD6WW4b5ofEXo9gJLndJwqEz5yvAQtANlliCaDgrXnLQaAqF20lH6P7hfrce
2XdfSVwRxNsL0BNftOYzih+IU1L4RSkLqI6uIJYGAh+BFATwhNxitWSeU1KL15JaIKGZ1fw9ceve
mrhCVEM+xoZpSE9VglPCAViOKlVrrecGhVoVOfmqIhDLC1aHRxXi1yznA/Ckc+U/qeBMuqBTse6g
cW1bdGZCYJJMXXEKHESImyvlGxNH1D0yY/rfjjATPhK/h7BfZ/64UTA0Jt5kfsZfFXqv7YZAJHbc
raxmT1uE2al1Qp9A4XM/KRtGxQpIMmshOXS3++bWupTQBEtBbIpdVE9jD1i5lRWKLcmbUcDM0tw/
OJv95D80TZZiIaWUm4FMr2qebKkojV5V3zitkE4+5/Dx2RCwJCkYUW5LlfDWnCTp2qKLEWQE51en
J/XltQh4qltWxFAmPBqI39+g8ROb07Z9mbGQ1TqouWJ5IcgmlBpAWbZu9/irc61pW7aEqhItDlJJ
pIWIzQXyFvwqjnByItUs6VudJbp+teNW2pfj+6wNOWiY1NTcWzKiR0aYovAI7eN11v4Qmf0+Q4e4
wUXbVU6DHmhqwkww2ay5qf9HrmazY5Nch9XpGqZiZ6uZCuUDacCeCg1sdh0xSDSay2uk7YprAI2x
DuKAngmhJDNvTTg8i0wT77hC8yYCcOBz90WJ+4dMQSksIThz06kVNLZW5CVI3mrKHEeGHsfSUJYX
ZGWNMQNwQTcorG7zNOzP+mnCHCZteWpUmIj62Yrsz2VUeEOBuMzFPVCggFd0hfd4s2HZhPw21QA6
4B3wz0XC4h/eKnbhCJUiJWRF+w1Ea2OuQ+R+D6cw44Hcnxa4EgU0WJLZraY4YxavhyMwlTKLfKpP
G71slVcbzrXsqhTyn1uc+T9SIeVuXgWv9/001481YZEHY/U8F1Lqvc1yHTA2e6bzywlRKQQJ2hyW
EmXnfm2g86I4DGIPuysHk+RpP47TQJ/7s/p7nAif13Vrid0uB+OLkJOtZya+BJFg1H6c/ykwugoo
wZWEsGeaFGDrE2vO0H++0ndRtgai4PTL/m8Fbi+WFG3UJH/ImkgJjdFzXlXfnkW93fB1m7fXedAA
EPqdLcEYluIrNSS+Ro0X77VB8k4IceXjvzN6zHa0RO7UllpslScSmsW2tMvUzXJ6G1RaS52Xf1tz
BcbHNKp7mXjRNOEni71oB1nhh65nm7NnYy21yYTvGfou/CKNgQxttZ9o467Y42DZmJbLmVtgSasQ
Cg/XxQYzCfZEsYh4vQUeqsOn6Xd0GIO5rkJCk/6jms3cTcD51Ysa+lpPADWZ7icOLEj5h/NMcH2q
De9Ig5hgjjMJuzasRJ2x3lJa+1MTjhcJYw9XsdSWx88aVZvfP6OnsTd4YLw2RRZ+lFXhmVYetkg1
ydqgkJfmnffE+kgM/6Kwr04ULo0sFKlrXDbG3BZU2DN+JFE1Sa2P1m5ZpXilgX9fKoxB1XQEr8EK
vSjzUJRl8F2UyXlgYerhU4lVucJ2Gpw/0PhdYeOU0ZmSWxfHX8BlEdvUQzetq9EHBxiItuTT9R1x
n+no6S6loVHj9qHafDEpMMnzsPy5uQlolV4ycgHPcgAxNRCzPxWcCeYc56wKsf/rAtEPaMJ+1QJa
s3Z7dBWBCOgOqXVEf/QDIqqdW/JA5RpG40/BwhSX3HJaB5FcF7JvfffgHiKIMoWitOd6RhAL7v3p
4IdtCbcHPeZk6vAz64owjARJBfuMe4c8q9Xa0uSyvb3av745KLAOp70k1cwx/cvXgi9bhQN3ReGj
PhKd56HKQ57ppjKiiTMCpja0KAk/kScAUnNWJRAHVlkbObTRziD/tPIOCiWTjWX/rFLJaXLROeAH
x+nenCJUV1+V8exwuRCMUCcgxdZvKM5K8k8XLcDl0fLi2WHnDN+POkGSeogQ6/cCx69C8NhjHtHk
LG9sFpGs91K1HTIHCq0HdXlXiuKQt/KDWM/rGWP17UiLYlaYwmNXf6v1CUbo7YVfMhI+A68pRh69
y5I2YKH/JQQjadG0bR8vrN6BdHRCyjK3fCnuTxn27O99GvfSaQjyIBLKUUsDUMrwvi1jkeRloq3j
lQcSUoFQG8cZaKFbKnnZGF2KrTIHFpZv8/ep5YFil5AFsqCXqhfK4UDQjz9YRlERMxnWIuFAziqA
vPVKGr/iO0DpWHGuVnaho8mQuGd3J1icmU1sGwahqtEBYucWCTWtWLpcYk50GXwjqWk8S6ZySR49
5WaEhY/REQKt7BCiHfPkrDHYKaHZQSD6AXX1skQo4nmpJDvC80/OkeBNbB/ds5iaUAbJuegdoOVK
pqRavom0e3Fb8aLjzu/VFMbjpFdoLHrnwQvvIjyzVaSn47occthN/trSpWaGzii0YG6m6m4SGE7Q
uEKD5Dk1AUy+kVbLiHJOKELCgH3IunBqEzJ/YlGreVLhXd8Fzk590AxM8DcTxfqdBqle3sSzKHgL
cKvpKzctL6dIwO0tM/TBorqt9dAX+UkqEdhmAthX1gLRA2DfO+kq6VaYC+VeG+XSVdokmitXntxz
v6rGqCDjyDqORDMSgg9UCHRn/JRxI6CGOMb0bECGx4uNBHApycYy4K1rGBQynnhFcUk1OF53Miq0
h4OukCfRg6cfre422436iZETlB5AwUtpGTKy/kFQY+v2seYz5MBbIVYgnBTQu/p2wwGHayRY35JA
cnA0FVYCcudkkuZwg/q+3o+lA+wKFWf+DQQ27NZgjHqGboSDvZ3jD+905E5PaxDZYCyHvclPTfjV
PCNey7qGosBC5JhZbUt6ElK7L/vIlsslrxDunZlg1GkQ5g/XXLEOnQYNbzBbqZBB7mdBlTDSWabh
MBZXKbXsiGmWzvQ3Sbsq/Z5EBtpzFpeH18dgS0LdMrpEm565ehHt6XEC7r3CiY1kCJc3hcKHi2KU
8rMjHDdtuJ+M51AGKJsXrBFtJ3po963RpLZmWJpR8GFr0voSoNkn2wW2j0RJmGXC+3DfgNtgWh9y
ey3ZaDmikqxn09+Qc13WeUgZYBBMoD8eqANpy6yog+QZoq5sRD+bBf/wW6YBn9G7lJ0BftQupw/U
2qWIia7UYfAup9rH89KzU0OgtxBA7Ane3ttNtmAtx5LUSTaQKdSoTc3q3aU02HgSJZBxsXQB3P1R
30BMt18qmmUh9Etd2xsrfDUHLBtxpWPDD38R2CuulMRpC1Nnkb6hMbZkJSDDRvJ3mWDbDagG4UcH
p8mbZKE19HfdSsTG3g57pjYysdd9dvtHpBj/R3o6KNtQ09+hr+5XvXQl5Xg5yVuQxJMbyX6jJNqr
Fn/2y/l2SP/sQ8LD1A4BsahpzOylcffDn68ChpPkFQVZI/s52OT+Vare+DLRODI6N2rw2JtHBOX+
pJPTd+VP7qYTftnzqENS1AVKCGI7l5tiLfWWh/kSBpawPX4p9r6vSeTD+23IszXwl8zf6Io1+kvU
Zw8n4YThVqhhq4f2ELZkhAzUoowOBXWi/uu1h211ltnMnwvM47bBVZlRGcFZ0OmWYGjjxPoM3/Yu
U6gMc+vJ3B1MAR5W+p2j4pLK/6B1gxxbLy6y1nfaN179P+gn5V/uhkq7zQdhWgmf42AxaVbqYSGh
JBbMM4IRL/Wh6HAgfRV8nJOFXvGPji7htIhI+Sx7dZy2zBL1tq8QXnQR+KMy6vHuNjt7mPYNm3HZ
YVg78EhR4ulIPxaErOM6YV/ChJGeStZuFWj30IW0P0krRVuoDe9d0nogcV/vRlFvv4SrgLsZ5+A4
JIXBql3wgo5qSjZnrU8gq3zQ7CGFq8ju/IEc8TzL7VoDwpxMek9OOfeBjhfwTNBsuZKZscVbab2h
8yLqvEXwieLLFihDsvmpfm2ksReCJ2YHyJLMIPziB8yoQiD91rODoAOpr9MOhcjlhILh4rSVIg0O
fjyI8niZqkKMlJrxloH6cm4y1NJxko3LIP+p780ptVKNUqAGG7rql4ZRQkgxxVNFd/8CipONPEoc
C7nlB4bs+AjBSTTPkxYP92YcODixlBJ+St36ffFSPMVk4malixRltwkeH59tbJ0E2YuXDeJh6xN7
KMJ53HBP05Sy7d2pzdhSwtV7ebLMQbcr722fEFrMxSa+dufPT/qYnfCey3MlkTOdK42vKd8shwtv
TKg28xgWtzHb5EaYkFFrWfVU7lLjxNe62ucwq3BaGPakrJW67fLUlBvIV8njYuBMpa1VBgQSAqcX
kJNkM/tqfUQd+AC64ljal/QUl3y1vzauc7VGEc8zd5bDXyCOoJ64IOS9V6zReQO4ycmcthhk6i8S
M0NrdqXtLtnlb34qwA0BJe2546jm+hgIDHiZgpQNqZImdFHtcZFhHePjqQv+m3hx5ACHioBR8yg6
f03U2lvQtA+yaFxLZpW9fdJL4cgbfP2RPLb3CvsEj7uNRLDZ5yzvjFOCKiYbI92sVPdZG2Drf9u7
7AdoxBFajt6ZakMR6VhpLnk+xulHEf+W14LTz60syMXbYic+bJ/XSvMNt5MTrBcCxbx29P4X2STF
uUCcR896z0Nifb6tvAsqPPiAFaF5QpDOrP26GWn3x97Ie8tYaE/Bd/bscVrrCD8EKg1aCXgJzUN0
a47okFz4/L+rSknV7Ri9bn+xem5nKp+vHbq59O716qt8XLPed9ABd2gCOC0XDpe1u7a7MbBF1ltX
yXMGrUCocDguk5pBIjlU06d1xP56ynAaeMSyFaP3JOOiGo0OrJ2qduOItcb5ccqDJR0JPpT1bi4Q
BR5sRfIFU5HB2MCc0GIGr4IIKR00jQPCJK6UN33bMWyJSZCI/i2Vq9kTVAX9w6aAdJEQNtq/fdaZ
pBPVLTp9cdojg29OGr2YtDSphQXXD+P7/V1AYcEY9AVo8TC675v8QvIyvsz68ImR66otURrR6FDl
amKXdugIga8g05DGkxeIioojEg814LCH4bC9V4/2CX7cgw2dqtHXcw1al9MMyVFxg/KFrzpQa5ay
ECjyzLg9aJq9P2lycfiZaH97vaQpdDqvHpI3W7SVODMTS+pmeD8hPzW6dfjFF6jMK7aiw7wa1oh1
A5wtqpY1aleBYjGj8iVmkkZGVpiqMeEF8/RknV0uZIs1QuE5x2y7g0c/NUd2bLV4vWpb3T5C07j/
gSLWfTlXZcStp8WnkE7UKExYuyAIWO8jVnUdnvd9qRwho1SgUtYhpGICflF4quRUJFNiGEIeH5iv
ytQ7NY1/HzK4LxlkMZR7nX2tKWhYzLuP0LMirucsl3Gp1n0gv/jYwBQw9BHdz2gd2do7lzwmlqJF
+lGqUgKWwV08muaRgihOgqDDGsYM0eJ0Z1F3GVAI/JSs+OPnFb535YOZL5bXQ6+hp5nJJR8Vt8JI
JCLvoLFkwPziWOZhCemqgSrkCu3mVXiDarfeP84C2XwoMHTLqAlisIPteQCEnvzmWx3p442eCQY5
NquOPUT66M69Lu0hq2aPjhmvI085aBXF4U+CT52i1EOA0UFaF5Fb5Ux68JLsMr4ErMuobs0udTyJ
o3lVFuP8dGuYGL++KoiPY8kWJjTEje130tF7tGOLDRpZy8f08WD5YlWOXhBPsS2zfzhOMuE9LufZ
9YZk/raHQxM+fprUFVkw/0x+czFpocqhCEg49woRxQnzRCzG/PLmVlgfqvzVtDPqhF4dM/ZUR11Q
PTu53ECIfYg00jE6XeCBzA0M67/LPA545+GcrKPzqxjwyFctiWKkKt5JBGeKqZy8bJnfrTXadkAH
QNfy5U4l1C52plAtn6Oi9wi0JG+Mc3YtKj9LKib8rWztrna/YYeQyzkyvb1HrtrpghFyB+kBbAq5
Nej1xlvZEvtdWQ04CBubwT0T/VtEXPlE8+nNVUyvcsyXoA1thsjZVvIdVQrcfga/oganRMxe+bji
XvZTUlWi1lVbcJC7Uzh1u9UWg1VX24izcRhrJEwpUn190hsKm/8ZUGQY7urXNkvMkIOu6DvQatgW
b5IHx1RvYdQt2MmoJRh+DoxHiHgmOb7i4RAG2DK3KN4037EvJ+PtFUCZfY/kU+qfSWC/+IHKDadO
UYKTGx8OjE3inTgdv9abYZW2bQHnT31CcbFIU4AY8s3eEWzFBuKTWSoV956dW8xv0EIsOBrDoc0M
Ukrc/AgBl89S10jCTomTIz4f3oFFGi3THpNQWaEtjG6+Ml7JRwp5cqTHuCDESSKxeLySHYr/Wyms
28gda1Pa4eOFtFkOFHc5z+O4dVlrOTSvHCTACfG3adEvL+vi7mZK92s1/ZSW81K2IQjqhtgyV03O
44VQgxWpQdz8RaRc3ZH3KlKFYANTp3OycmfZ2or7xRpZyGxBxHUQNzK/57dSCHhQbbcd0ng9ysvL
3JRYHLNMRojBhpjAcChO//AbOmuvRECNNzHarw0yES31eCSjVS8SVUTCfWqI0OXNT0haCviDDtaW
XSvidhx2Trtr3TQKjyJkjDHQZxeZt89ZnmfcpNTY6wXjgU4KbWHjj78yHjhgXSovzQqcCN61lQi7
OGoEU9sZfG08xV3wQI+8VtO0ghQZaf1xxxvBEdtgRKycv661Y3GJny/WEy/24bIuB6x7ZLJJ39eq
MPyLYuNePDXx32qCR5I4fi0yMVzPQOCFD25ivj+p2c5nIVOqDoB8rcGCj/2if3O+yiJEKI/o0KOA
QoypVx8gNA4YPFifAxZGTEQWRr1ySLBNVI4j4JDcs854ORpR07RUZUVvB8avdXuPibeQSmaKm1rW
M781wnXWRalFaWQoOx2RsQuf2jJToZpO+Osec5J+2PuDbeiX9mjGWPvA6ldUVKopcCczg/ZAf5Ci
E5u6lhw22g1eHs6mnXYZwcCNP1csv2ewcMPQ8q4Xb1YL2a0vJfRktAFhOP3LLvxb8N2Nb3xxjZ/+
gBe//YWKINInjPEC4R37Mor8TnoGq4wunTDsuPg3eXD6mJyoolYoZVJxAy90g5xJtks+OnzoNAw1
WNSc6CKjwkb2pZVi6JjWVg4ikYmlXkw/pb/RcSUJMT94FSxKHoYkaM31/K3/yemuoL2gKhVbeOli
VWY+RXEVXn5o5ch1I5FJP/ah8S3uVPKymTIoZI1eqrvl5AoS9M9r4XKsX+ZFAYF5AGrmsUnXtNHg
zEyOt8uH9Qni7M2FDn1sLIQEi10lsDgEcN095i3KbUu+qJ/ydpv/WneDsmqsg57vmcrjZPG8+HBL
crI/5dWe7aqOwRZ/F/oZJUHXCylyNU+GQZNFPrvM88EsBRCqUUOG3Cboev7ZQqNClUrXNoT6Ja7H
0RsvUxdaW7P4FPIpYsGxl8pzu7F6dwCaDEUt1d8iLgdOMkWY2B5fatDJFGkdv9wcfeVAE6G+62M8
+oiiYEZOCU4Rkp1J1xA4YfML1I0Kg/ana0eft29L8L7tUMpbE4NQtw+5e+VkYViWzsddr8nlBYOp
LOqBuAU1ai62hhGeLTXu/5Ox8i1/08SK/FxJItBK2OW+HmkN6Z0vsLNsvLEq/6/73UppzQUywO4N
vA9+Yi8g64635zOBJZawuDj7zEnDoxX6/IAEWasaSVB0jp5rwMDLGMd8yjoKsFQ/72O4QqLfzw6g
fxhMMPnvgEFCkwqcVI2VWgMmKDt0s4r7RakJ/Md7+iu91J+F29ugl0A7tWzcMtspZzlF2Q6dEmck
xaJ8cYkLbC3hwAEKVFbZ36xi45k8ti6G/ZfSdGig8Z1/hOAL307dEe39n5nWgc3HjMs6cPR0Na1v
HBYAmoi9PTol5HC80VBBUuMnz0L5klSxIYTJRFOEo6RCzOd/IjyERLwLD04tjpeV9yhyySHPImbK
atEEC2qxNyqszpsRG5MyjaXy7orXb1UMvdWUYouKh7Qs9AQYEjXxkkdEdHaCpEdT0LnAqt3hPrjT
gucdpW1VxRPEqTL96Xekm1En/KwdLDwmIcfbdrf2aWZb63T2g/tqS3eclB4i2Eqm9V/Qd9mXjNKD
dlav0EOj/OnzHOpdTM26RvnubQ2Kd2gL9Fqwos3lX3yDtL+m5xBco7jB5UZWuRPNcWJCgnBA5zVd
CqxjHok2A3XAZQ38/hPODO62UTEEbQ8jVQwjm+VhBsyaB1M+1SjLvPLrgRr0QMqCXxnsKyeLJOQZ
aNAruw7lVnkAR+D7gljy5nxrGxhLWmkrkeSQO+aER65ihw41kQIC0KPfPZ7t1I77W5bCRhYv9gXc
J9C6KV3aOZA3pPGszNGDUZRw55NjBp54XwUvof4cXqdLKQoWwR34OvBSo971PF3HbxXvJ4MWf0wb
NZVAodYKm6BTV0VdLeYRegPgMkwTWyGuBUDhwQlQcAAv0Y9Zdx9wraHe4xqP8/2FOIcbZwpDeXjv
69OVF575dIFm71EPJb0yjNLzNdBharnpkLmrt/LxQXbO1J4zeInJlUMsvjhskiS2QS9deyikLOCe
i93SooXN2yDnWm1EZqTAO66ukCHeaUW+/wG+vVpwxf5pzH5+Dz1Us37EMDC88fEZeKOO3z6qSut6
DDLIzVAeDDkbrnAmeC2uev4RR5NglmJ7TTTx9q3jO5D7i0aUlI82t441s5e5/KpL7G6LoiryJXwS
qKlD70fL121JLKxXx/2s0anJ2OIBhPe2iwUsfo4OEN9XyoWhS1tr7BAM1LLb/Xr7gyAed2Yzx/9O
cybBOaSo1Qk3uDGVYWWE09ovVTTuuHJDlfQzQHmhiWOXkwkdj93um8bnKvUSHEA5PMqegLOpYN3f
Rgugu1mbX+KOgC00xlwFEa0dBqiXbbE7hC3LAbsedQqxpsaPE2Tpbq7vRg/wJ9ydKzxDQQ4YCap8
jrlYg1/HlJNF4qyVJCicvCnBawGTokCXYOmVpXh8SbtUn+sCQllQL50EJbl1tWrHf+/m5kcERrXE
k/bxm9/r8uWVzwa6FZWO/lQA9WoA3Q/6C0GS5OwSrH3Q7xpBJkOpimwJGHCg5eVnKe1B6mbc4isX
xBkEBtghDcNrAn4pknLR8Qgz1uoI68BdqsbTFLNTjEXjo0E1jcWy1mRKHNSj4ehttUEAaUhtv5Tr
c9U8JxlcYW9M3EQmuI13mHM6c5tJ7wFkyARZ3RGXmwBEsNo7WqwMQgj30PbynGIwy2RdB34Sk+0A
+bSQuPWZAQVe67/4NoRR4NvqDZHr+WVlqrsS/+5car461RP28ofT6saB9I/JsKh8g32G8iXvzR5u
y6cB/2EH10uwikmxk4JFoTKywrzTcK8wXrnD4GZdWbyLxeMcPL4hCJSA/Lp5lm7vfreK4PVxFPeU
QRi3PteBluWdTfApXEepm94bJAokSKoe/u+dJ637/blqmGUmNXjtggTToIRe39kJflXfiN3GYfLB
gJQsmZYahx4Two2k4rf/6i1YCn5e81hWbZrjf8Zk/vVOM/1Z6gomy7ObwRD8QZ5QtqK9Bfftywqu
QWf6GfJYqUfBJZGorENJEdlc1sZ76l4MJ71C+f1DsTC0ooZgnLINdehaZ7Psx5IPIyOKOu+5vuRY
vmnE5fKECKpDcovoAeNR16p8Y3AO0le1Ts4MpJjmyyDAJPl+M9McGZbAQURx/G31nqNpHJFGHNIs
dfrI36mPNM88058IJvLnPHGVpxLqyRUzPWVm5dwYHi+Wl0JRZY3VvJAT/MrLALzzaa7UenhjhVwW
DH3bVL1F8fUTyXpRbS4CrE2V6Ea3pJ8p0cRVPb3L1lqs84hqP/wJ6pFlQ7KLaaPLEmHPBUtDP7hC
uTZ9bW+F5X+PiFo5HgHc1pR5krbFT6LPviBgS9EzP2YocZLd/Co8EKjpspFLeMxcg2AVORi80Opp
PDPAEFPwTEkdREYHFvt86GBHx+8M8C1winIPp4UeJi02/Gc7qnMEJLk3rVrD3rd16flIJlBKx4qp
FnCVQrAMmMgpxxichgLHjDfTTu0AF4aWkD/rgm9PfYmOyyiSoKVxC+RreuRYdnIQfPQUT3qgUQFs
GQ7gLMEZAjwB5HtPorKPEMIHEGAIwfWQhh5YCQZM54jhRhR1WMZqNwdmSn2xQ84gg8xn5fpYKOsm
Pzdt/w8xYDM6LQgJl/sUiDD4ScDFcVH8J3R6M7wAxrazPdloZ5yQ1atVa8JHp74EKuTW6+6XbTm0
T75F4A/Bght7ddARZiK/MCADEI1QZL8tczSt5P+2zUTxZAPWMB7X9xZfgOvNrnlnjNN52Q03ByWG
QWOJiGhNTeC8QrHYUmeLPCf1HWENrxO8pte9OtJg8rajNc/BrSv8uLBba9HC7L8UraQ3EerBiFjm
CFahu9DD+I015ctVdg/qyq9yymEy0G4eUHuU90YBBTgLMqaLtOYqDxGn7xpPosfPRVV6BdkSGGDY
TLYlRj/X48uttoI956gvtcLVKESMVroRha1O8l12dOOZ8kmFybAS7YgiA1htearLVhPKc1s+OoPe
O5MK1TVJwBF8Egj2e1gCJyHw+iJ24/WFopOJjnjMSPx4wRjYTonVWEZJ/w8KwLp9VXBR0vTBI+AC
+bNpA3B2BlHpjiGbMOq2ruoG5qvKoAR7l3s8WuZk+NugpPPCYBKjtWw1ZTUx2uhD4sQFCnQDCe12
quzZItjdm1s40BJjwH6/W79FOJTrCU8Lfbqji9nRs2haL2CFq0TwqREZqP2NC0Tkn15QsSWHXc+c
SxDxFUTEV6e1fFjOtvd7hdjaxt+u5Wd3Puql44+jDjMIKzD9KoPPwsrS4aK69+wLTusu2wHdxtkj
6wtu4PU8yETXFQ3Zx2EDnJabHMOpmGcVn4PI6vga8uurp/uVs6DxtEq/dZ9YdIH9Y7heFuL4Ror3
GmdDMwIvwx8f3xbz8RbDez4WtK0lQzPY0qi6kW09K+TNEJSvDUa8d6rLKqrXD2ZzkT8O8ir9YHus
N5JfY1Aia4lu8bQ5tbwl98ksU9kEHUnWYBPBx9jtHH5xezEOwpSmDJtb7OFaVGHzU8FkxrWQ3Bge
0fuEzEJi4DZKU/yfsrZT2naxeLrGZzXUkBwNCquCAAa5qaub23buKhuJM1kJoObTVVtUFhdcg9Pd
sKCKBAYBXcfe8oUwtPm8gEOhVSU+MWrkSDub4MEyV34gg1aLj4r+jldm1CrI+AQDWfKKTixeTw7I
Yni3mATgSrzWVMJpV1EJtJXcttDCNXn3QrRVmS0vNqHMenmHCFVPMEAralyqjQjtIuZWMtQvKkMQ
MVVqDGlxswhW2FF9kHGG76UkFhK7aqbR/gnAydigWeJS0eaKJ1HG0ySfFYRHpsa2A99GDmNpC4gS
VnE8YQMqriSIdAuhXctDNxuq7P56XYsCVrFYOyZRWgAmJ8TNJgAZM/R+QMuwpeFflkUVWq6cMPj6
a+NWDrAzicESA0HLnRU+/tdHtuUmgfgXeQ06ekoZiLYXXU/CTFqBg2k3mSfFoV5vVqgEKxFUS5Vm
RJ4hqP8VJ7v65C5+QLF4y85iJtAVcrRAeFhtDBsFz41e5WEBcRZGwFmqbsZwpJBZaSQve7mU1xqN
cROQDROk+568mZJo4VIBY6BQ2sF8BA4lWYhH6Bdzcfd2/vQN1X1po66GaZKcokQpi/OnjBUkUHwO
q3MeMppiH9+HnleRbTV7WCHXtEb9Z/VrrPzKdXIkOFN9HLlQt/uM/Tkf0Nqozf+gQ5E+0mrxWTYD
ODcwMSGClm+q/wszfKaaOvsEtDOBS3vAm0Nnrqmb+/E4cIHfVyIvVfc9J8Cai7PCAnnuqQ3Qv0ed
blcChRi8Vm8G2Y+xcIFAWEi7tEulvYxWzNflJ+YN89lMDKEIwo4uQ1vNrtnW5qbiovl4/2+NOPp7
/0xYK2JbtZmmqjSJ1MFtaer8PeOoTal6ifLRW/Ld8vrJs3jCbCCfzGPBLpDfEPp1xAb6hkBVFXcl
Bw8BwwdWSL2dV8j7dh8f9lnBWZWqiT6p6TMu/ipIqB3m1QitDmLiKd4ZKGxJfQGqCGJDsVFyBgaG
b4nuCRqCddnYmvGdqW3mLQh4IUfbfWST9S8Q3vMCybQKyuraCuyWr//6+7fU1mTrUedldL6m/iii
mDTIsiN3IV2BsXESSLliQcYiUyFvVoe1Y2TBQbMie/3yGSCGNolPLpPonKbDRiWQfoTcIVeoBzsg
Okajj2bz2OG+rtsJT3UvjE7SBtq1Q8vKkE1q6V8ITU4Boa4XJpm3+g0ACHXnfocYrEgHrCgMNV1W
dhp9dAhkI8NFXTOInPlp+yU0qNk2Pi4p4PlfFlIVJAeEzxCa6WNqKdmdg57sYT5f2c6J1EWttJLg
OXlpSNPZDLtV2/4P+VHEhwPIMVJJP4oT3BCAiaK06dJdr4Wff5Eb4ukk8wZ9uleZCBKI7fKWJ9jS
ZEAOGDS5yEv/9sp+PDC6rQhHKP6g4Q7iAvun09dWQGEvLOT7oE2vu/dm/ia0P2AK/VJw/gBwnY41
F8LguHepb7XzrhOqvoQOE/mztn7viB4GD8glsKjrM1of62A8hmPoEwauDIHm5Z+42bTtC274NWZM
1YY014kSr+O64XEN73LbmhMbwTZvbq39UXVY1eYwDPo98f7W0olVj6a/qZ0/BPXND2uef2FMZfR6
FDDgRRAP8mnq1///9ZryE1QiBAFaA7Ms2rzz1Mccxi1P9Y38skys9NV8sl8byhwCuWQiTFSOJO81
xybKfg4qw7s6LQgvgTgfJRNbFiIUBj7/zOCCTdmn53cqcpsfuhk3WNXKKWQIthSRs7wnrKrKmr1/
NIeZRDdTF/ikRXzQocw8Zb6HoXfUKFdApviXYdrJTlt4D7V7tVWNYK+kh2dsJMrUvQe8gDNnux+C
tr3jxHuqEhUZsKAk/Vk8kniGeuLFsqViTAqTcW9UHesu9Xc+9+5NHUiCN++W39ymm4TDBRR7MOZc
BiMY4h0lhQf81avpv8+pbuFaInGMnHYZavIFo0oF2qAWustmZ3zKwkMWeHSyYM9SjKLB39HUjbOs
CNcPm8gaGMy1xlVdvUi8S84sxx2IEXf7rI5noZjHHJX1S3wMmjuM3sSJdnpsOQxUlNwcyrGDyMBj
wARlRY84biK6sVZndm2P6rcyqFhLlr5zwqmFuTNB1voAQNmVlRc7ktZ9hnecrctP24+vnCJwUqP+
Cv03nkLLryk7OmDD/UIOJIe6+TOtIvqqyIpYtGZAfiRZQSHuswiLS4FJX552lmW2HsOgFT5dfw/I
JKjM/LGzhQk53P7LqH0taZ8PwsIozWld0IS0hzuSxFkvyBPnoTRNmj6uwxM9hYZKSJ/ZCZOBAhDF
YOkJNl6BqWSIpThTk+s37jhVlw7m47CRYom4uyFf0TJmL6eSrckS6IE1ifh4AGz7vXmbDaZAExL5
q9jR9mudn2NYmtjFjBK4WJekOZUfG5OyBOnksDJf8ypQkPXJvbUiSlIsz9L8kAPP39QIkyBwWHeW
NUjuVNlZLpX5PbP2UI0qQH3UmAtdIPnVUghf1i31q8ZTDv7pylIrvnjS28IUkKC1AxGK731RoS45
hPxTPP6c5Ydsoo/Vrp9smKosALioA/4+hfMu4kpWhxP3uUZBp1A4nYml3JrfKxnj1CBroi0gnJrM
ty+LYF5AcFytQGNEbZg0j9vzOPnQYVlmqAtYLkeiNfpgZpRIH32gGxBvpWCmpxxs2Uy9KmVYHzJl
mge/+GTcN5GapvPzTPpx8xG8uSaCeXnQLfpkCtZQ/gqXlntT5i/rjPy2U6l2Pk9r5RoY90ArwYER
K84E/iGbjlrFdQdoqLr1mdth2ez4hbKzMoyma3kP2hLBe5XhNxAHHAm9FPLV6aJHRw3QV8DG0q5W
ASdrK7SXjm6jnK+OyXzZHYnEuE640rHkKbHTnVYa1tbr6RfJY1KI++CwBxk0dCsovRqi1706BE17
VHYnQYCmIuo4PRlZAagpXv/65IL+ZigyHtiV3eHAdkBKNxetq5scws1w3PKwll8ubf6jt61iqRYX
g6wygubhryFjVj4ESm9YZM6VyBVyRbG56M+MmxC2koVEK/2G39LuQdUfCeiKUHtuadQZUIr8CZeQ
EsLXeXVCyZR8N1IMcEIQa6zZK/dvCnp3U2zWjiaUckMq3UBSAFylm6Mv93kNlQT0Rmtx72gkVheH
FmxT8m0+VCbDeCXXk+So3btVWz7JS3hR2aesVlonMopsKRGKlKclTn5NsdVsUZtL0KiTJhOgOyBW
7ScOCBGFIjOnyDGSmSpn6VrOIKpMlsOM9Zie6uhvfmV44S0Q/bck8XwmKo8k5i7Gq4NldxVogOih
wtICpGzKc1718Nl+U7xONLqTJD3isPkRUA3ECI1hdmEAHeXT6fJymrtfWZy5zLs1HHpRzoEO1Buf
HIrLge6kMxOE1sy9R96GrzAqPSm7Um1Ez75XJc1U27CwRQ9563BDuTS5CJhjV36N5DG+6PP0NbM4
HNiaYVppMrRxphztouJfxASygMQpaO+UFE9g7Lmfrflyiv/GtuSAh4UpfxlU9Qah5icjTTCzwHpB
dSYgasbYhNKVxqYS6fVz6BX4EoBUf5lXlm5zOXihw9W3PvK8YP63qRRKqapjPqzV+aK7HT5mnMTz
uMU+2HGO3O2HbGqNTkpAnEuT6B7Ht49KOi7DXv+13ZcpGz2Kl0NrE/qmtaXPtQlqMhfSFTqrOemc
nnupiMdofyg7JxEFXmYftbdnJVGmwNhEKwIO4dnTHQI3h1BubQID3ViPRE4gZ8HmPURp1V4SUjdq
AcD2zvOqTj1Q2eRHGGCKjA1i6y6fqHu9m7Hygv8nZSJDCfmgIqo4WePDdRhdPKwhD6NED8jQaxeQ
fl7CRfMQGYs34PQEaT23+U6I2VUzhU+4DGsLlnSatqy6Wxo4xBee3tnTg0yRMGwudk++q7icbB+0
+bC7cDkBVl5AFcgM5N/oiaFRWtMwssNoI8e6dVr5CplDoBLoi51xK9/3+LvxQiaNkTy30fwWDsxW
702v3rh9uPfbFD/Sh00fbMB7fFpSxm0ZyVPiZOTABwrx7e69A7hyL8gTrDucV/8MZdttANQhehYi
1dq9yAID/BmEbO7uXq6TG7dg09wtGKtAs1RcEytfh+hACEOdhD+dnCaVz2x/wvS6ju972+GLKEkh
CZwUcvpWNH2Ymrs7olPzGZfzO14xzNQTqJf3P3OBhNM0bmrOszWmJFjoNlTl1ktqoHO5GLd61GgC
V8oKDjuRdzFuoUF8aUu26j38yJMsFsk/qD9foDnhQD81/1r4R+bxCh93h+2ZiDAw2U1BdzeBNHcc
S/GGgxGDseyG/ZWRxwLHAb6v1PFYcXNrhB/ngP2VI0PjW4ehpokhjD6dHI2xGmX+3J7qH3q5KFGg
4FyeffF2LEoo0c3tP6njh0wed2+3tvi0H4sNEMdqhW+1vS6KWEUjb+6rZT6+wiK2pExmFb/kolCv
ycR2ImL7wc9vwxYl6GvfPy6J8VAlclgp3bHjjvNrSN45ODK41kIXvFQQQVylOHQT0cRdRPOmbGt4
RQaPkZJ5wVGrzXvexXnaENNeOUeMqCjL5QqnoY6+mFcCf4I7/FeaKdagUYmXlDU4M1W72cBlA4T7
ocs2hDcItv3kjIcMjRt3oZyvES2ORh2LfspFtaxjTmFtBYx/iWwWIt5pNhW/u0jwRnhrO6EOI8Nj
ZsY9S9djDnT1j9UR2vytnliEFV6usCgZeqRTuRmsFSD40dpzzlxnpf9Q2OZ8Mu4IAOCy2rYKVhR9
M/VIzC3I3HW9h7FTnvLoRIUyGhKnLBcoaHLjAPQxiYW7+gQlUWLM3tcl18hilI+L08WVlfhMVwQB
G1iM3boJyU9zAL8ZG2Vw8pnHEZ6No8ukUWdNvA6qepPjR7M6qXNrg/qDOyocgg9Yj2fxdmHFFNEz
tsdAqdAUSYjuzFSDH6XCd4JL7tKXXptvtUAziDUROVknZGyJVFou0LmktjSgM1m6UkgOwXxeOM/x
XS0FSeJckGXjzAJH0lrOkK3aX9KLhbxuRO3GJQBTpLV0kgGv3VNoijJRlEdaZ+ihekt4G3fv55uT
/Xm4IncXPkYXINMypWzcJik5VmwhJHodxaoAs3pFhpsI1uz0Xs8yZGTBfpzlCTti942QQd9IBUH8
DmA+ZTyhvd/ACye4CPv01saXPcX2sCtPw+hhtjjESS7cUL1D778Zqb6SW7deqfCzMD6GFX2gidFd
LmeJ3CyVMxIM/YJwhQpIn1fG/4F0yfIyW+vfMvg4oeCfPla4Rn0CrCj3MnW1aQCXhAr8Uy5k8Mc0
yhB0RmJaZgTmOtDVb19jO0uz8LZWAsbt2AFm+enkspj9/7H6nzX8ZPRzoP4r5cIOTBEACQqFm62H
rx2b5bgfMKIAtnqRXk4tqZrte8Q1+8iJBhWOKo1R8mJHxDnLD7pfST3INbSJfCrPlPugZFyh04dx
Ngw//7bXAGTGtVuReoquTh7HP12zfM6+HUWGKa9qCA8tUZMhmAA7r1uC9U2NzDetyOwBlRK8K22u
kK5gDMP9WOaNauNIAZOob63oOFVopNA1gToO3NPyoHLNC3QYejhqpnhFpOdUybrWPkVM3Khfdh3f
hUtNMr294sMF+Un/sxW8SqkOXm1jq2pkKzpznPS+YEiqlihVQyxnaZboZtqRtYrzL6gaxHJuXOzJ
UlqiZrHElOCMRDuFGg7B6l4sqOje5sL+/Ov768zlWdXFMmRAay94Y5fsMyITNQt9gEe0DOtnxXjR
eCvWzUKyq5t8MgQ5T0k85LpPI/Inc0Hk2fNVxbViOFRIwIKtkLZ50q62DsauOi2QRcawJ+p108vx
CDFbN2H7+5hCMaSsvIS66eTrM+4oE/5ngBdsDzg768e6WvK5+N0GmAhIxMoUEKLNokbqZKVu0iL1
GEYazXtLx3u7TEI0j50qXn9615lX66o12t4ORSNfQnXWC3nIHo9BayLXUXeVI09ezCJIIDIljHnx
4A7XUAJBbo3wcRjI7X8L/aJxBSxpvmGHaQYU5CgHLXEYV02G3OdmY+xUqpLMWo+FSJ0bfqAggP0x
FBJfsr8e/4yj8eRoowdBhZdqgEr+XaQdAhQ/jTh5MKHLiCaPJjISmh4vAwGTr9DeFory+Udtyr6i
vpyvanRAG+uJvK4IpXY7REF2hDg/RKwbdtkd5DE5vqoAJScG07Hw7wy+S/l7PxGKYa5AQZDvQ1wH
Ae7CDAQcIkkHRVJ5Qdnj97v3bJqPFVyF0YnkxjW7JmiVPdkalTnUrvVuNKBdNYms3SA29u0xiLbh
wYm/xwcgTioGri3TrBUm1+p3U9B0u4V/Sei2HbJBQ/amyO5YY7UCOHtt9uxWVAKOBLjbTROvT2AT
SXZjRPdacu+QPkV6RDtjbNrN6SdLXB+Kkv0I1SjBNz32LH9KRpO60wAud6r3eUPjq+zCUZkqRZVW
sb7yWuzI7cW0LOjboqygCvetN4LD1CLKv22cj3pt2pfB8Y/qVlcRy+DluAsCaXDsvF0WwyN1pVqh
VyIHSDxBJYxtdFZswEB4RfUkygLhUbqS0yijFPTEqhSrENfJPXuzO03Ps2PKj//S5BPHTU6yRPuV
GWGe0d6u+ClnBFvxFB51OeCrNhbCTg+iftN6K+QV+u7XTXRTOBaVriC2eqZCljNs2TwtdTdo+RZY
5JBubXvlxbMafNhO8lTjgeNwOvoz2kpJDITMhGVDT3GtGv9QMLJEw6PBYj9aS1NVl4rfq5c4Aotr
931EsHx8Jq4QS8JGHRwXhDvaVyhS4f2irSFWnoum7U04XK+app2r+zXXHbs1LkjlYuc8OsbwBZOz
2+6Hf3v9bo7ltOF9sSdZjuBeMirViacp0Jr+uVBhdu8eqc4N8IfDf3VVqq9lxk4RuRAKFFtAQFtr
17aGnhDe8oeQu1BQMwBlXSFyuuEzApAZt9jf+l4DsFSwHvc3VVPxmvUqdMFnWA/Z2ueRWAlMIzMR
8LMRjAN5MkQt8QQ2+6/I3oIYYwC6lm/NUXOZ8bKsvfgNkolqs3Lqz+CA2YSLyPx2UPskmPD47QGg
icFUEXVKXIRIavFRoN8h5s6OaIgI0JV7ySg+BVd+lphyaVWeLT5IhDJQMl7XXOFLVvS+Fgg+/1rN
QIRqTrXUyBWpmF+qnS0EuBYwdWjLx2m/AAPRrtm94grYwzTx+SSAK2bYRgMOy1F2ld+HloTaMUjN
PwvqIN3QNUFMt/2T1hBUSV/FBXewWJ/3IldsdCnUDpK11KQ/5dqQ3yjZ3YQ9+6nh56Dn6P5BSqRr
5WTtCrcXOw6xqoqDB/DkE9Z0BXJCCnn2BGSU5TS4IwZ3ry2OFimL50MPsP9oKlWsOIAdEX0gFoD/
akfns1Hv7V3nFNnHlTJhnfZMlSJEh8YQYmX/WpXCTLNqxg5KscCx1opm00CAOW2S+aM7sWOx/2aO
smpS4+sLAn5/sSijT73haLDRbSO/QzhwOvXxt2xrzsboVZtrVKAxsI2z/0Oz9L/weDGEZUAAtkb/
vxZ+vzDcbpLSpVsH1isOyjermOGN3v8n2f+igLtzxdsShOSEpHqq6NKUqyWGRBO/qU9yK52jMlqk
r+L8yeA9KgH3IH0fb+B/Fy5QNlF3UmZSFETXzKflj7TsXrk8rGAwIL/Sm1FY0TLXJFoXdJdrdt1V
we2UWe7VX7slstLj9VSNmUgjLtJWGdw8kkmVvW/5i55AIXMGy+2ERQxAR0WDIjDIXwTXESg952gR
ApkV7xaUvdExRtQDj2LJnCWQgR8WJ5P5hYCU5VtN/dkF9v+4oHrxK9Dc5IhbsUmWwqNVs4cktZqZ
FcunguvN6c8S7XlxNctJOPf//Sqpa6SfAmYVbMxEt5prQHP/0EMTDMlL2mn4nmBfzglllYXYHAFm
TkDDGgwsFuJJzf/TCHpIq0iMTIdPo0oC88NB2Xhm/gBXGUacCeFLPfwdVqDU1vyPoW1DE6nX7MLX
+vuJ5gbJI7wk0HzsAAziOBEr/j4DsV6OQamxxkK2RuSc8+GrB8LW5JsBFwxLj7tQcjHK6GU8MJ0x
g0NkbHNNQHrgXO0iVRQzX0BgTZpUePJ3nIH9sQ+MWndfgbao9dQ9QlKfYYD/maDjlm3lrsdZK5iA
uQjVDEjF9zt80+MampoBeCjM32Y7eYOQotvJOL2Q15ly/Sb0KqWb6bUb8C9H+s9XuXh8Qg6Wa0l/
rgqDOFCEzQwGM+wTctnJP3s1oBdzhT/NLSwN++tr0e2TEcfD+9sB7JcC6mNN9vuFoqtpIjYwwB2s
Zlj/uNs8Ykjl71Qw176xBGN8MEnsTb+6/A9iQmWHKx0lknoKwiLwaEXL0mlDm+GDxIlhdGGoka4K
CRjR+1tGsuGw4rIgLuP55mCkvc73UwSYIBdNGtm0y6gTa9gWLV0HlWNC6QO5UrC9ozhlihVFOCfJ
LPVIjFtRimUdV3T5BRuzum7GVqAc1aD33/Ci2kBMYm918TBcLBYsVwNYo7UUJ55zVAq1Mr8QjBu1
tvcA0MrQf3tOE7L2BtCTJoRToaTjBHhe1aotgPJ8sLD0Xl/jNSs3eYyrijACy81SZTkzZuWaaujC
6o1eUsziLPrtDMLgdLISvK5UQllBJiKOsw2g/QwXeGLWynylqjAvH9uUMYl2+DfGj4U4B7v82Gvq
iwjy5Eukl15ovhLqi7FzDxeQU38f/yRgiME01adnG/uPTU03sZjk22xstop5ubyNL+zwwLVI/1cM
aTBXphAMdk8wFeFqioy8LtmlRiut/wOzQzEY2deX1NqhlOCqyfWC5iBym2e8YPvkICbafNcPfhcN
Nsvh5JG5jWGzEnSNuA82fh3LOPi/G06q044crKCRaXzLi7kqblm8WJCYs7gXEPMtiARrI7iAWjak
/qBLmOz5AUD2sNAFtiPbAII8iuyr+GQgo9cNzxfowPCVRDM2UBEE7eS+KLqlIbx5ixfOOVpUaA/H
LOLVNJlNa55vYqKDUhEm9tbmOekG6vaHKUG8hlZQj0k1JvYnXvA/Po3zrO9aMVMAcjak/ZSaItl1
2OpLg2Zmq9iDcRHXjdqoB1tvM//KEpEi8n22mOOTzz5xjPyu9pIY5qt3h7YAxHqRp1y1Rkgnyoh0
L/d4QZmfcbg41e9Boxh5rlMEZJmKrBZ5mAuZxCSJpJZqnyYjdhw+5puKjy09xSD19BGn2jJs3K0y
1kcjBWw77PQh2HCrMKSL3gemCSechE/aYUFQqakV0jLlywSVDt291n5GCGg5OOTBUCbO75dAyuXB
WSU5R5JNtUJvod5l7H9RtA4kZyKgZCHQbtSVmhBCE0J71UnzK1zvTCvUJBqg3H8ZGRHHkHcs0XZN
T/S3Xd8wM+8d3IYaicVbN9FDGztXnxZrO7oSm88vaJAttiVSUjDiOwRM8YkIQNPj1nIKBETrxBll
qaWCG6gkEMvzdNz+foH0mZHNnSXR/abpqTJHTxpkHQpBtXgS8KiqHkiJVRjcXVxCHhJBgcrj/g+G
qWpFsHaJkOVgpHlXJog5u044NYNX3kaJB/cGaFBPuSMOvyazUwqfO7DqA8LpaAkZ50B1gl36PoDB
8N0KPCWJ0wO++eDf8Evl2tf+VjBUbN8vLip00uo7EhRLIKuazrR3Vj1vAeTs1V38Fw+5VqZ7Q8dU
iDyl+TWI/pQpt+NbDOuua/JZWMMQKRstP4jl+e/1wuC0Hr5mbCJtLUCg8YhdxuD3bzHTLG0qWgOg
j1xZb2GOfGtgruNkQcAibSwXIdFXyU2C1DlzcdIu67bgH1pZnjsuHrBiop74Yv5A2LJqGcYrN3nI
gviJ28HgLNqN4QrhiydF31rC96/LpNtCz58721pCiW5ryD712lvKO8FXb5SbBmwHyCEss45IBPMy
rsgvq7oTFLAhABtm6A1wgGci/e5xz+3w1lfXt8F/OUu2nrgp7JFLr43qy2VIzBagw7iX1SpFZej/
JS0E2+2IST4ZiGRYk182UkAzet9UjwsIWTYEBCnInF0IthtrgdJRunW4y8yI9kLZeTLAOCAUzH0y
wBntYGWJLJlRtq3RrrGO8CzGt7wS2ARlo5GTUs2slBm9f+SMxmoDb/p4BG+p06XPN9LbYPQ+PROs
F3R9g1ZTYN29wlSDUyD3x042LK5HMyRwyJDtvJ0eb6KIhHTXrmi0ex7l5BvCt/HyTAkSYgh4/eM7
76QGsn3hSWDPvYOnm+Tz2G1xY5qheUdSaurE1x0yKPvnOn28Gxoc6Tiz7wr9cRGm93Qz72xhR+kw
fByMgbOCKIxJ8l1JPrSCMNQ173ROyLNWEzF6SV15VzFds8x5JrYuy7yDew6U4Pi0ttNytzC6SsTh
C42dzPCZYg99SdiyZSXIAZx3h7xyPmtRsA2Tp56yCPllzAR0fTepkRUlGei28x4Kaagvxey/ss/D
ULZ0M70Wix5onGafBZSZ3Rsp3CxCgINeYtzK501pEWTv7bAsbhyw5X+bhUjdDRGH2BhbCLc2EUqG
InWeI0d70PzEvRQDXNzOEIPR8NeIePC6CRo+2oKhxjVzP2+MvQ8lwQC3WzptsGv4nfBUSTROIx3M
OkkTkHWLDPSPosrHbEvJtpO22zUw/J9TzlEbVy0jTYEWKAWUFEKzz9fxd9A7WkCgzTNPmB10j+fU
6IVcD2BIQdxuJqUTL6boPsFYMOlYpEr39IUsWu/vL3MstYhXCoB10urqyZAdERMOIxtFUa+ASH7A
Lx3AhCY4s16K8rMVoS8vE/iZx2rwe1KvDZcMeuHh1DFgZf2HuqUkbXwVbvwYFF6i45fr5DAduOwv
9csfrQfhuie0QdcPmNPg77UVEraP7H1GwqpAPaFGUpRUtT49sZZ80ZlRmsfIysrA5tX3saKx4ZZb
i9zkh7icCV7hlrKAtvVqZJVCMy7NgzrbwgY52seGI+GYDsU+RZHPZUOoQmkTQ5bhxqKc5tgzw3Kk
WcgrMcejr0ytL82zdjcEEGxdzv2DeTb+4yIK/vNQk1eG201r1hYzEvJOrVpH9LXz+Vxg+zZkU9CR
m3hexIH+MCIuuPm7ZIfrZG7u0ORPJ3KUzVItuTjp/gOiUzSsb8pAFy9bDcx3tNqq0U6oSkqv2WVV
A2y2YFV/6BMeFkQuO7h51LconXz2qbYL3j68haq6ZZ3/n6Y9eDdhOJ1DJy3nbo/t0QqbHhaEhZZp
j56O5Dso5z6VwKsKssyVZ6joTsWNO4qndYnzhZ1jgjqGwuy4BuuEQ/pt4CGbOTgo/rDD55XlYUEY
FHn54f6QEulHSLbydQmpa0TmzX0gmFOxd0SQssiDJUnMVZy1howa5+GwZav4dI25VZqOQYfEVp9L
zXp4G/tUGsbeUCGXisHNMwlgE2nWgx/tYKm5HvTerd0M0fTmIDbbrOEa0UoYvFEVL1j+7U7M+Ded
h7NVYBwJx+5j4k7knCrS3DIlD76+f347W31NxA9LmUESfQBYPXVwV18XxVdeVaIHdUUR2+vKMXyL
Utfj+bMomGgr2M74Uhowouq9i9VP8XB8XA82Vr2CcCfMkm1cSvfRkX4rUc+nW/JN7paqY8Tm8PQ5
2KTsrwLMnnUW1+8n0rfLQA1xl3gwXhDzHfW5dmcLiCinTi71aIkADHGkL4XHRMC/kSURzPpGAj03
bxSNR8sSDYskYj26NJVcy9vLsta0by0vpBq17ah8LGfcZ0zASz5T9Z1iJfxtTw0JEV4Wi3RCJkZf
QwSIc8GcdMxkBmQVEj23nc6bV6J2+nVUlJ4ekMWwgTNzTgPki9YDHRnXMka3KE07PGeCDjDN4VF4
3rZQb3cfQfA+H1wcutTvMz5aE4VQHhX/riV1Egly0HYgYnaMSUTAsj5RACoWTBNtCsA2lZoQ4J9M
MlbljUMBpwEpovYDW4bfUzJU6W0BXskhV1nr6xJCMh1Sz2HHs2Do+b4iDpzdS47iHHNiJvrUSj+w
yDubeu5Nd1qYiqMtBMQxZ3VagoUpWLia64XlFtAwD54itZKeiL050WHBFOSSavvB6qCfnPM5mHEQ
DNF0+Y5cDt3OEHoVAvUE3F67fMiItIS5NOVNLueKUSNL+qT0V6lwdCqEVwxqdIVGe8mEbt2TZ+NW
o0GMyEFPvVtIZs/vUilrC/++kHw7rTebIePQl1E38Ogwt9XjXUSGL+YdsNiEl+AG9KW6u7A8C/yT
+9k/lmF+VNbZkwcSuMnpM7g2ovf8rk9jsxidYS3kagHiv0Zmd+vtd7QP9JaWNuBcVOL2FqSj8H1/
lWUOjGB5EUoYIr4il0AJRaVVRrjH+XlMOc1lgttjm3CnsHx79gGrWLDT7qkCh8rnBVv7pzJO/LeV
8g+kBagtnU+oCRi3lPCG3hqMnB3CDfJDw5naFMJE3MhBMN768Qul0fKfUtMMcHk2t0hSx/Oc/7cH
P9j5ujUorpOFUefhTTa+RKT+86rbTb3uBoUAA2GJeJdJ4jDRAxKfVHNCB1KoRkiupKjoSgSP8k/x
lJjeykrhO+y5nv2INM4fflo0PI9fCHpQRzyR1Ou46MeYCOgXF0sOMIBeaKPI6lIyf1LCeQnis47y
U85gYRqFO+D1XfjiC0uCMddGoGSxijmtpbrtQor5zHSIws4m7UJKx7gTZAP9Q2CyKjwTeY/zCGwQ
G74/OVuSYrqdtTlrPXBlOQpE/HOZ/jwASKxXUkva5rPUeVws+ZTQ0frUEIs1B1ReLNlYWBng2J5B
0UKMk+/dZzkzNQTWxU8L7bgwvB0eXriHZDj8dpXTrLCLISrUN+IRTZ+W5V8NVwe1OOKYiJIw8/t+
p7q87js+C0UDR+DGhlJW6rEMKLts6ULL0t+Rd4Fwv0FYJKu/i1hCOoP+0t18hyJihZfa07fMpeUQ
GTtDgi4PbBDs8cieDJ8OK5zOhyq9/5+UHvcDtzOZ2yLA+3Y+T+TH2UJ5f6XYVciYVin1jBtWkrw4
KHCZi+LKxQBlhHJZMpvoBFTigrQAOEH90K3TtXnsvhvsQVIk/gIfc/J+x/pfNZ9r3TQWc3opiwI1
+JWk6UWAnauIDjihFdv/SkDuWR9BuV4hCetdglYAtWg/8nksbmNwbnoGg2mOMoVobLuC8FPBHayK
2KK0BSQvfqq0uVYA/mOUbqVlL2GwvKHqN+ELlh1o1n6W+EYUTuH3r/+3UE8uzjUVVXorWvp4H045
qYN1IsJskgHODUlhWdu18QckWdJmYH9QoQtblyoUSbTqOxt23e/nggL+JWTdKnXkPRb0UtBm0QYL
3Lm1i03XnjXO/FLs/wylfEtkLUQRdDiMdLrrGCR+6m4ngXkLbPfOhjgzBb4tk3Q7aS9S0N83rAmu
ssz54l3qvoQCYEjq8WNAeuDzR1jlVgV/qJf0sswxfUrIqubLpwVxbKm99RS8joe58f9qVoyIQxpw
BkRtkuzgo2hBHYDbvKStH/sAfW8GRDgpxghDb8N/O1FTSo1jI74JhNiBE40HRf7r0SjW00cilXdv
MTRBlo1ZHUZzI39ZpDERrdlR0tIjk0ebsfwcVVHYhye3DVm2mywkdT8/vLIL1OfLZYbc1y+w5ajd
yeNDnYZIEEv44Ei8zUckeP4y5ubt2GVmPWRK+3sSAnFFFTfY0V23ahYg1lzV2HjlWtVL/UuxaBLt
H5Eiz0RM5eQ5YzCd98rP3CftloOkj1/QdMA1vKKE+8Qxuln7ufTz0X0l2cx6epiH4Pv/r31n+FVt
q0BZCm/nSmW+CPpfTwNRrAZrSP/rOuCNki1e8BYmk5yplQ1Jrav3d4+ptPmQwiB7nqH3GTULGLzJ
98Ea87SGY+4G6YpAGtZcrHqjf3jKvyAc3wo9L/rN6ml4DBRsilhLqFPZrwWAgPQRbArTP6ySdAHx
wS16p5QFPdOC9myJplQut8zcUqUaiw0GAQs2QIh4m7gtxb0eFGyhRHyRhx217OU5sHjp9NTGBAlJ
s0R3cpHznkbBnMOyoK6AYm2YUX5QS10Jqjlq7+inxS7kFRzD5uQhU1kkuWkNmB5ZHkYACEXrXxaw
+T/yDEVHxiFIKb44MxgO4ACeBSmryH3R4fPb/47MN+WlQAsN9DeX9iPZLkUNezkyRul3KSn3SHR+
S44IblV687+HzlenXnaOCjtAQ2HgbHFXl9BSuzw1zm5Fop8XoL9YQ9H/o/qqPN5Zqdx6+0ANYgIk
5QEXS3DTOU05A1s86IlifU88aneYfi6Yfx+j1GEgFPgiOfrmJdk8IeiuC1EHjJ07np3quh/xNizA
rXoUXWuzWKh+Ps/bD/SewDNu7b38dzmjqaSrCC8ldEugCNDJYgMkztnGacPCbLZqQ9aHW+ecZ5Rh
KIDEFeD/xoYniHkvbGzsOAg0sqabhyKho/3+tXMp917vZ0FTv153aMgpH+UsVgBElX+8tr+t1I0g
F1sznD+PhFG2JcTeNX79Gt11q4lpZ8ANm1xKVUJ9jm/c3KliCFa7ybN0PZ51ZjztgFcY9NDD/9Rs
MvfjU1LV2lLPa1rCCOpKY9+shYo9PNeWU5M69tmIkfHAXcKkXjat07hv4mHUrJZjJtATC5eAaLQ+
K6M82MhNMOkljqoj4mDT1QHJP1CORcHQlz8y+/JqRwvlf1orbmHlBszrwooCDkXHTenAdE+SzPZl
H1RFwsmdY1556h+X136yaWwU0K5y3kpdjBcGBdNv9ra5Z/z43eKE5NH3voKz5+zZw64nO+sT7phS
K3PlB3VQG7K8wod8iiXPYH0GkP2KfZ471f47KJpgadmr7ns8B0kbC19+3pUwUP0/qZNhJ/bU8mYk
Vd4YjlBxSBn7Ud96unQhELqbqWTv2mOGpeZYptR4s8QX4BlbqgdGz8dWYKbYL6HGUw6weO/ZFyIO
9dxmSXdNSUKjdgoRgNvOG8qq+5Z7OWRYFloi4lV16WdB2YcJhjRejoEuZZMUzcR6GYdA8uEL5Bfd
4tEfJtp01paalVhWe9/nEYbhkqa+USk7XqVcM883SDU46rQHZ/0QV5Z5uVCF2s7SL9nwfUoHLJG4
FCUcujZqH4m/YWdBaa5jTet4goCeHcPwqG+PyCJNVlKvz8nIg2zJ9xhYNhunkMmhemw7lu+WWimF
lUUAUybAOGlPUAsT3KZlku/g6ZsdWxgxVWk2IPmwfq0G8JoClGxx72rEp2H9TfTwd6rso2VSeJc1
/nr0FBkw+ufRrBI1++6J0JPxQUCOnV0b8se6PQITY6AdNuZdBbLTYy+0C7C8gfPKBXu/J0rzi7aF
neApuN1pBDXSHxbIxXLx6FFbde4U7djfBhseLQWEEmNmMYLLC9z/SekvCcilWX8xu0ilH/G9JrwM
6q1FcgCGPgGywW13r4bSIgNjpFy3sI9jGMf4NgD5V8bqJ7FlKvzhvaoykOMV5NiMOPYN1p4QznVg
JpPWi3B5YYtwpioEQWaxMEuTWUDk/rkkrEEabLQcyARNYEzDsFIXz8DUdGUjypaZjAbSgXyqj8HU
NGqV5o1uCeSazAbZd8epmmTkRYXb+CRGh+CpQdLESsk6H10pKin5uM7uc4+gwlZv+wH9+0fdk10p
TxiGGAVhO0tvoMC9jwJqIxzw8Vrw9TCqGJUzLIKPwLYnJB1GAgm9MxOxUVY3d1Hd2xRvJxus/Ae+
KXx9kdcCWKoMYn3QFM8JAITkNtHWw1Jqu7iUe278EDhfkFNW9JQ5s21Maw2qYjFlQ2CfEzL68PUz
R/UVB3sj5QCf7shPoStCA/Vy8mQfJaSXYPuRfZn+4dbqEXUQV/Af01Bg3zvvVc9jy65BJLjCPeVy
g1b3/pZp+Zm1PCReh+PSija7qCSoy35OPiGak8hCqXaYuQd1vEjZwPXBLoaUM/MZ5HkLqHeXGlGn
wUBFBtyqoMc2v57rT0i4FY0j+oyhNYtRyHIW4I3XAutF0La6pPBQwBsneuCHTm5xfInB7chSeIK1
YLO+w9v58QcPwypJ7iLHbxZu1kdPNQzJH4Iu4oPxpGaYmEgqCru8xJfVgSaGNxeLQqAT6dftR2DL
DBSOENbCwTchHZn6P9W+GwWpT+7j5gJSDdXNByBZKYmWVo1tmNZCxfmAUFZ8LWDrSiEZX+jGeiNC
ul7nlbH4sluAj/B7/tb04XkcUruVvA/OmxUTEjIUgkfgL7MM0IStI4y1aVWDFT8ByUrMeWhLUrE9
xmqQsmkH65hdvcwuLDVVOy1lkb1yXaAYV0bbaJOAUfVOZGl0nO1OoX8mwRmwy6RT7vC9QZUWfVVu
qbWOqQKgUShn+EqOhc7x8flzFX9d++3YcsIYMj3kANRS3v59dUBOYHno6lcn6gVyPl2qeVbl9Uk4
PTR+iH6kogd7CXzfNMrksRaenVQ3IHhPgJZNw2t8bYHq1bw1bzV9fhaDHMgfTyS9pRD1X5W5iep2
MBSnaJ5zoDf7XGUl4BDLkh8Fs+ahjDCN2g2l4RrqfdL8eTq7rJ9FnqVb6V5DEoAS1CBlrugN+SK5
9QVniQcGL/cDVLU0xIBm0tbo3L2x6ksOjLxVWXEAVRjzqZlXz7RkErnTiLndlSOp43LjQSnJ/ocb
ev3DE34F15m4hafQ+LDlCX4GrD4BBqcRWOnbsPU5vlmNRh5nU4bQ08QMD6XpxbBO86UTQAC0xoHr
RK5z7/h5g957VLFkVLeWkFahfzuxoXErz6ND22ybJK8CHzCMGpxp3Igy6EFJYEvx3pyKEZWcIAXd
c475s/qMOLwTnXwbimx4TtVLktTXrWsXuwEHTThplcw/hPwrHFoHzNmujlTRxvR1+cFT2FsNtG6D
8xzQrsmVIXH2LvvSA2OlsphwQ9E5QMAdnukisU6z3zN9s3FVLw8977wCv+oIcpmIYpr4WJHfZyrR
X47rBmZJRyNP21l7GNEr/WSaIorRG0xnVkCks1gNurXQM1TIfJZZv2lhZ2vTU2WvxwBDgxVVJ4Ms
4YYybl8ydRaJYrXOIzflr8I6mYll0aSm0ubVYTKF2Nc5RaQKblqxIA3HAREKY0DK5/3g4leuLUIg
VoZQA+Bvn7UiHcbo/0GXts8to8B45F5WztUiWDt/g9NE3x7UWdbpd3snIGrNSR0AZTwM5dyrxviG
4xT3pTMAfGouCmF1kjTwa7WoPlBVXss8oEYxVY+JcXa2qz5Hb7pVuNJPrQvIgxdJAoFY9amFF1ED
50qglE0O1ShWcfrsO3JRbsYiF67rRyNWSWr+AGZgfibfOE/G54QmIca5iUvZdr764DGc7PWhCy9U
Zn20mX0cEs7bS0mKxcK1A9zLMzrYvwjRg1BHjG9cVt+tb9NrP6XkiG0k9r0DWuA718AACTprN5iw
wTJmJm5vO/k1UCYMprptK1iVFPicGKQd7jPbSE976SV8ww0UQj8OSYIEVvDwuctApOymOswGFH+9
73SfREnlq7/b7kChiC9ElRM1rUR2YFLhDPTJXJWbCmCAd2M87BuXB04VExZmlQdZA2xDwQyM4VZV
5fOUUCyVTm3hb5+mbkZnITZzNtHirsxSTa/jiyWD0ZAXZy3IP6LaL6PgRi184Cil9i6XW9VwMcAR
7PYkdWlvDCeYGII5z59Z2N1dehw11jU1KKIN5Ymyvc0f1FEBTYZMk0sjphD1cOfRoqKQ8vvAb7ZQ
xpfjtwhl3J8UmMEicnFAPddXIIIs2KYxT7tEBQiz2d3aFMMVeQWFy3KGrhMCNzL6gsjxV32uRKpF
N+XXIR2liiZyZn0ZH+0WQ5KkQ0MlySp6zzhpilPz4fbMPxwQOmAc/id3KTvvA6eqCY+3JjY2V6Ab
CPpq7D5l8gzHJByGvtbal+q2Wxc/Nd/JaxCB3GCVHHN7Ifj6ZxC5WjdHvHoETokQvMfiUtvJrKmI
H3uOVhVMdbHntrmk+3LCAMVPx2aST0L1CMHyvhVS8SjjnatRfylbDZCVXhqUdxxvDdScmMCPiNu7
YL7NXPvWlxeC1ZuIuQdJpdwjegJUBJytX2Ya4oXOt9om0CAM/GHv6vEp0cNSxsYDX3vqaXyN4XD8
q14UUsQIFG0iTq431BlOcnTrLfH/7oZqaMChfDGCPsACkVZ+uxgBSEomUxW1Fsaan6apWCA5Ixaa
hX9wSz3zYOmh+HjAx2yp2lNP8fUTgwRgaGLrie+6NOTKqw97gZE9GYp8rdZRG0KCcw5pwkiAm3kH
AioarnUdBoui+51UbO3C/Sw1MdDU+f3+HDoXs8ZTF7s5xwMGCfoaTA5wMxl8xyMH6yPSUt4Qe5/h
vqjfgvl0PK7OTatwk+WCFcrl1SQTStNlXPO/ba6wjziOq1K8o2+ykvk/7pmnP2j+G2HFVZB9vUYx
pbpkyShn0yjTEqINO1Y4H/VI3b2lrvllxSQAL9EeisYzoLutRhXevdDKBOaQp/aQ54ZYK8V0MRmf
71kS784DTpCwnK9ZrlRWo32A9Jv2nVp2tGBuZvTbCs/9dRnSjlUKncs+tfLDeB+BKh/ZqzQgPxjT
7HRoFRfmW1M7xQyltjGHUrwqKGUppRTin5TLOVMvnXmUm9aB8uHrJjxClvMJgILrJYDPyhZFBPGI
zi/njfjqtncFAk0E0hUVgqdMdSNZQux3hUSRdqbMKyNa9Vk7gd7PCSw2OIzVfnSBBN90JGJOTTSq
ryHAIImLqwWLuA+WunZbr4ZC5t6H/IbAdVjDyaDMejg1VEkIMqJWpazGjYUycqo3TNUmOUQNe0Wx
PfYxfz3BsrIEtaZMJwWYTc2+6b7+KL6K9qgxjYWxs1BS+X9KtDjiRisYkxmJQ4gjJZw5P3lojOC2
ggHILkM6IFhqmPXjb+bLqSRS81hyKokRINZ4qWf5Zw6BarokbbNQCYy+x7e2NKAsoGopz13ab6qh
f5hKCu1Y6ca7hDMwDiELgkENquw5On6IkqXS2PqYUIQzQPZJIkDl5m4pBVLqmShvrssvZw03/It2
f3CZwOwpIv5rmgn6KQPmGYVb3O7kISkUcKO6nECYyZciJyS29US5tt5eNGo3We8OCedXk002ZfgI
r6oYdiiBPKKDiHF+zI4mnLCD/Ez4KJDGHQZOBwQ6FAX1lu8e4QiC1gT8lznS8KKH2rfWv9iCrgnd
TVimTBHGr7wo4ftg7XT6l6DdlV31e5+rfhjL5eN+3A3tpfrJ9+jgWX5D17YD+CxaSz+ZjA3G6Xu0
v9Ud0HZy9Ct26feK2cz5cxXH1SRDbzrZjd7qcWfCYR6K+8kvTaQC1UmNYJbUB5zIzZYLyNLn6Vuy
9r2/Ipm/gmKEL/JMPoQ2yLLudN75rKd+SXP90gNijmVDq6EssMnjAhJjZhaCOxvWchn5zGL4399A
zi0LScNYnCEPb0eA9jTcfpUeXOX2EH3TeCZyaOUyLl+olyh39stEs7SFnfH4KW530cYFshYdX2Wa
DR43+xDM+zC4f6M/U/YSl+MOnK9YiiAof1RQyk6suOrJP+hgMBqe5A+OcB0EJLKtl/dTv3dFu7We
9ZGoUs7JktG6rzAiIFyLnhhCjGT65CwY1505TVZAnTHyckroMkJ7RGCMviDlkI81lLQivYkWeL8y
booixyUjjx2lGj2ZuaencPb0v7VzDrRzmpNYSZLy4x0ooEwz0+s/UVfLe5Hy50b+dBn6V8Jz7qMu
Rd2txtEu9s3u+uo6OCaxpg2ocsZgEZX2cdUyoJA1MM4813IKOAUdjTej+1i7W2yDb25FsjLed447
7+vTrT4tK8jIr3eHHO/9iB8G6W7gb8I8qe2MQhNJrdYFQhzj+AaYFDyq4SspFGubHVFs254jlb79
BIkWnS1fiYUJ8Kk5V7EFI0nJBA8Oa/tHFTB1mdPxmdrNXXhB79NmKeTr9AyaCOx65OMh6mbSRGwy
O9h4ud0HyogXUlEFKzMhwlUQ8D5QDt1Tyc1eswO0cP4DdqyUvnZeIu6Bhu+awQ9lZfa0zDag2BuY
HzT9qwP+saR0dgntK7GQRndt2Mith6+bjdlgeg8otaJN3asy+CE1T6iBV0oZRy6MHQhqu9jPlr7U
yaya0nDUqghQvUUc+CbD/zWAlAfliPbSBnjum+E2+aqgnFOXL6jPK+4kpJqDO5yyTNrgvMIavzTV
Z9a64oTGTcmlsfZn/0naX6weTMCOG8ZKn3UaSl6zAVsU0P520i1Ynj5KexaBm45zcj608wJlwSIy
AzRHVxvvMGwzhtLt5Q80J61X+yp/Embt0smMjIjXr+CoyLGEgtU/kjkcEM2ba/lpqKvoE4ZMmdVM
ZKNgOYPmLO6C0M5WcaRWFMJkgOfOE5p2/nrEnJd+juxoRTSzK6Nyry+vgjOFBULNWGcFJ2MWv3Mj
KGKYNFDaXbMsHmLrrmlKTjxJNs+t6JKx/MlaZpJos4xwYdSQfxJ/ll0BZQJs8o3ey98tV1aQmC8B
WhdlwLA8apHg4Xh1yNoraiQj2rlnfgO5OB3qAKIAQrFTu0fXhY39GN+kQVhF3JOefeZamTeqcm22
GWeVoH/LppcKPuAuXVq/iwlRseM4jrw9BLhhJ4CjQ0H/75RX6OE1NeRrdsTgOxp+TkpsSEKw/38i
OWJZhKsxwUU70Wf5SXk38UjcSekCp7Uq9ucolAYOiybJExUePCMwM+8ZzzSIu0VljuLU6oUh9ZgD
4xB41ZxlDbrR8TRJBt8b03gB91AVdIC3UR4QzSdNM8BZoRmw2ESuV0Kozl09B+dNdF3ToIzTnuWu
FhMuA0PtOkF7XH6yGGqxJi6VyMCgEOGmuFy2H3qHve1iv84f+eJ2VYblSEhtIdOU8dqANqF/kGlC
TpDgIL0YCJRI2GVLzjz1Ey2uHTYtpEKoqCzutXV4bxHxI9EbENKKSOSG9oy24DnmUTHnUtSBhIJd
MtdaNvJ3pGEdv2fqe81IQZALVhSaaulLzUBYmrglgF+4HBzV0q/EfOQMa8DGuMPgIksx2VGgs1Ap
AySiEsNNGVKXUo9M3m5UylXr4ZsxUGNpQ3npsr+8Hlck2taf1GsJ7wwqyoO1Wk44zA/OLkOUlH1A
lWZIsfE3BnLcHtA49Qbwa5jB0Y2Mzo5LN7Yy4BI/DLOdND3Izkn6S3SPdUPntUhY9jF1hDD2Eo2Y
+TC9TnXgskFopqURstPgKV7TqWMyZQ3g5Enz3IecXS6J5saegRHgAGLLCIre16IoYZRa+G5xLfhd
D7dU8+mZYjDJfXfTK6bU6XglHOfiXFePoG6i6CXDBhC6wvq9LXimni1AiAm0oWHHd6wPM0f9BSB1
0W1w4HeUcq74zv4eerj3UGLGSQUC4gXf7qsICGZS6dccni+qd6ertl3ON1Xr04UEGgHPgvnmzCDe
Ib3GI74Xk7CMwcVT8O51Q/Ki/LUwSCPzPJHjDydUguNaOYjd+lrtOA7S0mLqdxHUb7znQ9KHrSmn
vbThySdY0L9WqaiL0/mxCwerm/G2/SHlCSH5mbieTn9Qg4iEs0gzaA1yk7t2Pf9qAtx5MhPFr0Sz
mt50PVmmtiBBVc+ePu5uqDmjsKbYUxhjwRshG8AfLlZnLYFCyaNwprNNBKza7LB61vfLnkGQvM5s
ARrf+t7nXaefIYEj9zs4QmqcCGEXh3sPEkgaBiHwO6BDskBpn6Mm+MlzeXUgiF7MuQZF3lnChVXL
MEumFNHcxWbFh/Iz1WUGbjwikDyA4tHMXVkJlgw/ubiFK7tFe9CLKzFh2dWOEbuAjGIEvV9JnQ2u
QxmuZEsg4Z73WSZ+d9Y4W8qIONCW+4EfrLZUNEjUW8zUwPldQGdv29ViOi4eqh11iQcV1JwMHttd
GcYStRs+znGYtdhgmOMs3EZ2gr1p+otM936xxKo1ngUA4f1Ni+ZvxjZlI4ElIsOWKpifS5qP1FGi
OgnwhV34TfvL6fCmLs5/GqiYJm0Y4J1mrZPhWztTTnQbXHiQE6yNiZump9h6ocpsr+orqyhbo8la
Okuz3LhXRINrXJ77L/z3MVoNWofm+dG7HzIdsimLZiYRga8zJmX9m0wWPR9bgflxAum5NrfthG7z
hObm9gL0Ea4w49AxrYRilAKp8tpjC1nbdnPwxSUthcpeXavSbTaT+kijDGHEoj/glkl0Tf/tJzYw
SdK2sQa3rRE3ZuaTukqo7q/NeYn1ORNfmpOrkpc4JtsKe6jVwkvmWnZpn6zkp8JyQq0LI+ougC0L
uqL60+F70cw2mdb4/yAF0Cb5WnnABzJ7ga5qB+KwyH4FbPCPhZdeKkhTJTZd8pDMq/P5NVqUTIAx
mwUfvnsvB3dztrKR/hBHj+vD4mrz7+xN3ch6kRYTqnD00zLUXtRw5ErLrpzoILILoWFmU0QqeLpc
7LOdVHUTNxsmJU9lKgXOTx5H2AsMSTCEzS6+8EENyPQrCDr7M0aG6gaDCdxeO5ssLG+F4zq0qQ7S
hZs9ZxvI0O709A5R1I6tItaxINA9U8VT16vP6sudVy185OZC6fabXldCYDeyageq3sJwRfyh+XOl
hDB73paxCgGvW4R5h9RmXxcfyvin8LMJZFj4m7WmdH0Hk+gu4BPuvMQQFSKlkymrSgiEs4ijw9W4
pz91WM2ZJqCGIkCBh0Uyz6vLYDjV91yZKpIsG1LsvSDSxhvugzGZeF27OuPcYPhgS0LwQSkTx5J+
VrUPHiDCskkiHNkG5J/9zN55sIBXGxnOeziEQE3XSvNQVy3GdUIATKPU3q7hdvu1NL+1j9Im0WnH
R+Kx/diWsFPdgd2G/2HySVvLGjkhwd3DOZmYGGGsQ6OLnih8tjFCdBx5XDXq3i7uesBZXF499ywV
YzCYKoA8e7CZBatvDdeq2helWJhv62wURh8WbYvLuuYNsEnDJwsmwALEtnIdmC5pKBztp5hg11Kf
QM6RCgJHapN8SMO8o9jb/jBjJ3UAkw0YbDdRNKT+v2JUJ59yqUUGT3yJ0BX96hlfdVXISXEPB6X4
aIHuvys1ecjg3qVMkO95PjToCCyOofxBTgpH2M0S/wnWTEnCXlbjfomF3VGQPWTA7A4uJFy08asP
xoWB64bjoLPSPLW4DArct4sOYzUGu5R3D05UJZvOsALWogi+LrM8/hqUBtb209nMNYhegewmj33+
NjIYE3Aroboc51Klv9i0100/sA+svwxDEV5jRb7sox4IRa1YPkEiw6eEWdy/NTP5EU7Osz5j9dtU
1RCZ1EJcZtHP0KaHRAyaH9RaxRmBgG1DFtQGFOcWTRBsMhD9+GWk1CjMdMMQ45yW5qhNKzh2QMSn
0l3sb8y2ikcHpuuLUxc2BOe86Lu4eqCsio/BF9nqf3BcknvQ6aS22L7psVOvFKrmxvlUfh0H4iLS
6Oa+gm1slugMaDxJPs5a4LdUR99ggzqNOo2T2EQYydxl7qn13XkF1i/xDdCI+eykLKyGCHSPZEdD
vs49rJJ6rxh4jRpVuJaaBnQLMDpACM+OFoZbCQn+eQgNRl5gNiBVNyUnhBzLCmowtYNqsf9V5K9E
lWO7eYCO3HNAmyCo2pZcnVkDjFjcWkN9w95PmjeYVMOXszfyYLr410Z8/Z5h7mZGDj96KwscYysK
k4XvrB07wZW4LpOgYRwn5NTqV+jDa2GoVIR8AtpMHqQEcc+gpNzjkuCRMcmBRkgGZ/F2fYpc0/dU
U5ADyWPUZzAXZvoUZhaJpIWB+oi/VCL152WSlX8+QygMEqsOEYAmCkUrxw859fei3EO6wh1ucrOY
ZAjFIpKD4L3H1reUfo8ROwjSrv2RwoC2COPQoM+MM/7plJtTmDLjtZvD9FkzPAy8sXysKVTZIN0+
vdr2RJuQg6qG6rBsbqgR+9Pzug5/ff3E0kFRzNF6U8BLv5E1QGToUnGjkyZyD6wwxmWH0hdU5Kil
bMLesujuhFJ2e77vBWvcX40R5mpcvL/RRzbM0f6wapyTbTchl7blQmlDXp8Q0sD91AgbMwy4P7rW
9JnFjsLW0w2b1RoRCzg4peJoN+IYRqzjr4SDDScuWotlu0xmSCStrvIRsIHHU85mmRTSbFq0IpUF
ZrDfI7agypE7QLGPWru6IKFO27Z+9T6PPkON50qmyHYM4IicMie/fp3AzE69TlVqKCjsjQOUAlMp
rgCk7suZCXNYVFsUcwT2cQm80diFeBzLybY6ihZKgSAIHeUvy8u9eMMPhuXQwxMxZqK1svjJUTy5
gF16oIr+6/x8ETyNbRcpmZzCz5UO9QBV9fzmOijzYhd5gy3gY+LhKx73OAJpmMoDthq7pKkdDlHW
7SUDHcOaPb9+0E3RV4aaqPYCYG8p3jXLWVHoW2XBH3b0D6I2v057WC4j60AHORfwx83YRd01AjS2
iY+MpecNwfdSYwID0ttQQRBDL19NfQIO2InxPdq2wrjySH7JuMjoJliedWzpHZAeGBR5R7NxhWhg
ZwsWOjUN5RTeb63xgaDLSXUIlnSu26qGHk9Hy9E/U0+ySDYNKbsYbAVAjZSKXUEKV2n9pxznRe9U
q8+deWSrgRsxAn5aaN9k16mXVgzHsASwL66zVgItKpjYIWv470FUZSmv0daOV9JmtjcK53+IPz/O
BvCielj2KK9dvZalk3jM4TJrEMJkeEZa2BhdfSH2KW6N8foRNvGZLmawlwLB0chN94+yjzMQ3mEf
D35HX6Jfb6rHC8X6KFNmv/oKyCUCo6BymYTxk+RckTqLtW+dEfWcGb0LBhsCcCVnCtmdMs5a3bh8
MPFvjNOu1bJ3LWO95NIfbrhgXjNwJHfcKqtyNJpOrUfGrSQLJj7WYX4teupMEaaUohil2A4EhNXM
y3MGzCiD5wfXHcxhMbTo9+m0vGtTImabLPON1WQFXDzO76PnQ3R707AlW+C1WKzkMGu4VCEirk3K
whMcBCMFjrUJ8QVN0ikL9uYDwnCzgxkjo6lCub/uccZD/WpiULRFP+jZKQwgXDywdugn39HGyMhW
wDiufyzuoxdSPOgEx3dNTghGLLNZHgB1UfeSgaj9kPFjOcQkb7PxgihgJ3vhAXCp158pAuOKut0H
HyO4vAK7kJzwQnU07JOjuv0se2sNrLRWS9pojmEne001q3Cw7j90dHV+pMna4DELILQNb8AOljAa
wd7iUj0a2TJiyYDXxcYjXfJb7ySWkYa97+Swr8oXCAFGQkjIhio7db1CLaLJPlTJ8gllobYSPuFY
NLcYynnaz5ZwwGv/HWDHvlUwEvPhWnQtYHH1PN0AEPoWmxQQXugFIULWh8UyPZwDO0rFnCn2hgcN
5xgKrg/JBHJGiUmt8Taei8Q67ip8INhincDGiL5pxTKmlClMJzuqfaeL9FN7FPk0FKZzqHHTusNF
F/jx8ReLFgASK41Og+O8WxBHxT5sixvWwEnk3SV+5+6Syli+ozSaIy4FINF0QDobk0lbCPEWoLDv
uGXP51u0uLgWgKVH4X4hbGqo4BbizzECGQBlDjSMwmnpqFMOlguyCrCXEueOD/3DoV/H1MqSetIo
04fQFR85uMmWE4gCrXB0WAyDT3TmrHtcQaPwy7u4frqE8tpgWDy+2ZUDNMQIWpy78KknOlbb/IV0
LntI6EimJXlAUhqJjdqI7SJrPPbu9rcCihurI/SUuXoOmfxzoTX/OzNSlsv/Eg78ZxcA2IJOrzsf
vqyrFKvgZT97glVMvZyTtjMo+u3TKIeLrofjbvyFQSAgNJsXThXAAkA2GZd/4s+NhteuDIvkouZk
IPuA8SoaxSPzG/SOAoCJdcJr8RbUXRF8l2qTqOecb5dt9dJaVs0obBIZjaymuJjIZcp9YG3+6AjL
A0lJZiJBlR7p1w2Ib3nD5F12FQWMifecVVsJwUWygqcGKahq34D2i1lk7iK90oLcXUGHGzannxmM
sZWHGqR2D9gVO37GiIDLKtvkNuClN6orqtzRye8JVYFLAe1bv3Avl7x3G7wDbxsQZUFwim44OJd3
WBisiFQip6nRju2FAg44iJ4PT8gf9sC0JKKSb1cz4cVsFkA0gDTopPTRoTofTq3FgwWdaYf+g5Qn
p3/hYb/tE5xk3KnkY5eVVQFitWTg3ZNQ7JEZBLtAB1lMbbUf0o+msk4apCCAHitmCgty89s/viCx
HwQfXQdqfP6YvI7VU2Eo9MQ6zwBnhVqj3V1D5L2Dn+ZLjiSxw2FPEZBKHiDGlDAfif5zh2b8ZYQf
ggM4Tvw5Yb19Vh2CSs8nv1BaCwSk5q0GHgdKJt7Oi9T4Rd4CNZ48Fq28xgsjFR8Wa+WYktIiZbcy
S/6Y/SYgfbUc+pdio8nlbCeBiUTmqgFIibpDjF4bfJvkiI34KnHG3h/SDt2aWAQk0OTYq37PmNYP
i0V+kY0L5CkyonBSupS4I4OYsF5Geg4NDuV2P0ltFq4gFn+BJ94gDVMEkEi+nIbZgo+hZ6SloCr6
3zeCgI6LVYIpGkfSxBF1Q5WcIZ/yDXi+3EFxC3Uokfa+HxmNfA4GnLOu/IBNq3rJYpHCE3wU+RzU
YA1pK9Du5uor+ibxTcUuaUuCpgOf7UWw3GuEsPbNy7nSUJCO9NUyB6sDQjfUiW5xzJ5GCyYyPztt
cOPCy+e49oFXWtfLPopk0LErVtlWaCZbO6ickV7PqDij4cMLD56EAMlpMveMrcXz8dopqKvj3kFq
cTq0AqL6aLmPGA0wGcFVQRBKvzaM1nji1Fxl518TZ8NblqMfkzUal4TjnlAmlnmkPBqIEP3dQ6J2
/u9zCyMCQ4G2ZA++lHgzEpuOSl3/MmKX4ZJr5SdQdZqJBRQLteayzS3JlWCTAXyp90kWLtrahn8s
oYp7Auy/AHgBA7w2nUdnGZG7ItqxiORZmP17x+ROV3tKu+FYAsxoPZgJfBFKgPNurqXU80p2vz8T
xmrbXiGgMO+OlThJGRrvD89i2AQQWDjcqNjEYp2eRl894R6ASlN/XMto0R9j/wQm1YPS+LJvNTtD
7N6iVoU3vKHZDT+CYK03rqi2Zj03HLepHciKV0TcNEzUf11EDHjyzmAJ2N22uo9FszOAzOxWnr4z
kFGd+ZQtvpzAgo83OURU6TUM+EtZc020l9FP8orcL25EfxRRtokpS49kQ3030rfuRFWAWyjR2zH5
iIBOLNZe3ran78drxcYw/cAKmC9ZXhQUaji7M/idTXtsOBmr5YIZmzcOPU0hdcVK5ElcTbar1/k6
eFn90ur5aAO76Swq3ZaqOCnIZiuOGVfjEWtoE872v1Uj82GeMTuhm8eOHWOr45K30ajCpkcQUbYn
CIxIBuq5/iRpCl+sV7nr7+9CM0rE6ncZ+gswt/Y1X3XzS3Ei1EWSpx/PXaNfGVyESj8RfEWNBLC8
98GwZAWCXLP55Ghp0Fk97Wcn0b5ZW7B6/OXwUwHykj5YMzQOJ6BbkjQGRgPwWof49rGBvS5AtcHk
o2ktTWN7RBAC/G8wxs4umftkjwrbsoof0FPuoxy325Fzn2lEWdiREEmYBYfxoIG+scSFLFOcrZN1
opDMPRU5fV3s6nJUXbXU+s2VcqWk8sSjo9V7xjf93GW169v3Jqah3oXnlXYuA/ki8IgxUNKMkgpl
h3r6WmeqWVyNjSgj3ms/90i1zdJ3x1DeNTyQ3lLHR4yMaFgSbX2I8Ag1eUugb2Um/EY/SZmVxSwG
CNYl3zFe0qd93IyYBpKejv108GUULSIcpa4Do76EkQczjFsDPvqf/++SYinupe8JwzxR0wM2vCJa
fyAkyYC6s3K62/Xkvc97/0JewwbPpSuM6Q5UgheCq6qDZ4xoPVHnstjR5qp2eICFeG45qNvFY1Jd
WsZ3j16rzdUHPfUSrtfv0Zb9zNlsnU/INoAKfdZ+jNoBLj4sUJn+j4UtKGuPNn5vffSuUfvKrERJ
6+dHFslXRnbuasRl2EAj1Slc+Y7rE/Xwj2ivmCJ7Z87thHcDzVO8e1lCRXXCjV9fdbVZ4rs+k9UZ
scf4WvoyRa5Y9b/lfSed2bhZQs8En1chL604LGDgrqIGOQuNO0dRTGqksbaaElcFjKIXyU7OoktS
OWjrW9DULaUgh8BUXy+oJ6erdcjobWTlzzyZ6ktL6aCzb0Hi4dymAdXBivhrKAn7n0oN9rPZplmN
mhBRWRzdbAuQcTTb4NdjCxu88oPaip1SntYfcSihXZa2ef5Cr3p8gjmBbvhoDw+r3KtIkzTX2UVz
usKdOzVl+hvrK/mdakvAJ4se3Fy51n0NTklTwOj9v8HdMSimdB7DnFNsIO5u9EUZhzMm3436WHjo
PpUhtZd7ZqQgiM+UPB5EtYddzQk63AeGh6XZllQ75X6N5Bv6rgDwzi2PiZbGI/ymDooh2dyd7WVH
at40sf3/hwHiSowrbFuzX/nHU5NYxvnnD5+PaWTRIjO/c+3IXFvqiP4jVWLRLzWFN+UpWsYZ1P9o
ENAHhg7xUmYNsgV54tfd3EP3D8o+50vjZdnWdNH9HM2IigYcCEpAVm14WQlgXpSmBxnREEgDBlu4
IU6xGK44macazwca5cloOgZ0ePmygcL4Nuv25AdLLFrqNk/SXK61rt5DWEDAEt2jYl0VvhbfvI3z
ObAjChp65O5G34DkG8Wz2EcCAFJc/bYWHRo5gTbY3Cf3HTGIHKl5Z8JQ4CFz+O1Uwn6GaNoyzPkm
5zGgiK/pKtx5JXWHb4gQgqZQXbxH3hXsO0ojo/e9QbcjHlv26kiEdPqzWeXW9hnasrS5xarg83Lz
KUVL8XNPvI3DfLoPwM3Il0IyC4zHKy1lt7vDSlfyGkWZEdEy6eAVzLN36R93PE4h0U0iXjntAxr6
mYCKYHLsie6I/9juM8cQykR6DXDGSkF4XJD4ndgB1vIfB4dKCx6i+qE4a4B9Embz7v6mTp83TovP
IGH/0Za6tHaDzidZCT7jejoNiQ8zBpdT7Mx4uwQLnDiwV3u9vvJn4lO006u0iBTU3/E+gj/lFEwd
w/dBjujyYky+3yEgtHRQVP6X6g3oA9KH5mSNfgJhxHpn8WYSi351d/JDwL7kmhZtZ++/FEGIxGkG
rQOYa+phcEYjPsDaApS3Ubw28ckh17JQoiOtxDYmb/X6DPqhZrv509AR0O3opjWxz5ePdGYyZzrL
RJAJCTzoZA2Bnnj+wZb1vVuY7JeNx8gguqAHL2nzALqHcxzlHqOHwT3Gtj7wulYbYxclL6eL33AC
JNKlxsUCeOCGcu6DNgFff/fTZI8e/w4uChjUyLaoT7fhlovI2tFbBFkzbQ0EMXsq4oJzjIZGMh3Q
AocMbq23inMOGI1CDB92ub28nyk0cewZMdpGiQNM/Ztre5KaCH+w3sonuSA0SEvTa0VSLeN+A7kI
OUx7CdIIQhg1o6vH8eJn9s6He/UExXO/PbqfJR3oTBShaKBsUOHMHnnm2X/hwyv9JA2CP4smxKqE
TivjD4kH4gp81vtBDdCPBojLEo0z1TK4XZ3SMhrguZL4Te+5t+qZ/CZ4HdVu3dR97bMwzcfSGIlG
t4d1joOsc66H8yiO5MoCjhRISXqkMfzE/J08O6Gl7C/yeC4GXtJEv6KSZQWYreWb7Cqpyd8N4ERV
ZjbDAi8d9y4ioQuyU4/WCQ/M8xRhKNjW+MTXzmBjZrLyatMsflkIxe0kdIvUaJb9VDcC9KjFKf8A
zvFvw3BuJWKyFHcTK2H/hzgG8sjy0/hf+H9Kk3UOXfOq6iBHVZ8PUtsNlUIsiZAP9xu7PT1pkCNc
Qr+i4+BKZXBkrITCPMho26Co+cKIAKebmwCoanpOdYUuPUH9veeWj/4WvgGaG4njMS/y1Dka9/CN
4JCjSnBEbpsWvONUHdrnB1YA692WEPgqVMsaybF+pkLHUQGAlazuUkGzwYxLETgZxaIoV2Myw68x
X+jlg/ZVkXXagWNlEngaecFNpDUIQ6IOl+uACKNBOF0YZmn7IhehTQ19oPwKY7/q0y5i0qcgfyB5
g1qfCKETG6nC2uqLjZv/BRVOdl1Zhohzno4jUR3zzU+Ud9jI9gSLprrjjo1dnrcf1ehTN27YtGLN
cn9Cv8St0Wcd+bKlQR3jFF/JiUeToqFhMZzVfVIp1054alIT8a3odHsGBZjGk9ZZ65wICLLqpeUT
09a3/k2gnpMyOqe6phRrk8BQpNPHX7QWX1PFwXhaF3XL2eNoRmnSWXaPkCq5HRdTtzlQHNLZ8fN/
7dmZ7+cqWxdNwQkdhxTYrCLEahHu0GlnIZmqAX8XJMnCyn3kusZ+CL+QRskHCEKJ/HD3qjKIEyre
Q20eeiI5Vtz9X1AH1ctXgOdtWN9rSg4jdBQYbehQBB8mxhTLHHDgD6JaH4VUEE+4xn90Ho8R67VH
MXVq9AjXTomr9MdNntMGU3vWjWBveOvRgpG9DZq2OzqiRfHUBWqwLRX5dFmaSMLZKyBVL1Q2lxGi
IgWUEZlWBZ0wA90QTGioNN92OvIr1sfpSWk/PaQZfCzLKyxjRssbrJvaD5izvLCn2/dAb2gZEFIi
Kh1hmFSCbZBhyxzJbuGZ5XmRIZ0hG9wKEHV8sLLMtEG99I6CMo2xQbIIRbz4S520rLzMXKj1dHyr
fsVhxVYxoiwb5XR8/9Gob2OKUvTSzR25lo5n18jtfGTcLHvsk6AERa7mZVbRb1y/xJcKzgjmuPJc
tLgWF808hHu3Q2g7NlUcUVFpadApmwJS/LfHtzdjdXAClRVM9wNO5WFEMssP1KejeReclT4qo8Wb
N8/FFv2TAnzOfNHC25jdiEadv2wWFIZ4mGQCDzyslc8Fl39QnFS3WvHYuGRjTWlUx0IBGq3dyW5N
r8Gw+BrnTxjOGHkipSy9VJPQMHthM+U/rHdNrer83RBkjyMhqm87kyB+3x3h9p0qohNi62yPxVe9
p7ySJj+gSXiJbc5H8Xf5TMJsp5RzjfD/Evohw+bNLtA/HR37dWO3N2GQsJUhjErfGEu+aCKFVijn
WYe7ynJq05S5mUfQ1n9JpT6ogydxQbtPVF/WG6pRfzP9doj/5YO76JdXOBg6F7a1witetyrfcPS7
IKyU0xob7tJJU0X6ByRfJCUN75f0kG0nRh7g6dXBRh7N7nQBCVwOXT9ok9XTBV3BpevenB/oX3kS
LqmWN0aHSBb2AcjlywYMVY9HXZ4s2xLUxEr0mhHQLNBHDozG550E+tuGzms6Ele34fMWkGmcXt0V
of6Fb0yvIdSdpCqFRVSmtQvO52i2vYOTQBqErcJ5pzPGoZvJe84IYlN7oJcjEZPyVVyonJe2GTYi
l7MK6PYwMidC+ekSf1bCAoQO0fbFFi8PqKueXeBFgKMPyFQ15a9tK+NVFuRm4GMwb85Yn75+29kx
94TAyVw0DyTQ60j7sSepN/UCY7UH7Fb6qHrBGsWLq8DFT9Is3qLDIiywV7dJPL7DqGeaoM+OC8kJ
jyhxUVoVlkH+/faqdTxYCqm8I+9Rql9ZxnOOQ2zxhFV92AGhC968nJAocecBFycoAsgqGPtZj92S
yNj4rPMh/ARXRLRqYTE2RDGL52c6pz3gcaI+q/D2QwYteP71OJqHy75QTFu7IZU4D4/vNOMZic2V
x6QrObXpFxI+D6XHWBM23+EdkMeb8iheJo0ORav4VAC41aIbZo2ljZtI+bwbp0xWgtg78HJxTOAP
MAXj8duDM9u8QRBWq6JveCNJ9FXo4TI+GwuMommpEUNSO+/DyG0iIYu2hKusZkNHEMYRRu2B/PKZ
I7yqUtu71Nfqw0KTMoHzRInqb2U+jehZY8Oh53z+F76XvW+oR3FIB9Xc131EEY/jVhZJTQE7BdV3
HAeH1vWawqjKE8Dq6SiaNt1TYcJFkFJjfednbLbX8R60EHyLpitbrIsXUdnjqXVKDd4MT0fitqYn
+t15dEF7/5axxr2h2O2eO0IcxHrBVD+lxA1+VZ7fbfA/9Wp9Dmo4PZQs5gQeXMP2kvBQWbg0dXkA
RPuMl9qScXtHlO7Dt0exMfnMXzAMgmLQlnuW3Rqls5oJ0ya3Voh7QNZN+elQVUG/vu5uAXfhkexZ
yGP+3GC7xgoh19Rn2aPEbLfVV4fAtQIae9JRv1bk/kxGwi5+1M6Uekx6z/uCf71zcjroBBM/VJm+
tpdWVzxTUCcGV+hF7GpqstMP7ONPg4NaM1dDwv6EejbZWdMUWxPdxlyJZEcUuWOYAAR6uiM6ZJE/
KYa6rPdhGr/yOrFZt/VhY0tHLTXFejk8Z4gx6qScqHg1ScyftJyai38k7lYHwGk2ZTXThnL0K77l
uNnocTXg5vw4jo5jPcbYWMwgDvbUBHTXz8QNC9iMtwJC4l1GvjB/Ct6l40aIpY62tirOke9FkKS5
pPg1N8kB9Cs0k8ZQCJB346H66vIsAu0b/pm7z6qKUxPsH8+UrqeP3vUmANWlC9yedEY98yVhPVmG
tdcKw8FobU8sjTIVT1yXlAOQwnvDfUT5FLYUDlfsRJeOwZ1LCyFWSLrR4j0reyMa5H5pm+wIxHmY
IggM0B7FEyuVjGPMdmAfQYl5lgyfKUoGJymrRBblOcV/w2VXp7gxqRNoiE/f6vm2+LHE9ZXHdUH/
B01i87QSAj0GUV/ESuNsp5gRjxR9YgbOhdinqepp1/YAwOiEl78uAPrEHexMelYpeGUcyfZG6U/e
1ITVVUeuwHHFlU3DmGtsDb0/vjZwunGaFXWln6vpOx+Siu8TfbOw28yFaSZJ4wTUZ2IXOdT79U2p
qR7bSRMnzOJnxdNvkLtNBXmzw1vDavVTlHQjb3KPRAN5ksMUTqjqKgZGci+lZ6/UCdwxVZz3BWOx
z8dreIoBmBjdXVWQ4G8dGe1DypPLjGwTni8vO7klwwdjExe1YBdpb5wY9mNGQPoE1Myt9LEjQKVI
+jQxehFMBmHu9+Xmo4PXvBFAj6gVvjP3yD3AaORvWsr/jZkg3mm8/ULuTeC93TLvqa98zoVi7EUO
1sTPL4FrGpXO2W7LrNhlFu5JlP32exjvXnkRsFY0czGimv4bCSuEhA1ccJVsKw/ImBAm3/EDmyQY
MQJHYjjbLHOKalabIVQx+MjA6kNR+jL54QliqNOJPbnuX/Gi/pqYg89CDq70wAAIMy6XAmskRoYJ
MjEpC4jHIxhkH/B2js0J6Q+MO5b1pA+9RqnOv9OnxqgyPSIqfeu3Mz8cDadqsa4FI2eq2voeOZ2D
/lQBvdHNXHykK82pL+dhQJABVHEnuIDNJ2KtdQZO7cfE/U4mehGPsC60nPt8nBtbBEPhAEWvQLKl
7RuT6bK8j3vv2ScaBxi/5tJB1fsbD2AoKpS2hU51DB7E5cHPO1jK6BaZ1ICQRA9ECWGTJNUL9Pth
O8OpyTarbhIExA/ktYDx0ziPSOrVW7Mc9BaxQcAjgle3E/d6mYLJSHRpELt1O9P5+LZYd149apDR
utlgsap0zPIStHayD3pKcp89HQzlSwFz6WlzJ7/yv8bO9iES7eoyhinVPWFgwafXKu+uT0wXoy2w
j2b6xnX89gpcbgpMHo9M1OA0zKZej63Kbd8bz/Xwb050fhK2WoNmSVtkKDIN+akFX21I+banONfe
33Nx8cAtNN7nV8y2lgD/TrnD11xKOBFp+ipB0ft8MK9HXvB6q0BRmqezFnZ6tNIAuapXRlwigO4w
lMC0YjCyeS5ITcKhCblOg012vBQrA3M75pkjyLIiGzq3OxFXtrNjOdcCtjSXEAL09oLrDnWLvLi0
DGPuWGpAxcs04m/TVF2kGlfY9fxBD+90Z09DlomnDfZjTPxUzvV15f/TFkabsKjFCezrkhPL76t9
h1aj4idG67ov1RhpRmwF9S5/ftqWiF+sh+I01LUQoUAEJ2A4rzC4p6uY74BHkPob7kijVXJf49nN
iF5gxc0oDmAwjm/Skm5cvAVPUzfC3xyOIyWiHnSSG+BuoA3AT6rwAZVQ6VLAUrQluDwMhTspoRIj
bYu2/hfYKHmCJ0xvULpu0MCvkgrQFLqGNPR6NjyXx/H1jI32v0+KyWalkkFQRjPcWy4TfotLAm2x
KDpqff7jXKoEdbjKXcXVZhnEu2CuY1RK7P2tzIHM8EEIMXpaN83SKFuvoHYey53VcymJXEYXc4At
gg5ALNJAgey7bOx6kwuk/SqKwtn6uKRVHhdQ3GJKdueaUJwVzAY6Ho21Ha7EGmfVQ6cX0p0Yv9Qo
DjrACnc6fQKoDo4RkpOAfO4GmLTZVi/zAb0F3V9pcn4wcnAjDFQl07OR6Ffwa4KN3JNrKNAJce3B
pMqQqXF0akPyhBOSDO7e+WhHk+z3AV0gFBOkrxVnTY2lA4a3oRn67YLl+79DX+KE0p0FMp62HZmF
IVQV8/oKb1zcjndkU3cLdhGRDLBRXtiFDwFFps3Vlex9k3dvTwO/49yZfGiiy8x4XN9zQfI483XY
YjHPVfNXgcBwmqGc+LB+/xspebeCuX2U5Oc1t/gLBVWnt5WiwS6M/GNyc2nr6VTRE7LmgogPnZUc
lABZC2DHFfblc7lI0QdF/sBmm7yZkXlijMVYzBauc6qf/GurOKZ1Z8oU6tXr0gK/nQs0IF6KsEcX
IIOC43oN4jVolhmAvsnII+10b24hHYOT2AHsr9mCAWCD822xVlNR/t84UwMp03ljoYOF7HifIrvR
BNwyejeHlkDM+byqRNzE6JfeyvEuC9aNIjfPyOH5zHixtwB49MWsqGM6YtKHyvQVlgb/4cvgPgES
uXP1xeQqLEwMvFqo8o2wOJKBAeAAJgnkXmjP96l3BlpwQcEFheyGcQCjXdVlRljxtFeVMvC1Su79
n7XsUQgeb8apciJPK14iYdCdbItCZordoreF4SUu9glY2y14PJ8hur/W67eU33K7ZNJ7smAcRzOL
IXj/TQLUuZZnzDp21RHqZ9PjC2CQQJYic7lNsEGYclvr1/X1TL7Oeh8UPTssjp40MEZQACQ1Uz6X
62fjFzII98v/ViPHbzxYZ2tl3NiAmSlGMqrkTxLGIFYZR6zju+39AsMu3KMiFQ9vDfjx1wszzmR2
Gw04F1k3vfF2AEvd0Z/YO9guJ6nVI7xTYqsztQrFJkTSyDpS9UFc+XQQ3YxMB6DBBbyVzjr023ae
RNiIFtisubiPCEiPoVGHhRMEy3raKTklKFe1ci3YndSaS2ahYUMnXCk0BV5mXwg3R2i5NqKGHwqL
Tnd92sKTCDnaH+PRTM1DNwAczi+tN24b/AfuiuvMJOJB8LNgjvpJqtgUoHF2EqjFtRotKT+MRdGy
lNGLxD7iU9GmD51zgZb0Kt7DYtlsKKf4cf5X7aZ2iIVW2PDbsDP6SfDx7XMSXix0Bz+OnLDAi5D3
9yQQSD1ikRlBa0NsZBFVvhmIkwMSjvmU5hWhL9Ufm8KwqaM6uo/rI50POw7AbxTin2dSMSUEFhEk
uyFLmGapIENSu6B1V59cLq0q7FiBQhLK5ZxkYTQVKwdvN6khhdvWZGtxSqY32LD4GSPM+HDRdAVj
SIOqWy4HXXEL0e2KZ0obLB9DE2F2aCTPGC7OE4qlNsSSyJ4Xo6G1hkiNjxFY880H1IXMfEO7kSdV
HZh0gCmMuwQZcgIN0Ez6hIc4l4U+cfukebDpzbYcFVCR3AUv5EHqEw+IXYs3zpJVvOmH2YFodsZC
cRDGmaOCBQT7eDjcxA1Cgiw858IxsEcVALsVLBmzi7vUv+oWUDqd13Gkkc3jBfXQaiWiLd+RKDKv
b8cWTISZvI3IfbJCsI2ReWRrlYZQYAog0pFZ3lfSQn1NMNtE1twRb3JTLTmW7fCAShl4gcB/9/1P
qyjwtfUoExAcd8At2EnGGTkY54c10FrB2Zs+LigbcfdFhgqZSv1U7qn+jzN3rkfdRiG4jexm0xEH
Mq3JtPcd1YAhomCWfj4nRxsivq7WJ31lPyhuk3j9LRtgiKA26WqcPmvm7a11hZvCa6er9J7tUvaI
ka7IAmLWiJFxAprdJlLsxrgENa1uVguMLrRTtFItfZolW8YmCx4h1fPlbQA7h5VtMO+LTiZpEJLn
f+7BNYxnqO8W4UBOp1G+MFCZB7piK/fr6x5uoEnmqP5WUoFJ8vWhAeum9U6XEtTF+NemJ6g+hWJj
5Z3PvtlyF3R42q9RRegVoV6wdsagT94/3kp84ClvGKExXVXXLuqnUyebGYfmWfrGDRXl54OcY5xE
Im0gEVe4oiydgFRyW3pCkfClmFsvQPxPsMdakvdHYEolA0pjLgWEKcmLeT2/dfRt7SVMaEkBhLJX
8x5XZch69IchjeM+tzwxbkUE1V5jgmooxSsO0G/nuLHo0+uR1bkDULlCPND5jK/TBgARso7023bI
BY9lq5+9j7ssvQm79GT6SBqF+sNktO4AEwUUSCVrBIjXDU1DrZQtEFzRMyH6BsyxssCNMsp6gYje
P8bJpaa3Jw9J8RYXmMYKNTkqUA0iPb4YUVNJErnRP1raGo2dm4ELvl8Dh39Ul+ZSlY5C2xhCBIrz
qHBHNrr/2mp3nqOCkUHd86vn6uhuQKxVbcZMaPc5ITTj4oiiUEa/AOOi/lul0ux1v/dKd6VuwS1V
PccIyFFZqRYloiI/3FPobqLPlpmV64RO2e9XL0DM9PaEjBjBzrwaglHPG9WIar6k9jkJSxxKRpSC
CCvTr3j430W3P6CTLO0Vo2TbMVD3JW2/gzBPWS8xl3BvusGs3B1iVudiD7LketmqQRZ6r5/NYJuG
BPDhlkwKnYSlWoYTU9jKeE/QRS5uPtTwGOCx+iG00fSsQTsGm2UbS2y8SrxWgv/Qcsx/txPBrXOE
k80zVzaMtOVoruXU/1ahv3EN+gxEV3bQdKQzo9oec/4M0ryKr1Coy3XcdPqKVkiZTDwim8QmO+4Z
95/Tb2ikgBES3RJuPTEszn2BBQOcs5jpYfkH5XGL40x/scvVnHBwwbTTxl3IMxbzEnBSsClM5Ily
twKngjuQcQXfl8RhmFAojpkgXbMJmB5IkONv1208oqFZd8JeM2dA4LWvT0MFOPX4PBqAU/aHg4HF
EIP5b0ZJ8kpQkx8LlwkysZAIzPe5dsFLFCetjf+SRS3h8Y3ThNoWET0CSCfZ/kCp51FFvKVFqQeV
gR2faAa21W+2kLjNFbIT5X4gNWju0ZFBkIP9j3WMkMHDZ8ELVQQ8PB6p/8wiDHbAZS6vHSMnQRHA
BHht7gnrjK2U+Yux31brnCduZ9tj8fnd4Am3QQ3EcBTJJGe30RMdNZ9J6Mf+wPDchVSlqxHV2GiB
PGTiOpLrdrMRAPPJZm23RLNiYm0amgy4+SCcMPVUyuluKsnYrUgO4l9+EILK2T546+/hLaK14gVq
u9yvAM2U5QXudQ2ntZYli7vaTxNGzODJ/PO6jBTZvbmH8RUUEW0Gl+T74/azmrYxJHK+Pf8OhvtS
gIVyRnQbmsRLMzKWBYnMoPfWJQyIdTVf/TnPWwhraBEjVIJLB4mO2xof7g8dh4Xse4zsuHgsbNR5
BWFJuo6YFD8m+4r4fGmFbotW8ndM/NsIUDB+JD0Q5s8mkvlm2wvSBXfnRPtUmwWdtrrbTgx6AD1T
NcVIT4y2zUJfjH7rpsb6w/tsBuIDprjMaO4W+S0Fcz7rSS6co4r2cyo9fFzKfI9NnwPOUYzS8yQ1
9UuLisdKylqxlc1p1nJhB9fbmqNFbYctg0RiVPKVqFp1Iaar98MdeBzTGMldl/Wm30qcWQ7rSqmb
DQ8+Xl9Cl7yK60v3tg0DttQaDxs37XGLPGclZLkYNcNE3P1aVqXVPIU/kOOYSubfoYgDcZxTYrdH
kTYseq9S6ywL0xJM+gwfdTcKmbgn41YgMIUlKKaeKgDYHQ1rcUYtQx07PIK5mtbWh4nGxS+uhicz
YXg1Pd/tTaAv/Ib1mFn+emO0Do6xh/3nG/8Lk1XcGMJ2Fo1f19e5lA+SytE4CtdxbTwZ0vLDrybZ
+8EYSA+Ww5ogDGxeGG2JqrNpdn0XPb7QeOwtLBSHA6BtAvTnoEBtj74q7EwCcDeQwns+0ZnEpdMh
1A6c8eIlFB3dduf2kcP4iYVHgXKdnWToAEZg+vBArCrb0YgRtxa9gZ14zYMqfVhgP9G/FvvYgMdF
TS73SnBrHLO3CCRVOQYXDI2v2VsPV/cdsP6l88GJDbzwG626mAvYucSG/vMnkLzSZFvL2ye9hUDJ
XfNWfDPmx+1Upqh4EYSBTI4MLirWTEjjrCAU3CJIVsXjj1qtonB5VamNp4PVKkd6Z3c4uEVn/HsR
9mZDhm7tJLxwV1VP0sGI82564/WWHWnWOa7rRHnwYR8SsnBA3QTEi2GKFUXwE73qffPJjekJnxN0
u9BYuvESosp7YeG2SfNanauxcJxoDeZVv+5H+luIB1tMN3BHSJbyC6a0dilIIjlbkkGbLjjC7Jwq
3uvMnLjrCxd9xGx7w4v0xu5BfCRcN7TZQPW/N6iY1CbJsmfnHi1fIpYnbetIJjyja/O06HxL2iW4
nbBVauX+R+NQlcpeFqau3Xy6cEnEia8Er2YEl4UQoGxkMafsfmx4yu/G/svwkrkix3KXAPXY08cu
ddxPI75Yc09rd5N7wpsFdlkntvI7c9/vOuhn9qURCO5XcAtOPyJL/KAgn5WTILjEIyo51gxARPoB
bLfUzSphV8OZwNTJvJWlIFaiWavfv6/wte7pe1fXy6l05VzyL+9yxVlfS9aFMyxMqWpvc9itdkyl
NxA3Z2EKCbBQONCczN4YZ91Q6eCl+D/KCfAJdIxxRQ1s5UNF4UjNQMdXGSNGCpvuKRpMSLMXdOXN
64sUwOVH/yi1Ymon7MnQDjJDqgbKhoQrT6XlAxQpOK+CjOmC3Jb7ixNn6mi6rFYPse+cvga3bXui
squN+8rnguz3/dnWehMH83nnIlsN4cDQVVv7kf9sXpF5mGgLUG/CF50LcvYZSiwgEPv6ROmxglp7
GYzwDfoNBYeYdwcwWbEEX8jhYGd4BuFFd2n2pU9Na6Gu2Pwgk7u7WKjvWkKT76zUCmMFVcGtjf0u
RvtrdcX1hUC/ARCRIOha15mtntsE9VRsS0pojfa2qQFkRfwpEwQUPs4nGGPJW115JzOnJkPACqr2
d94+N09HxChD+tsp1tdgRc0jVFb2hlDJ0G7ohsg8hAZLmTf/4RzJNlOtNSnDmADytIP/z6G34IFt
lZraiT9vhHLjQltF/MfXTvkAOB3SY97ULeL1kUzpoMp+X5IVRaj/za1A00j2XviT+J7jY+i/ZPyC
b3RvNre5y0MOI6hbdVxOfjKSWqqkzU3WzbSYiOhLV1zW+e+pZncvhf0QOhVLcRJi/T8Ed4WVSXLt
fPp37BYSTKFv0Fi7rrpXaMDx4CHlemGPHvCsBOg+/+p82mVXiYexTcQv18xZI02513R8DVkvawc5
TCLwQ4KIpc9JrcOmMeH4d2IVfdSgv+q9tGj6BThrakCg5N9dpxe7/5V/bOTRBL2J0YBg1YA40sFX
uMjzZW4UHa1k5heM8APgMHnzRSjBlXx67hXMbrSP35TnLjkudORVcZbQZo1i+afYfVv8rxpVY0+C
QQvN9fP9MRmpqL9M6q0LazWhVKntyM853gBGqJ3vNHkHPO2Me313ETpDirvFelS1Glk2d4f/UJ9n
o0/y5045xu5TAhVL3yDEVLR+Sr0KejiUhDuJrUlGVxr+aSs3394Rzc2FRUAGEey3gir1xDCNyIG6
PSJUBlbGzzVmiHFLCmqK5ft8Z3zfafZnaoyJFWysQWxAyMF+Ar4xfrHkyd9f2BdIlqhZ2hcvcdX4
nnbmnHGgWsVMurCkl2Y6VgXpgQ2/BGfLRdEhUPXrnEKGp0lDLmyj3ShA1PayxT5mTnbz1i/Mvbcl
voRONWiEVH0IBbvq1EnUYtrlmB0abVJmccrx4ulaRqnc45Zvl4FeQJgMJAgyEGi9dDAppKKLSkvC
Z63UTjYFO3QDRoWnr1d6j2SN3OWH67Kck8vUrPJe0KnDJp9BSt83QUT3sZehgMT5sD40bcC4vAtS
8zqxKj+irOCfIJEXtjvQreUKvKCDvedEGslVt+X8uPWi8oJHPCJidyuXVrYFh7RpvNpUGspcqlCF
DiZSd9YzCRRibdJchLoLNI65QQzFDmtOyyYcZVmYdw6GJgbiVJCX4DQAc+3JG4wwI9pDZhVRQG5h
9Qsc7Sh/RjoJLuNOXFaKZDIZk91n4PxF0aqhw1CNFOpONGdWt1LLawUSnccTIjBflOYEUVIkjPLk
UbqLZTGU6547oIrcXm+c2SLzMtC9ylaEcnawt4yCajzuJ+Csyjmb6uFvMyeqPX1hmgTy/eoLjDwr
Rif1YPuECDGCL8jfdezoxLlEQDL35GtmcJSxc5XQzHiN+S4fOG3DxemR5uGXiela2QZSLeNiPvd/
1HDedfFN+wBwy/ofPec+QZ+GImjh7fFTcrpFRgpiME+LDHvAtugw7DJR2AZS41dWPir1R3QEudYU
gh1n+B3l6RRFUFCv42yRO8F6sGZY6xq/rADkmTPRm784CWCM6pxw8EroS405oB0VucRni25nvCEl
ih/qxjPSvUsZsCe4u1dFXfHWty0i5UbCjecb66Km5qJXOXzs1TI6k6AJWG9FTFWHFoOzZL5bAQI4
axB3Em7Z9gShezEuMCfY1XXtEdiwX5Ccj2TAaf6cvzezNiQ/IrHzPRWC1s2DbzO1eSFJpOayO11f
bd5ynp8JJsf46TS9wRm6VHi6M6H6ntK6h+X/+y/o/VxyZL7UktROo8kfY5ZlRZcIXTuaI5NVvp1F
cqbeoWEVqU8dfbEdsN6PPk2Jwq5RbHYwtZoPYxu6sCVmGId+wE5RgLFoFlGPxResJRvRPe3eQgTJ
EJUQ1ec57SVWosyJ02D0Z6YAEW+P8zwXG7RBxbmy3tlUqtfhoBS72v27wqjTFmMFwhhm52j9HDSg
bgqkkphBs6nH4klfEcKP5qGlwx8cPJMNGLNn3GYLllAr2u1svNUzvhkY1VkSLXN/g367868r1bRJ
yL13AhVwWT3FmZz074u572Ymws854JIZBkVaPSDfcD0bvJ727eUQWcmWg755qbMKRIgnKmBlPW4P
LM8LfvUGDQ267mW9fb6oxP2gqqw4sonaIYumwvxGAvzKCDmhZ+PB6QP1l8PiAA1pd/l4ZPPPiBSd
HaLp/ccThCyVSeXClgE2yd4C5v5wekb8t5yr88Pn8VGR0/++J7/gB75YuliTohHTIWGIvSlb/AKH
pKpunJ3ESoHlnZOQ9TrlQ1tO14h6BORHJSp0QYN5qvN1/3WB3R5+XUayl9IlBqRX0CI0pUjpMHeE
v1noMozV/3eBhkixFRICTSv3L8+NH0YUvQMtP97UmTZmVWD9XTP490FXZDuuS/hSvLLurYgke/jj
mk9yKseoBS2KlhMY6mDR9AaHL8MWrx0O5WRYsTMK8Or9DsnNBAnitfVjYn52vVEXe8+V5Y91yIdk
yPeI/0jb5cVuXKjY6N/jmH1ndpx7dzB7X9rSW+BN4D/PEB2KcLQ6lkwjGbsIqHcfaNXcZeLSxIyD
LqQt6SY75fz92GlwlqE60oHDq8phW1syJ2Jpej7vk81SCpwv2PnGq2ci6StUMFe/pfHRB7M5e8F1
9Y8qayTnW9HuCDhzcFUEEhD+nfGXJlmLk44PTxzcNBZeWyBufYsUjjfxXwXemqJI3MfIdMfuevrj
D9NzAc4vd3+lsHEreVyNuhwuyth/TEbcffcrkZ6lTGumaTTAIKymQjh+SKcqLNkKqbXUQ4OR/0fI
wEfy5OHkde08Pt9KkZOiQ9OZ8vWxFMInuWfjUe6XXlFI8A1C+vSOnfnD9KHTewPQHdixYuLMhJ9c
n75cQ96LSmjMpMAiyZdKw+xiqNJVOOgd+eBFBIem1InBLH3JG64tnZAmdHcA2mnQPa2nb+VaIuja
vDv+H1tazzcBiupAfPBECj/VGzSQg1c5uSi4QvVXnl7Y9lzQoHhPM0sBWCdMhsHFCbnKBapJ5BCi
cYvANaD47uRD+cw7gyGxoh5ERXM63Z0QSJ+c+NnLO0i5V/eC3oSPfyd3pJ7KXH4FCHbP3u8DtS2+
a4RoACj863luQwIeOyAjKpB9wNAHwa3Zom6/ycfY78KQDGiqcge5VdSkCIhqF99NL6LL58W/hJ9o
ZYnwoNdK/upbiREacp3oyYxNWedfodCv7NoL8mbdkArogYQ5iWQBq/PsPI9xRdGyJyIPHDISesuM
TIBKcakoW9JYa22dqXNXCmmKRCMbxBZya4NFmuAKelUVaQgol3+OALxED9IjsV5+9y3b5JV5panR
jx3KnfMo5xOnLC2ndCbV6HX0hDNr6lPmuZXXKq6Y4id9Cmt11pYpu+2Pee+TUPIp1aIyEqFh3/uk
kjqTkVcE3JoVcIx7pNkkF3Xk2S+gKnO1k6kvpPMsV0wi19vlYL1/2xhmGzRrVCVlsshcJFD2PMyX
9Ox6qQUcHX1ngQJU4vUDxUbfQ2G9KtIA9ocMlwsm0TlvToEc0CCIS3IwxuQztuGmwGOmcJjHfeK1
bwOZLFrrtsiI4dn8GWE7wIlxVe+kjry69tW3OgnbsWqRNzB6Ke4oyItPFlXBCRx0wzqtj9ogNZFV
1NT08X6rq0jYAFulllHsZgiJ73T17waG3viSB7pIphnstifyn25UWWF+i/GlZASiGeRu1Fg5WfFU
FeJV/D1yPqM80WH+wB4CM9fT61btArdFtP8m9zlSXVCRn638V0eGwUNhrZyb1sES2bloFOa3oO1N
bivuOAUFTBMwCKutm1rFIqfE+GsM81fMQmGaAG3khSwhxG3ZDkawTCGmX3PGRIvVoqhhz6nL4X4H
ajqHVMW2cV5nKUmgXOt7iK2Bhx5/r9mRcHdO9QvFtXcYpr1p0nxOFGoo8F6eb9dc2/CpoWK36uGB
4WKqS72gE/EeL72DhPkQ4JGaTaL8NxYDXciIANgfzllyGElcoJRA+T2flcNBrwSFI2cFZ51Iwya6
o+JDZq9UB0b8V5EOcXM6fdEkP2kmy4R9Xy81A77QoKF3CIeAwlBGXHybBu7vS+BrLmtstGVPsocb
YAuYOOMFNvEuuuHYZxsyBD8CHdOU96uExYwn+tSle2gd50N+Z6s1HvbMbcnByG3pl22uIeikrkMm
5HTawkexxl2FIF2v3Ex2W0udt6XdL0iRNLXETbmcgJD14DbGecywVJ6S598LHAHOzf0EiHezo9Hn
ANy9MGubBc8EJeqZg36xqyBfNTIv2vNXFikfX6cDO7jF8Z6KmrBV+KHgfvJxKuIoNMwr+3cur+ct
O5HQ1T4ME1CgqkfM9mRqWg6inCJ5S6e7EbMUc3qXJAIML9avFl1WOHXBXeoR/1cNpCeWM6zBXvLX
AsuRdOs2du2F2bBCL3OpNBfk4yklaUWwMsE5Ny+34YzHbM/txRrPSsKXnM5TYWcRBBP+ma5Mayr4
TB+VvYLGUJGPgrgKCjH6J/GojEzOro1UypwE4rxpl2FD519rlRy/WJvtRtM8y7cBvh0MzibfZQ/L
JUkJ2lAqavNI9tejHiRb+VIUKAr6oRAwfjjwjiEQbGoKmcraSr7B9syda1G0itpy+8NQZzfEm5rj
c/iK+/bWomMdgD+ZTfAKY/alyO92R77UKrvw8KGarWMlT91+GkazWkjr1ocv+XKPfgD4lceSOrvH
UeLSuMyniNM203KoQqzTPw9lUDn5l/Z4gOLYrr3IKXRRjCd1ydCAaofM3cynWx8v6OY5b2fapbLX
uyfAsVyDz45n8zx8VFNx4ffjGvCwbRI2tlZF6WNOuuvdLFKZ4xe3djFYtKLh97Ta/BoheY56tVVr
+i2tzGUhmaoELTPlGcCo2sA9VRAoLb08EHOlLXQt2vahStM3wy23O1h0iugUQ0U71CHaw2meDgxL
b67IGXUpQtUwfFnlm6wogAyGfZK62m3mYvEjjaTtdR+zy6VihtoRpTBQlXJOsr1fp6p724FLSYFN
M11TMMDWWZhSQf19vm9rsE+PCDkZCHG9nH6+M0QQWGeScME//tNSEuBmQ6ZIdnL720E4tYq2ufQr
NFamT5DHJPoysdLvYPucarfAvZ37o2g6TOkLIJTItUGYZLAZaQljSfyLwQYHWbKlx80HR4Gr5onk
Vadk6zOvPC1kHMqaTeCPCLgxZNGXQJ/RXDhoX9SAFRXJgGM1RLeiht1da2jPRePzEGxZqfYciCxy
6LKfkpqIH509pjPnV2q9hgJENc3DSHwaXYLAXZpVgeFH/0A/1THH27KofOYhefRave4aWC+WYpyr
BfLXYZeCoCukRNKKZspx+ILCKAE3bt8qG98etXP9t/v2tjvoisiZmWIKFUnFoXNL/S4chbzNBjj1
YghlO/Y+zoaOlJ5MDBBCdP2kg5TJegfzvGSvJl/54MXlySCARKoFZdth32/TGuimCFfAcyW9UJDL
8xi3ezjiMsxohTldN2+8W+9DY9gYC0yiJrYFg3igWVkkD6fUH+B33ntNoru1Yu7a8MsHfASjGnay
iMGlV/u+s+QRzYyZEoqZQuYLyevvJ7UZI07coS63UxFlQI9vePHiMoq88MYuj0RBkzPPHua35QrG
KNjD2wak3AJQs7KkpgjYsYxha+XuBP6Z88NQuAZnFTThnqe3Mmi5/TCSNn+lzKr+bpaC5WjAoe/2
/Urg20SiRd6hl0/lK8fU4m2kCyU7AxkDN/0kpKEfYnPvNI9/2LHXZOWi0D+YDQOp+HNv63TDO22V
yHo6t7vDxaOUZNn6FT8jjorZU4cGbB53TR7PLbT32yu7mL6LifXmqYYUfO4apuPeLoF6xYB8SOi6
fS8/5+wTL2UZK0qPy56zJ5KKL+QiYw4oK7p05Gt6jBDytMAxkx3y0My2LVyQ2WenPcFzcftueXHS
3Hcy3r1k1pr7g7jUoih8o8mGaxQwRJYQPXVqIAPgNr8duUMgPUR3r1UV6VW7RdW9sox/KtcUaqLk
DdAGwTi+IDpY6LSfK/WmLLLksR6kbRfQUvYZwi/neQ7cYxYmBrFXhUHn1MVChQTSRJOLDo8YfmSE
vc9sNe1cqfNWUjk1AYlyJcanalVR9SmtL0CDnlfvx7/6azF2rFM4VlwP7+h8Nzq2JZdrNE8TOET/
RcaA3xxocvePB1yL7cZfZZY9r607AullS8f2QjgZdKVKJKJqZPRa5E8JqFbftfH6iT6EZUHXiSFY
tRpBwiLgLvS1k8+0t3jbERGPtnmvwYI6lMzq3ieJCRQv8JxLvrTq/55LdpjG+8toJS6g3iJcdVV7
SEI1z9ZgRZPn0w0y3Tay6eb7IoHnqPNgfSFdqFqvImxQIrHwGMX0IiGbHAqMWv7hQBLkEYFltwNy
FZr/E1m3LcGvqciHrr5CPPdcvcsY3Aqr0l3wxwpMi+sA13vU6I5nlV+DnqifP+HvZgEG4ZMro6rt
MMst25PzmFplX2CDcjKjT3sUhzAXu/cIvIXDMFeLFeuLKQmZ6AuqrHPHngEeA2uPjiDpoCILLQTS
glxoPlYfr5QbgoTd375gJNLV/TIbovznXEf07VHgceYWWYIfq4/OQXXfKmkQQelvf1rZhxdozwbP
cdn+y6h5NczXdcYVss3yzffYtjMW9jRg3JxLkOEYpQCceLDqpZXOpDILeVZErrW2cGKKuQOOmj1K
y26nD/VZoM9rqKqwKT+xtPaBl/Tt7UmAegf4WZ0aSPhF+kBVJv5CYWsdC+9CsqQ0QJYYEaEllowV
ZBjTjELpl3Rct0vQxsSOXnHQ2I6gmsN94/Han9O/t/5BiKoX3TiDps3L1R1u4z1yJ2livLoduwkB
PNMVX2/F8W/qMeh8e026bNBdbJh0+qO1EJ7V8dOemrmutTTL27erkAyH3DVSlWcQQsWcs3ZwwXRD
BiLdRgBhKLF9Aa/wBpoemU51qXZZ/KVFVsE0H6ujqgiduxWIRTMUha5xyavZt8xHPP5Z7csSqXBG
Z7iGaFhLvszHOPGv9ESGuGF1t+r40YltHTK/f+mdWJHK45fi9SVMYJSsImqfxSkzxk+ZYxDoR9XW
V8Z7TyyGzLYw8+mTY4paywrTD/K9xTNH/BRbplDjzqvYgpdgkF63EU7sRxujT4wZQMqK90MLcNgg
1syB25MQJgdJ57K6dKn2fU/y+mUfSDTJKEKyAm28sR9MHygbXtRvXrbFMg2COacrE2bwHugxnPSn
HzCxjrsmEcaJLv3UvCuskgdKN6K6CdDqNY7MPsYgKxc76DowRCZsOXWHc6wzr/HDEyBwhro5NQCi
mlZ0/+wlhxCLa/ftHs+vYiNumdj3ANOdcxOYCm0gy27WZnxt0Sn2CpF69QNpcIPJ7I2egwrdwSSd
SZWGbHEoF5ER3R5nwuYAPPOzCz4y5RekarruKVhVmSpGWYDe8i3os7OyyYfHKHodQtoQmXPDJhH+
18catfmo1WZzfCUv3EnGWxYnFZ3CJbHebjUC1VhUGEXhK/VEH2U8rZnHTJsPfY44L4m24UCj4FB8
PXxMRqwYqM98abylLlVko434tTtfTf387DnpdeTWEXaS3L+EXt1X6IEua4UHNcJBAUNTOsyNlsvS
/WvKX1o7wobxsClxhcUrgt6osy5HXQf1w1t+4JUstTWr6ZqjvK+y6z+Bt0zKLjYoDfnzfoUE2W0n
2ucm1SXtJiwXHaFGrmop1SfabHtotEVy8/J0aSV1xTgD4pZs4G6mdYEQLaA9XsLATy7sWvWqHH5p
tDvJ9ML+M0v2rArd7+JcFTnwEF3kGSP6sN0wiCwU6mpZgk3EGGfZZm9RrBhZSLX5QzY92EI8UvzL
d6jDtVJSaohrt95x3eClM9p9fx8YzVhqbLXKq8ndO4Xq+BiuarT+eKU5e2jmrGYaZNeFFfh6dmeJ
jhnXhw5NFs8mgB+soLqHg4O/YmeeQYwnn2s9mCoBcBcIOSTD14e/ULYEA8BgkTmko4dHyr4pQL6+
sV5y0VqXpWhNNqNeGoxZFiqZoBH4AiMZxRHvrmd6TfxMrSph0WIB34ac9Wlwp+pZiu57MoEplWHz
ZKDh7eqPUsmJQu1/3wt0YIQIRy7S2JfCKImyyJOOlxP/5Liua3MvmKZYLhhSJ7MMLL7oEhsul0Y6
rMXwg5Ufqs9ODiX/oBwJunteoBZkDa2BHiIDAQlewGOqRt6k77LpBZLI3zFZhwPq7Gi38SA/rnny
FZWxxUpUOJ7HNQdp0tsQ0G3GIliPDJWWqzokOkCSZXLXlcxPelQ8gmFHudSjmTZ2E0hojJHsMmGJ
mQEHFsj/w2nisQ/jF0tGZBdfq5XR2H4It7Q+CsxQjBSHa6QiPxu0bTaP8l29yKL78YeF2IWD6zzT
mw8+XhWyVc6GxMVC+hpQi6Ladc+osN5Qg146dN9Bh1ZGeTUOS5n3skFL/17sZksrBmX/18u/A+E9
7m7RZ9Gc31yXtvtqWY+UTsNlt2bw8nNxcI7aBuZ1tYcbeVVYS3hXHJBfPT/3CLx0u70p7t+RVNEB
t5flLK7HQAgs/3EkrEk0Q8l/5PUEiXNqiCqImtfKtC/mUmUMAQoBFHGMQ0tpZASHpWGty2PqBrNe
hP7Ll4XYzQRh4R4Tu1f+fq7INbZLCBgcwq2Y7QS/qwWSUgdlqo9KqUrYptd0KBPocbIjmvz3QKDh
2rGySSCGIqInWEMyvPRG9ggzyQWwNB3kYKn4oUhv182oWSvtsYlJBwgjjCof3uPcTkfqcwWHdoyw
RJNpiztzkukFz+hSNnPt2RYMJRhM5vwJS2i5y0YYZ11Qt2kOZWf6opjk/+BxtCQSLMzJWczKTLQF
Am2gyVYm+j54hDBqwgQrLJqyewhNBUdob0bwUWF0ENXhDhp3epfrCLRROsXUruKeWHk2NA5cf9w+
LF950uH0ShptEOkPuHR/TNocUXOzRggh7a2WKlogdnvReWyIo8czbDc6asWAbUsPNJqzO0VGP04b
feu8g3hgLnRgFZYsutyRgYyuyV2cnbNN3feNusXD1HFsa+Obn8lsOq4WE8ym9PCt79HjvfVd6+nu
0rEZoAAnKrJXfiPmX2OkVDokqO48eohDPoeHwg4EvTNi8SQq5T1rhXGCDQxMSJQg3ysBd/xeAUQF
8JCMPtncjiJQUrxNEtXToNCqLD5UYniYFc/LNk46MzS2SO5+wiuA2mPaUUJv6gi7HCsiJx3p43Zw
dXnQlOIG243NKD0mc05sn9lfd/Waprh4r0YT1GVHovhaoLTPDIPiljnFCw/RHWsjCw7fQdk5icx6
y6qYeYA3rmlcjQfWL30Bgp82pxzBkQxku+8zAE5bjfhQf6rEAjuKgVvFi6uErlUr/TeZHcEgmTYD
b4cMVswkKX7gODP/7Ojwh6A5N3eUQ7LZ6oFre0nOE1fWhcWgoQy9GXcOEmJZysdtmKrX6S3DGq8n
GHNjp932GmTmp4/CDWkHfp2/G5NmIBsruNo4N3HopBxKH0iACWCm0B9YRkQugnw+pDzh/H0Ks+1U
wuYVXOWGXpQKqxkC6YzaSqXMXitylA3lDKqKiCYEAfpwo+rEU2nNgA1xOBI77jSjq1un5ubQ1rxo
jkH/4KpcsO5EquOvEGiohfOxu8if+JeyUHqJ9oZWx0faC6X9rdy3JWhr49QMrIHDJ5uhS8Xdtj0M
ZcggmBmXUgjON5FGIjmlmcE/eqwq87aNqbC5pPoIJsuauSqUlIcGI1beyHqlZkZM3ycURR/+73JC
pUenUmDRdnkBtIPF2YEz6wL4zk5JnYoJqbUpDwF84AjxmZgasDPuXSoe8v9fJigFPhujwRtoLJr0
fdjoynfwdbeOR/Jk3xqumkVkD+sRewfoDX8vJGfawBeQFLG7+RTYvl28X3mYPfhSFvkaBFjoMJb+
VDQ1i0ZHiIb9UaxBZdbNyCGA0ha7E+XPdsyQ8p7mJkl+/CnX2qeMaMtyI1gEbYlVvailFxajBITe
+/MKfcuj2SZtHfTdAOpOi+NTBSl9XrmH2aT8vhXPN+00pGWI5d72Ku70hSGWRDiXWj4xSQQ0ozI7
A60mL7YN62oJejsBn6MRqfnP4h2uT3vcJccy5pdUkYqyRCKC4iw2LNd5bfVzQko2cxy3nYXXsXMc
fo/J/cVl7Mlrv3WxOEVUnYNFl93C8Z/tsxVVQZdseVf3ZemGSrkc0hZpp+87uZ33R2f7Qb+aZC1t
bHIWgZy+bOXsluw48Iym9xIL9XsZiNtUGLOjgXOg4PRQVbWDFkwFBbXsIbodxTvcZd2GwBp0K2vZ
lNW77e+ytgIkJ7lskwWfcEj8FZyyzNO/qiAbHYjEqMUP+3C4wEF9jw7LoSPFf93NRKAbXKaCz+Sc
R9ffyCl8q86hc62Spp3Q/bhXo48KcrT8So+drd++sLYKW1df4YBn0GybtpsBdvVrcmqd3l0eIU1e
LyFifAxuLbU8gnFTN2F1KH206C3N3cmGNcGo4HURTl8rJqNjNqAHEA+uSBA7ue6jC9Kg5EMh9yU2
wYu/NcCLqeUDssSvkImmDwtP9ryY1XLKu9AcIW7rnKE8LCp1cOwIu5pv3/7ZyJQyxOoxO8ZTTBGz
NJM3+ZHHj6UPXT4x7kL+0KzVzeqejlFwOUZ/GgmhPqvgCeqrpfQqAJONz52IjeOtvywqJws2cvbM
QQhcUUYqm/HElikSvnh23EUABNWQmAUrfW6OlwN25OPzfTUlQ7Og7XEmW1ATs2Kn+ggWlOULhwqt
eAB0yJwfDTIvl8CWLCW0LcGoUuaU1mnefOIvHvo6bwE5vC+tL8N4+u65NMYGGrdvC1fEg462a3D1
P2wPOO4afUPC/BNIpU6R+Y7zACEtuRfkbw+nI/Nf6Cy7TppOHgdM1utrZYdSG1Njs2QMG70wzrLb
pzKBgE/A0aqnW1seaz7D8B+lWgVDbrA6p6mXk3ypvyz6kGaVPkY2jSjNNICje4G+8xRSnU+ibmzt
uQgM/ZGC6gjsSlKWPRE74WDWUs0SRLUwzRKdrzXTREaKw1Me45nLX2dn858rFRU9J8ObCtlJnUm0
BaB/4oXktgzeao/bkFQve3qnD3oMjQ1yObN4Cyl6SM6NdXSZ1DsQh853X3KRazwVrsr5FjP8SXzQ
ZCrEZZYYhgn+5T9J9MUCVUjb1q9zeY2qxs7sUVTAehk50ElKFU8PM5upUNfY97tlszIhngoh00PY
ED4fAMzpp+PgoFgWWd1qUjjzbNfKPOq8bkS9XgtNnsaWfYGQvO+0nLzAwWUkD6FqvF5Xky7FmO/O
th98zR5zvjgu5Ixa6c5RVTEiEIiys1T7WO5enqH1SEqGrZjphMBkZOhLSJoGMjvGes2w+OoJ9CNz
YpWiDgFz51OwFaVk2sxi3Uh3pDx27T/Mt/fqn33E6drZ2AVb/KSXK/HdyPc5W77vyGWWpoIIWgIX
M+MSfSr+JiOIIbgau/IxiycGNJ8fya9cZkpTXH2VuTZb+aUFigz/+KJDtVzVD4hBbgG2xvczj/AJ
6UMypnmBDDiCQ5t2vRx98+jk8LDSdj4kuFSc18dw/I31wHkGg+dekghgQOCjXhcZwHNAe0PbMwq4
WeDduo89vFEPaoGS7uc7shgjkEmI2zYvn7AoSo7yZAyYVVWKzpgAG2EfT6Q3nNeyaDnWcASDmTUp
aANcbjx7TN8AFCvk+PWiPO9vFyGrh64qR7yjk19lnATlT0n62rK+Bz4/DAjEyiMl2BM16SZ/wLR/
pLcTpDz6suRNBFH1WkRnte5EV2n4D0ww+IoU/raxGjrfvJ2o4Hb9VJTghGh4bIGLRR9u2R70hjdt
dSxWip30P4+cJMHM62spkbfvkzjd5rvSLrwXZrVyS34WNhhdFvTcXhbzaFy/JuJsTuhOGref0n4R
QPQVmHnrDOq+rzZ9zljkm9t8tAt/XwWtt/VXmSXPenQsz4XT7inCqgN4J3RBuLMXXccS3fO96gLO
UZZ/UHjB9+iAT6lRUNGztO6uAi31t5QY1BdYd7yccJPMluzynV3r4Q5dN7P58goTWzDFXZxlTdkM
L87qOSAMNODZImuPSRHl5fl+l3mv4X5/GkdrP/IiLeE4FMVIykJUWS+1JARo9BIAsU+6uaGTyNxI
Guo0PVxExklpJwDRgD2bQcS/nDUNwq2QOfM/FNX3kCt6vFY84r2ztHsQTyoiLvgM00sv69ekABgU
llMrvW040s+mItD1l4AeX/Te7eiev/aVgBkM+OaEKvBYCuUJgKxK3rtfhh3aqJHaXvzzt7ILiatE
rqTKgDBevOJdHu4RoipjCrGAGS6eV36mHT5Ntsvm1XyovKJ8btVFzd8vU2Lc+dJBQRe32EMjpIml
k7cQY8nQJQCuiP/TPtdaN1gtYbFhIwZH+9IqrWUUiiG2c10xoZI43391St1ItqDIlq3wbETGEsWe
tUwvsTS5vb4Nz3ZME7bCxq3SCYBi/T4YugJBh3h40Ftak0taBe8AdV+LeTWBQJGYuFcaVFzLJ2gA
TsgWnswTlAyth0Akleyc+MB14BKDR91rKt18cpMhhjhx0pBSddqYkf6vk4hn4k92pmqAvIZRRXNC
uS2f23Qzwp61WENabIZxaLg46MiajTEZvoMw7a6zZeOi4RIwmwE6lFUv1gZ4VJyfeO874IklLL/P
30SknoNxB4IgozVNfHJeCnYyQKhyPTp3cTt3/92/yeORBYXYiMFNp5SqgxtCJemahE4H3OrphARP
KdsPj+lweoyE46IVwnckflEguj7w4lxLwe707SbLAITXGs3tztuxUlWAI3kS7AaQOiWtJGYB7B2G
aQtuCIxWJ8hNPG0+xb13PUMOiq9wq6hpFkvdeAd/XUgG5q943+CiJUsm2jwd+KEBhjB8GdKASfEt
d9Fq8RfgiLDwR5FgO6f54RdRKCDOEjSIksf4RayGf5BUTys9zEWY0So9N6iIEtZQmknr30dytGei
thA5WfCNMx5yTimyqcjGbsRzjXkUitsvmp9oYiiNMGzYxqb8pvFINoY2pqUGkQMZzmgikrRsNBuE
Yda1lSLuFU8zXZA5K2lME++1fLr5G1OBA5QoyhqK890dh2NOsdXcOctjDISpNHxVn0huTqPKylkr
88SfbwAhAY936X8Fh2uMA8+JPwc+hs4mGRIikFjPGZVj5QdJ6ilOKvzO8c8fg23zqxAxY3eCihCz
aWOoKgS/Qqnn7pFGoQn62voYeXG2G3ODlOu2t7JQtQP1V3xrFeMMrkEd780fpH/9sYdmQgDP37IC
Exw3iEcGJH3CMV9sTU5SIJfmOzHcH0fHBb5CXtn0xN2gA7T2U5dj1TfbCtgIbwKIn0DVBaMU+eNc
Onr/kU8ZPlJN3Gd1okdujAujAUejJ7T6K/Jz0MpbHyHFZsozZ9Zy7yGXe0rwpHeCfGjO9VgTtJju
2MgVsyIPBATMqwlKi1j01C7VqOJPd85OzNg4sOHDbzGNwF7OPXZuzCwo4O+xYzodRJU+G4d2Ymwu
V7WFDLNPMI9AbkX61vbZLwOAFWHSfz5GUyzaCiZxFJ0dRDYEguQjzkGmwcijGbRVG74VFwGFsNZE
RPPxyE/ANm+hwwaGXkwW+Gc3uWGO7HaqgBVgdJc2ECgcA06jFELxLgU6saTMErjtMAzt4P7yhr6U
AMtFh/rc9+PKOsyqVSPyuU2NaXLMNXkraO9Y/7rrnzG10Gc1wEp5zlKPUXesZ8tQQq8ALUkjK0gc
jg6WNy2UBIO8blusCT28GxfrMICCVqqqOnHnZXxf65I3SRO7BT0dKOY77/i4CKzV0kzxLvUn8cC3
SS5wAy84JUcjRFUYMNQz38Z/kKOxLLRrk6B1v3uDkyO1q2z33VpZXw8ReueKIY3dbRVGLUsH63ls
gaXvSZDkRhmdGVbQNuaF3PX2E/XwooB1lAqw7YxjX0jKmkEPXwr7fXGFUzPq6RFAH8r4QhQcHrPQ
b11YFLl/r//4wMD7bZnm18KoU9SJWWCLs5ZTmObe5r3cjcumrak2vZt7L7KtDx6oes3TpAvm0ZQe
N0qwm/QHnq56hnkb4o7LilmI7XDKO+LfjLCussoRJQfIs8okiZRforQ1QnrDuKBmKjo/9ByQeM2r
7CipWUsCDdUcsqkP7halPS3aTkZ4m0J0+gpUgn4m2lUtU+qGbwkPCG+llaK+thmgjTlSih1A+ANe
iRPfFIBt68kql+jDANK4GSpy+MKiJ7zYYRcZRfEsj/xcMU4k1NNEbJHdEUpg5uKk0IsiHAaKHLbF
DzKnEnnrptuazEyxC2BBJoib5/58swyLOIIETFel0xn9soCocBzp4WcPG2gT3JnJ6uK2nhdyE8YF
NoRNZYrR1md7Iq6L7CmTJfRlv2oKTr7a+u+le1HMIUYPUpZFO/X7Jd4h9mApQ533LD+XKjNH+mYG
og9QmqIvnuRxzZHc5McXlTNuLds59qpCe40j8uyw+Kl1G+AltWng94CQkS1cFxBTWCJtkH47LdPX
NmRRj529ndImZBGEXLm7E/lT/458T/ZT2vjYHFAQBJt81+/wSXw3OBq22gISA1taTEa9wyL4fN8f
j7x83yAlJ78zheOiaq74EVtARUej7MWVDaBUoHy6HO3rEIARPPtCEKydHBrf6JjUQEzHstzpHfPi
UZm2vyPec8fOhu6cQUxbsDGqTcatVq6Mzyb+kgUMWmGqGB1syDW4GgoTdVF4LnHOrLltK/AYfus2
qT7cGl5vNkhbAuk60AjIGrl8trijUUq+6MjIopn7pPP4yRuuTfIF2lLp56PM69vNWGKk+iU2h+Cb
TFkacVbNWqnsstOpIBrUQ/phRChTguMwGeBnIgT6Q9ZMBp79rQeKAmtpLAg3lllPDCS1RBSm5s3C
bQGODUsrrRqV+nfLN26K8+IaNHB+xk9zJCJ9+ntwaaJstKGf7UALu7gcntF0usp2SdLyfoVklxDM
ZlUfBakhJJ97tInbTUa4eDJay/YttvN/1nDNYAIYWSq6vnwj5EGlOfOv9ZfU7QMwMMwEzJ3CTUls
cMWTdzi7LePrCatVGjEVh8cKbjy7oDaVmtd5PbeI/gELqURz/66sjnZaSmfcIwOYY3gCSEA0HyD2
0x0so8M+N1QPTOdJcwfQic1Qe4FV9JvJ72OOg+U3qRT+F3Zzxj/Jf6/Bo/3n/JxElN4BOh/GnqhU
5EZ21jkN6FbRSieyWAHk7X2UtyxjzcZol2zvLov7cG5DRemID7eB+fNJPfcDQlXOyIpBaJVpvywX
MItVJCmR8noUKPgATPwleBwRa3EakH9Skq++GmQbThBOO3WI8SNK2GWuBVGN0Dqu7YVmJ9UHc+3t
PhfA02FoeHNrX0EGq9MoIt9rSGXb2umUtPGUTu++/S/gtuN9mjxaBH7ndPmQkYg6fYjoqWkNoL3T
or9pSioy/7SfT0rFGMR5SBM4Y+YVbWCT2/WA2/DCeLAGSgzTmWGS2bWmApaNtA5aALsFii34xOe1
uZgFEC++OTDUDl0Tt96UEu0jcvNh4JtJKmdG+9k9qkp39mZSrwIBqJA3kYgOXuuL2ICdYuRC46Mr
Z4wM6Aq9qkUPOZDmnX7rx5CwORgsrr9UW0w2eCaH9QRtHO1X9sMn96j/YqxGJjBnl/qQAOy04xDK
0hz+zKsGFsmo/QY6jHW0erEM4wBMksu/SDDhWS9xKvG5PhBRTJv8W6oRqLCAYCoC5c3wZWFtxgN7
i3agEEjlF5Mum87Dw6J658I15HSkCwO4TdeaBBOIlddHMJppPCW2d95ocJ4vqNRVLnqHKa7KPZV2
b8o4egqXa9wqo8SLdkVwPaonAsOIXb8nlD/Ftu+hBAwNMuqaC5fsViF2NvwBz6n27txe0LIYDkUJ
eDD84vC5hzJOJW602z6gML7LbTPBnqXWnMmYn0NplSmX7dK+vsX2jLvJeicMVlLvN0bGXCHxRiff
/l4ALjMUbFkAXJ1iEFUhYuPAn6olF7n5TGUjEPF9f5FbS5UQTSMNu7oz35aQUShDab4yvldEJycf
TiDpgHA58BOtEDs7tKaItGb3EAhowcqzGMfeDWst7hlt7wzuHQTERbm3tBdNuMyjmiOfm6V46dkC
TW3G558u4Yn+Li6dkr69pEITC35p40fusQTiOqtnR494I4Veyd0GebMRs9RowMWFnX5/uJ+ROkBy
Qu/6qcSdsWfRZawX1UuW0ziYQjgf2ZSYlH+mGsNhojRHNaubJRuNv/bzBQR/fpqN8sXPydYjj31w
5x+XUieFDtnYsw2lmql8i9CmDiU+rufuaMXsU1Pl95zEykeQAJGikOWCYttiH5/xC182kNU5/Smd
DB/avvjRMUAM62fEqkGD/eskex6zv6jIQruf4a6VB6YXQ/JEz5wPBKPXkjRqMoqBHberwcZY/BMv
yBY0Q2aFo0dQnIz3/Y22Lxg96kIw3c42mKgb9b1H82KLNhfmwkXM+PFE0pMVRW8DXLoOFC/h+X+n
UrK0oPA/wUOS1VJjBFmkSVRol/pZrNCAKTnj2aoIopKHrGJji0h6S2HYsJ2LRBn4AE/sU3y1IsPn
ayYU57yd+wKFPIcf+Q9MAHKyjenfUHLaksMPL81XE68PdwS3fcZFB5vIpIRbQr+ZaCaCXtKguO8y
XXOM3MbIpKU0kJR0bRR8MCCtKoUstunD5XqpGjk/SNZk3EmaL1PKzDUxYsz/ie6IF59OkvTB/kKz
5oHLcLDhzFNONV01BE9KXKLMh+xSBSJ8r+iEdpW4kl+gEDFqIn8hxrbxWmmyHv+Con7zuvQHR8LW
P1sXgq34t4+QzJTFkqYS3wwCCk5rgeKgvT/2YhuLxq+Pi9tiHiq+WXgcFBRelCID4DpJI3kAopdK
54dUxe+ucWpULMHQkLAhowdrwdK0wsEz02owKROXw6WghOTUHXm4ihZmnft9GL6Tz22CdIAxSQ6l
ySxwujrI2S3u0D/G95qpVy4GGUBydyptKHF9xLR1HFb42XW/R3b55UBQR1C7G9QAejsQYs83LKJc
lod8u5dBL8WYBYbYzJ1TwzFdJcvBHYlcauhKMZ6vuA/L1wEpXHoKIvXIwjsdVvxy/TBT5/VuVXfg
0FnIeGiGF2yKZYzKh7js0OoNma/tTI0JtJULKkiky4CLAQoMouGYd9nh7LA+OCsSyJENFfPLPJN8
JJwXuqqtX2l8Wp5TIPf/nuQVTHzTxZ7qeWMz5MRMLUzoiX+fytNJfd/MWuxutz/SFuzy4Rb1KHTI
DT3f5VJ+oXudm7V9DBNXMg3pT3mDZQD7J79IItyb9nBA3yeFuWFPUYEeYlSwclk+AUZkDHFC49am
JRTSc7QjoGZMeFNiCpF8rqLKwxkG+hug2a1Slzyb6F8QURDWD69kPHgj8BLAkxLIs+RX+VWv12Ok
nq1QZEN/l7ywly//x8XoSsk/BoJ6yUvb9R3zNf6r1AQ6pfjElzw3FeUihzf5nMMW7Is5JqmMZA4P
5Aj6CV3M7PyqfB3mOqsdh4ga3aBW5QGddHt71mth6dpAWbqxrPPXzga2sD/w5ZEbXIbzK+f03vR5
8pVul+SULfHjFO8E4u9CXucMdOlSXnBuuonphAJzaVBMXHcpd9A5uuKdWUk5tt6ZqJ+KBQMuxKfA
5UbhkgH+FdejTnh7+7yqjSyjBdPyQhYokHerznn5bwSoeccHppKKRv8oYU2Hp8G8EhYSFOloa0A6
5gWNtVDN/FZN9GJWd58nanCyy8m8xkNQPE8Gbs87AzirkRjxpB/RqijfF07YxyI3+LpFssCIVTv3
Yz01AA0YI0Vn8MK6Cx3vhJ89YaYb0PimSACKYSQJvJgly8nIFpwbKGCjDeF/vEWmCWQZASh9t/04
MoJWE+qgZx1aTXvDBVKnWwJ9LpG/EQJ1RRzixcTpXOkcBbm8sBXg7yrcZFV+ydnuAxMuU+ybewPM
48GcnZg2Ho7fvbAOZokaLDt2mszTTnjWI6m0WwS0JzFFblJc2FZJNcdUeEmFqEtT5WRBpvlo1VPS
mVfN0uM2uNQFL8IDyU57DLB+fZSjNsP7MCymPa9gvoMsvAemlAjMlFbPAAeWw0K93amdvQvzubSI
jaRLuE4SHAonN/K0oypbiMAx97DN9zBA4lzLODtKjteL00mSISAqXu0Z21D0VX6eU8p1e3bKpQyn
eTV2Qh1/tg3u+05P3sWhXjMk7VA+IMExWEMr+XtT9wW2IRjJ6THG+P4vpVFzhFkRX+9yqYu6tIKT
h9OANj9Ju89yaCsqNqJ9pXnPbUehj4cQaTPtX9kb+9uRsyejX2Yls7zqRRUM4AI0Py+DDBve6wxY
1SWYuYZpWux96qObtfzF/gl2EXkoxzjToyCeqbwFEAxPEopQqU2PjwEFQS3mnpE9+tDvzl4x44qW
6WnPo0lO7y7PdOgVI+qOm3pr1eoD+z1kTpulBAVF76F0zdvEgzy2wE9cVDcaJsI6LCyh6QaAcqTp
HceX4JjTnlTK0zJITeeF6zsmfuVK5DV0MBN3Sho5C57fFywtluZtbLpP/HYUovLiAVBslS+uzO0t
YNyReOQ9xOrOQd40BBKkHqydJsG4HJ6shqw+PZG7QwnUferiUVuveWctfuS9TjgjTFHgYn42gpOI
idDTosh+fJdpJuC9lSnhEF8lfklzcU6qALchdpGjb8kc5mD+Vhvsx7H77I3CKP93wVoIIKthbaXP
BHwZx5jp2v6fpEaNSOlwS2tyHJtvsov0CfTx3CKkPdAI2HWveA941uKnDJhhFBmbvGKDGgMsxoNo
d5HsshS12puTggdjqOmKpb7TWrAR+k96S7wvXlnI2dpm7k4/3EX/K+9OLjK36qItOroqJeDTCkCJ
mWZkUjUJEOY1tKgEiKjF6mWUDJqhJhLbSWPwlU8e1ouXrLEHqddZJJpZGkaR2ZBRn5ngwaHnOiY9
VboWjqx0Q/oXLXppF7Rsts8yaXv5zmESTyt+ClnZmbAXMyfvosnw1UAh1acN0SaT7wNiuJwp7EE8
36OME3UbVw5uBdnJ880Je4aQMlWYowfwyrnYUL3u+YvDMAbf/W6suMxkXWL/pYDuM0ddGXCZKlvB
CXmH1oKn1l/JvlanUxyz0OpUkrDlasbdWIhGZ4PE9K1gxU1gOTy2nc20jtetQAcC91zlYFnnpqLP
jMoIKylMIy48+frAtris3vxxZdgpShSWc7dnTupZzNFNmqhRkE08S7nujRu73KtL6QBZVdujhl8U
LbgnjKXUl1TozJX2D4dcUUlj5Oh1oRJmUzFj5yTeceOQ96p+FBIdIamc33v2kor10apnq1zBMg0c
fbFsy9uiVeXJdyYHgTvTL8Oo9ILJWtiQYqCLntfGulowf1WDy7I/wbQGLOgIrLJrmkd9DuDP9RSz
V9MgL6o+j8QRk1HV5onHUVs+7bKawrUWIkVfx1Wr7pK6L+FkomZQgkUPemoyA4VwHUtnRR6dG3kd
b7q504+6Nrr+Hfa14PlOWLBq//ph/HKLQF7Hnh2KiuR0KCBo9WCnpsSLsnjHwUg365L1sNk+h8k/
6ZR8EkYl+gfj5cW5VHUmDg0CQoUKiLGG1nGZC13cTwwvI7vUrgLRQsKTuljq/CZInLXXzQ0fAkSe
BqUPDjAjdhtYqFSdwRnSdBvFefWD8Qtp65yzv6w2laooEWkIZGJm5a9tMxhosjnIkaWlLRA2+gd9
4ri7Qo+I79ox9XSD239ZTdP6Yxw5fLwike82NNmpBRTCX6+1RdbJU13fMrix4ylMxSVJ41kbj3cx
oeBs3AaKiz45OiYUN9rMvOadZZIlU1KWG4sej7J9mxtxlVntv5/GMq/Pdn+L14OxeYvCAe9oEpUL
68DCGZ1r2/TcZKFTXMOjk/IkPi1VYjJyYB3I0okftnWTDmsoI3Bh2pyePELsRy6yOEXa+y1dwXH1
UhdQafA4WSLjsf6m4zrjgkbDAHUyklvBvVWXJRcXsr4q5dK3Fo+ttTVE3xcWgJqE7IcAFa6H87Mf
4Iz7WdgYtJy3HSH4rJGbBgShJoAWQZ4IGkCI7TCbBY2Z3lb4KP4h01d4dcrOGNYLsv2HmCMf0gaD
3YR50OvWbYHC5kYzEKKjhUoEEfe3/L+kEWPhqAn6iMzDCYKHy/gWvd+0TzIiSrTBd8z4HAqnu4vJ
hCuS+DZiwYbHNEzV4b7pZ8P3xx3S+EXAQ6IScbWo8gy9E8K/v5qEwu0yD6z+u3ekuATIupg6E4vR
xbbvrj13MeL66EDvtRZkoqXlzbCHUxNgcdfqCMff709+O1XwgMt4tz/Y9p/T3EEB/BZzCcum9Vkz
ugNjN3+U8K91MrSQDQDR9tl3tTGTj/jPSUNM+6vV7/Ow2P/aYaXs/m55/YHOI8eVPUcILxDuIDbD
MbkJlnW6mSmFlSekm7QS90utn+8mAPNhZlibOLhOqpuGa8LZ6nJHkUHbovlBqB7TR3Y3lLqqKUUS
AOz1EQBjR+0/mC/Lf9XL8OIa64cgEhXrlQyeDuYxPa1RfzopeQy5aY+RQTGo6lnRLscwe/VS50VM
jvn7+d9o+1188UgL/tkmFkVf1qPori2Twcg2pZGKKCoavtm/UrfEW8Jq8bE3dPg4JKOvunokw148
g+JhHgfFBSc8ZMLqjE+N6zhiukLs+cICaJ8RJ007NrFoIW2Hob9ujq5F5egtZp6xL9s1t/h7BgA2
1Bjp+M8ODGcQWCkhxMtbqWnDceahqp4N+N9/O7C9D0ckfMe9FipGUPXpfgoiY8Nj0suEpV2HlW28
br2jPShIs9x3P6Zy2bK/UOeIGMhrP66Qp9H7hJce9VDDnf3tzLnh/Pz4t2sOage1DCo/GBoNVGrF
tGh0U7YKZ24GbAM/D5iJvBL1qMYZrUihWuncVdgAI+sgfqm0KBlu6bqhAZb32Vw/zdROPVanE1hS
/wW1Ub/HZ5MpN+hNAUioEIfoEeOrFgx1027F8Kg6pYNIPkWesWcs4cC+2cHU1BcIDRXxaXrHBRIN
t6VErAroATrZsj4Q7LLeMStFvlv0nycs7Avwg31/l6fbjMwcqaYpGSxtkfUUeqF2tw3kCO3gbkkw
JRyekNf10wKeOxvQSgtRxu6g8F7J5NuFA0sKxy/Fe+h+ywAqI/S+VWuxJTDtFVL0Udo6H4yl8rwK
Wpce+/3h/Kx8ILezHYlCuHadQQExcLCX/KVx0rg0f9iPZlOAHK2G05wykRXfQmvwrV9H5TNTXfK5
ALD+NEKR0znIjV51hm9YhgLo8pSLoGNdU1L6Kzc+xM5HsTkaHo3Qu3LWijM+fF/HX65xDRoWK+9P
Rt9xQVmsyJN948kR0YX1IfmhuJZsf15tfAIqqL1t2KehAiBRJVTjbFue4dpVjKrH0xHEbAF8KcF3
GDqNs2Siw5l+yXzLRd8PUFBtEh6EU2gQb5flRjti0jvX9auaG835AQd8Itc1bF2h5VgF+MmCX8K7
lZbOSpR2cKPAa8fSdQU2BbMCYlS8DKwiJzc2NPYWhQ/XQvv81THMCma7WSj2w2l7TtsjDoDzfN1T
6yUYwF5PEgWm72CNpJGTh1Ws+JWlAi0DV4Opsa3YaYrOaAotHoqZGV85RuzGe26hH8AUwTOsERKH
6dktU/wf9T/eh6FMQJg9NgniYSQ5I/YTBND1amQwG8svu19DdtIcOEw1zuXbRdrHezZ1TlAL5nm1
vTgVg6aQDUYRCZRA4q+npeUM1pVSTfBsdE0ME/bj7cRJ3YTE9Jt2O5S8pOvdouSiJNSLL4F7Peqw
zMkY+EbFJ8pD3FRBeNQw/+pBrWOG+zYgrNc5YvYEgmZ5/barxcZijKYQayhj2MIdcM5lvD4+sGF9
q5cUca22uSsyS1QiIX8UxQYGBWMPzU9c2h9+y1JcWKE/c4cEyd+CA0S0RQOmiCF4us70yZLaXkvj
IulESNdLyBpJ2iZSqHo8NaOXVAIN1J3FUO4/PAlcoPXq9UKPGmKb9dI3vOR7lp2tgQdwZtVEohtV
nlxwPtGCU6apkNWYeF5PFxnD1iNznjsxIMdiYyhhFidcTyb8XmLNXYkT05QB+vCJqzJqpXYKRLUa
lault9Nhzd9tqmQVQdhDjSKTocIHkbYuxpMIe+UfMJhh/TuIzJEsW6Sc1B/h2zEWjN9FFo/U0akB
IKLHrPPGjMMjQdFJXi0urVcwocNAMpthdQNMCRDVG14+cl4FeHiR/H4uyK8JbnjpZdYdZL1GFBal
DVXcAZRvvierTPYa6cxtcmGCZY0+sojsxRRx9wHliwrbJ+k6F4aXk/NX/agIWJw0Ijn3YNVp2zfb
47UNfJGGzlzOEDHXbYdrkvdYGHrtkwNmAcZXkstN3gzVaetdJCLetHiwTz+iTFXK0QZ1JwnpTFH4
VbuK6ZenpQfQYa7p56y1G0mX1zPO/mGYgH5oUJxvuASiEPryPJUmECMW4vm03VRuaBnfPmb4hCuK
NGIGMspW6yX+mcnLBfeFdXnV1IrFLIznUISNq7OXdq5y9GZ5g1Zz3BIMpWOvcdxo6lJ6Dqqkisfc
0VXk6r26Dmt4erJobiPwrRnWZ/k2GderOLeYIPBuJGkrYMXSn0kfMiJBvhStAZ2Htzo0cMtmCm4I
PcYa0CewZvM4tViBnoalz0wmaCWLQRsuLOBBhK78DpEuHzsK5Uv4Af9fDzfL9sUWcDshAXd/nBbu
orXVlyXxRnREfHuO9SSKw4zLDRch+sDx2hooFtztYPPcvwmCV08joZ+DBhnq3Ndej6CgQgeKVtVP
L8V79xyksLDE/gKw9Bd0JAdXtvSSpVbUBKvfTwzAOyZr/H2TFqRG+YYJzNzxQInpRIUMv+kWM5Aj
WXMFTevE91ZXA8wIZpn5ev/WFpeM8pglcKjqQnjOjVuVarfO21piSIFUWG1OIw/d+aPTh7/QeOCT
Xe22uo2XHRFgdqPobucBT/nEfDmaDWKEn72KOtLmI7F/nZLvBb+C0kBi8CtOGtYHSRzUxoid7KFC
k11mqK6LJlNrvZ9MjR3Vvg6VHmr85jrVlUIMgKIzoDCOqwZpsc9MiV9elxuzIDAZXra9UXsGlaKS
Er8NM27bOuUeDT6f0ikXN0wzbg+F+fTE15R3VHJmFd0TbPr2chZvR7eDuXoyUxIcJ7Cgw1hZuL1B
EUwUFSfNOUtRnonKxfpj413QMUcxuGonnUlmp/Nmf9rZDywX19zPCHtoJApN5s2twxhipBCzX0n7
Qf9oaWQrIdFrTD0uSsm92iMQjmt/zbykDLqVnBQrbPJ+KEQLOlUcO9TQboVk9SWuC2y/5XWOHOsR
Zqmdx/er0VFz/KUvw8fwi55xZNORTuOd+sWbsj0KpoVtECNMxaTeGPy236Ji81SBxLiIhmlK3opa
/wwriMO+e9f+vkYqs1obNXqvRiRHiWoSFpXpuffMx8rf2PfWYFCP4l0W9jNBPgVJF6mnd0lfJ3oO
JXkDgbA49M/SkYE54S9J2jxeX1uIYZghRor0FilV/RePA7nAUQgSdD2xqTjyUR/bv8gZMsyNBwJz
ge/YoL+dhuW0EUwqw/FK1bKMLgekgSpPB3Zo5g00ZfPQ9ZR/VP6htPaTxJ3uUTc4zFU7AKqyYZ3w
co8y/yNFvHYIyQ66nkC4+BZ8rGN0BPPR0JGRrMnxoFba9ZEJvIJHFO5fRpcsYeW1EdD5WQW8cEcU
D51GymJdKgh1sydEtZsAwNly/78VSNdZu200qvOcQB+Ikjj2vzPRQB+ze/HDhPRbhRbL2g6F+1pj
MFk5lRnatkQ78AnjZZ5muqIEkHie9afsPj1zfaMRxjbDUD8ifxyj+6vbgMihy8XSIZCVuR+z7DZG
G14f0Ccbx7QpEOFo/cF6LvaYQAdIE4deq8azzqKM8+CLGDT3ijfCjlX28WUn3n43tdYPo1qHuj+K
LZpqXLE/o7yMfNBdKk87gpOso/PfM64L4Xi4fY0O7FxTWm0kEXHcuTqEp6abHejlKG8UJYM8tJNF
FSgXLeugk3s0ePKZEMlAkk9mezT11m/b4FGnglR88aOGKs7VpvmTcGT1H4yGKTR6SSOQIUuQKSC2
BH6xPVgx9as/fDK7kAWb+AEOrS4zjW5DgxVjSHnYeJxGBQZcdyfVLUzKDQ2I5vmO9DeKHEEzxc55
XmMO/sr6xdp/M60XrBQu4m0CdqeIezTeChhGjNwW4Hac1faT/dx9X4M/iDwYNYth2ON1mHpe//Pf
m/Gk5SKStxV21lP+9JIYOjNdJrEiuacypZkjT8CAF89+OR4+xj57oHQKI8xHi/IVK85jyb6o23W9
bcwYgnEyrpr90IMXEAT4LjZNXolki81oszfvJlyvvIKohwGlS0C/g69YuONa4qckD2DbbBACnxm0
RDLmrfUlFYm4aOIXqmK4Jnuv3UVNaN7HMr7XcbHpyo910FwVRht7uurr6sdN6ponKx6JGJl/tFGf
uPkytAvOI/6CySTpte/70Dk7g4jQr0Z2ZlEI4EM1xumLGwizmT7wtmZjrOqC/MJizUnzmmpO9nn2
tMg9z0FwZgTs2t7BpZOZtlToG+fLrMvSYQ26FDDs1MFyj+yOJ4MJmYRDz4EuQKw4j7bWx9OrxtEl
VRp1bOjgt9mbStSQrfyOj7aW1N2T3Dk3LDX2SA2I1HkSTVjQABhr8e4V0dyoGa80aPcYaY41EzrY
R/xaeIfHmjJZPrXh/hQAtwG95p411N+aU6nzwTwvaPjfqk+pzYklSpx6aNIfPtNUTK51uK8VR1as
+AtdTPPrUqD4OgiMdaB4yGAt3itBb9Fw2w982uz0bc0qVPRPwUPk+OpLiJRS+Jp8GFi/F3JOsyku
dHKuVVhd9rkGHGfo+VpZL0JaQQPK/3YEBIW31+7MyQfef439ItJ41j/qoEdgYLpJLYV8HaPHiTLi
lpeNE0prkwTUSsFGu/D0isRg2+wsQsaECBPNzx+cQwzF6SeVRXUY9CCnBdhNm7L5sVlzIWcdFjwe
KbHPurl2PekQtTJd1+f2Vy6SZP1RiH3ZZJESVibGB7hml6mpcEPfRQ4pZbn1CZrhKA/vCvBHs/Ib
Cr+lCCdmKqKnnp+AVv+OOryXsejT7KZTxUuNd1XWkdBZzjHXuzoCBgtt//+/GSWRSUfR9j63yjyJ
7DotN4cbBHoQWcpJh4xLqej3eH9NvtyH/et62cO1AjOdCuYoZnQSPCMOSXCVQkj3VIbDK1TiTaHZ
lqYEEq8L0Atuoh0fHF60JdMKRsxsCWgVz6gXVMaOfBaKNqTq3mMoyPsbmztA9SgqcJWMtTcC8dn1
I9q4dLXBCPHQSHsZUdPWZNkgblwmfQk/uPiuYHV4POUnMLMbDXv4snyVr7h4dMmA92GpjF3iKgqB
mZF9AUCiGZ/G8AxuRzEI/r/hxA1C+DQGm3DW+xcqzTD2aR8Ru6Ng/6s7bMrbiM/iv3Ub+nntJUXX
ZSxNH8c2CBoXeVxN2LMMj7FUOv+SNQ9nO6MLRomjKznEaOjFx4/4try2lzDF1VqIT+FZP7UpEEvH
5h/2qyw3EIQwu9pYIT1BscoYa5oQDF/2BjgtW7jnPPT5h9/XytahU3vmxTj57egMfUzA4zWyE/8k
Y2PQFcT7HzgmUlUckNvz52W5TEmyQWwuDUxmF5FojKMrBb6qRlOUFvfFrbvBVXThFPkoLKGx3gN6
h7/Ay+VwTV+q3HfU8kieVmgUvOBWFHDDFNQddpxAyMoB4f4cAeRJkoG/pw+ofnx20S4rJdCSi2V2
YJ7ahj3PFDxCKQOL1rldioQdWTPB7uw5rPp6kIlgQJ3ONd2FwcZPsX5nPNDdAV1KW0JRUjTMCM0m
z3p0TQN4PEGC1qAPTByCkTJiUvYCr+AZzXYC5xRZTLMyGTgx/TT5vrZfRBPuw5U2R91g/HLzR5l9
tcRAbMLIkg2H/DF3JeHwrAsDApyBFYkhFUZ3Rx6mdYoGx0pXdfUTToukRH6iie+Tch5YLIYNR7OO
FNlh/9Nph0MHTka2rrEHuZy3ReocjpNThgBzq0sstCycxffmobyKpQgYRdaoRzCLcCvME8vXB5/Z
GoarTG6fC3YcQsiYWbYLdIf9zjpj+2ocNU/3wEtf1uow8dZP3l3Q0Zs72sVuW8ex/it09aTGisMF
zMyBz/FkyFsBDsqsInGRQZK6WNoiUmDFHaX96OZd2OROChUl8gGJ9MYZCxRNHw9IlryFbmk8A709
G39NuaSWdLub+G60kdYIjNQl1shnTyEQ31n6BSAXecD9hJ99MBI/Y1t9q7ZXyz9t6hg+uPo7y/d2
XfZGKcVCkR4qWlFVNJp2SLLUQjRDjUdaFzmDA/BBRgY2BI4mrmE/dxDRMvhqBx1tIqWzzqTfrZTF
sWqLCwbd7tFuB0ID143dT+R7DWt3Yg5y5h178XQHICiysz4BEVDF+jT0nGBhEKzTN7+RDVnM+QDE
pbGFtSKR/zIXA3do10RBsVktSncSO3dYRpP5csYF6ZguTgq7OUa3BLDdg3MyQJg699LL8DsBnyZa
mzlYi0EhChHQcf7ZYT7hb5bEnKHe+6Nx5PXsMKVwwlfm7vnkWaIqkOyYpLYDfAlUcdN1d/kuVMg2
vQ+o/EIzYNkFOJFtFAjZClbknOdTIoAmb0+G/Hk4C/WBjfeencdiSTMYV5xolbR0ILwHceRyr9/2
AtJqLhpFfpnfAlUNkI9eUK7F/d1DmgiZz0sc3GmCTtpHbkHdipoPHsJL2X1nqqFJAxjdSLYV0qEF
VkZwl9EclkOWTLKQvt7UTTYECYg4W8vP7TvpGw6O4ro/rt4NKLwFjhcsh4APFvHyWgI/owf25ul5
nubba5SvDdYxJ/kUV7zuMV7L/AB1wAKqBbcIQ3G7ldRDPb1QPM2UAhYTHFQphs/tVkVNlxCAdWck
irckme8rvVn2MXybEHycyA1mGnofSfupNJCWsbgA2dUckl2YDKh+7VdyU8xHZgneYXfnlbygMfoC
vTpS+Oe/DaFF7ApYf5bV1V5ct3wG4mhaZOEOpQuWS/xuMYRlFXthXQ6/wPGYMUgV2DZEqE5SGFYq
WVcANrYgZ/7NrdKqZV/VHgoZ0FYpgB9zUr+7cO39e5ivVlwRKlPp5VST4PrZsuL9mXD335mlQJ6q
bvtYVzRANEx9lzedh+OzBhvuUBsa0+oIS4pc07GCLEaTm7YRexac+tNPVK3BNoTlvmBDiuTKu80Z
eSvo0ltjQT1OUV++9vUl2ghMp+73XOquB5HQski+sdyvXwxjGNt358HqhjSrU+/QbwdiyNM6wG1I
ngqYe6oTpxGqqD9FHvBsLUUGyBeLD9U3nifmI+fq6OxEOyZGDF1HP3TZUoOvhCtZsSa2pfe/JbgV
Vmlhg6i4sIxkd3EWeDyLamI4Tu/iRHXTa0IgKmcTLjziNT7dcF9O47t0Lp3Qao6Jp0jJgWAOfj5g
rgA2HTf4JJLkHG7r9WYkb7zQbfXLxSAMZCG2dsgX+1SVmanmoTLwH6tkrXyzByTK4tG5oslBGECI
nowCfKM7zY7GAC9aHPtGyYzqakGvBloi+NLEjHVVTNUgDHuySos9rXUzQblyv6a8bLNvG2nprVch
5UP+2Z3nBxMqLjWjmje3HgUfEmK2aXjQXXavjVgdjRXFdduvpdnOCb0CRP9Mnjjwi4uVyNFlyWhQ
u9+8XlZb3Z1vVMJ3QWkQ3P/0BNb0NPh02Z8xfPcnP3HA5V7C6oFoqrEkHzHXVxnipYlCyz53Em/d
CRr04NWxIjyDaPyb9W3Rzd4h/H+RgPIxmQSHgn0sXvhmYivNuMTeDTAp6V4NXVNeiZbGZju4B8dc
xgNqxjF/akAZ+/5szw8Uke1KIrMkgaiinS8TviR2AbJpFiLYJkJNf8fdXdjAEOCezDJpO0mWm/HH
rjIs1vr02l04bje6AT9gVwYZosmfIvynB/N/3ZIl/BBX1rCpj3ggvXpIP6lP77Hz8zqnY9WXaW3J
wxDJ1R8ieZOzDd3P6sGV16pCfsLK02BBLGG205vHUNJ11bbuvtqLD+OmwrfhUwAS0OL+WP0sJshS
6Uov1wzowcrTD6k9qw7z+vDkEChs8zvqrMoI96aXwrxlFrFXK4MP1sBvrh0Wq2BTE9Ijq2zjJMYZ
CE6hV8Qb8Z6V0rJD29G4p7CLshFXerXAvE60DD5QWxbCzGzH7Uar2rLL18wKlDy5HpEhZZgaEKNB
7gDGUf3pgYbPmhsz+XYshcc2zZrBtOO8+k2TnVMFrkr/cbyVvBJ2IXjTX1Zk4DgwDH8dcEOuYd1R
PDaoFN5BaSiJ2VRwY5AoNWmTcHKEM4rh5517RNnze8QRxvgMfggSYEwlevtnBnQqVsv5AM/tzA5z
hNSCBy2Qxarvt9TTee8IZaVnmhtNOS0iZIbyO4cynm5drCwRIp8jck7M1thjMaZf5TUO5s+Lu+It
RzlrF2CeGTaW/agPW98UH+ncpKFLqv1vC30BFEY5ub/NEV08LO3zCc3aawywpug4yk2AYtHyGbKB
iWzmmtK35pWSl4dkEbVInMeLNszsGKNHKHSSLOaWhKDoXGdEsmhEJI34DYPz5YrTfyMVMAB8Vuei
UKmk7Yg+p3W2dV01crxVqY2K48BH+RnhtkPeqWvvUkzESFRTZijnjiwQMRXOzmvLD/dH+hdBO1J8
Hik0ormuZCKTeO7T31BtqCteI6l8kZW7NP2MQs9nruFBCBoSK3VWhLIy7oRptpqjhUBgxsyLjCyi
fue6VAAQMU29Ye0ZkUN6sJ5e8ulwzM173DtE4uw5NMAA4zjZeIf+cB0LU3MULoYtxfhBFZmOUHyp
KpJAkLcNF51c6H2yxsNmdgAck+pUeZgV/e73WC4dFsrXs+pqJ6ZBNlkR9a3/mNxFYB588cLutjMD
58JjIZh2rTGbbhwGppajpsXbjhGDDBdHm8yJcAIc9xw2b8EC6kY7dHSk3DmkfS3+dE1a50oAw61V
mo1+5v6IBHq53pCQ82yVmrGDnGYIwmVEpO6yLy0qOsZGHGwgpfGNsELk8R+nbCX7mzDekZlgKMP4
PKWBufGuxbz9oY2Azd7NO/xKqOPrxEoLVlpcX+e+JRBAJV760j3x6sb+QilwtXRfGdkWMqETeNN+
yqovCnmY37c0AGb7p7mKg6mvJVD3b5Kf9jTMwQ1xfE03dDMx7YlxxbB7hdQhu3oLnr+pK12lkKAv
zF8kLlWUulUxIlBN8gAUr+HcZ97LPU4djLa1GitsmCPttinO3opRKT8WHN6V+TsuxzzfF38fIakO
TYlaofA1V+WaT0UlsoXGTxSFBzFcbKa65WDuJa7rIeHVn1kt/lb+ona102pU6RM4gPJwDcNQJ7IO
97DA03YKsVSd3jADrJEmY7yjk7ZSPGER0bFPgdcElG80quRtYz6WtZ7g6+TcyCNbx72O9I+n8HUH
9YHkVK5qp5084hN+ZqVonLUGpiJ3/hpjt3mjH6/XEUdwVWEWZnjTfD0TyicO84jMfqnTmURW9YpL
ahYWrD50c7hLcSu16DAaNnneRDpzezv7TWL5PvoAs4R0i9GqTSIqJSjzjDj4FWUpnRWC/rAfMTsP
viNdR7bo8T44P4fRpr7O46EXAOuHoKRVFcGTYJd2yi6rWiVWatrPYHAjVvoQSOkKw9DOMOG60dKO
t9DPBZgpSNV86U/5bx9+lYx+mkhg4SbZrP8yYafOYHjecxDdM0gT4+Bdm9PxsLV+KOCjuxcgADF2
cTNh/LE2InEa1NoxcNvDDruY4nACf7w6PehDdwsnSp/0lZfVEnXcjB4IWs2di46FDJeqCN2emz1W
0KaGDkDKMH5m1/5KzcNS9s0UylE6iY+grGeg4YCcez99UzcZ1bVAu1YRjIbSr/79bjW9YqXs8jOR
r4Es0JrhwcLTIYOD9V4NUsHdaUAIsONqUyqvyn5OqMTr9a38jyCjylnR3bH/AwrAPOoNJxJcZii0
AwjYgVZE3aSUrIxqJGjhDGMFyu/EmYIqbXl1AfNePjDIStaticUQAGCAJGUpYdf+DHVwyXo49aMB
DprYKAwSqg/LTrfzMHe31NbGfpsGy7TO/6aoTHHrF7AZHa83Oh3HkiCgFnEAfWzkFJ5fEl3jmInU
Rh3uM2mbQSC0exjGRvUstOA7yDLN/Ngj3kDALzEswpizOhDbCu8bkDwCNWLlXQVhr6wtP9gFCN3V
gndp0JNhAEg2yWRVKfKxwxSzBmhtlOQCX4NRlzLO9BZDx87bm3xD3LmWu/XJja8xjOfjrfXRfje0
YsaSHkuE6qPPLOQsf7zx72VRiWP6k2QH4iYW6HjCTs5puW9uJYD1/J+pC+J5cu9coyK7FATBIlqD
yV+RLy39KdWscd9EsllUe3z6CxMFkRu9XeVJb9iRLLlfJVtwtBH15v9P5U0rOWsIcUVeWlscFRKI
qVCRx33FQFJMhGaYd+GqeLDWqjql0uA1gtkwKmn6DaSffTVkhSAT4+rRzPoDZpU7by7UXrLO2ecL
8dZd0EkmLPE80X+oOPsdxk0ZRGD5imp/l7WL8uj6qp+P+182aL5jZHZ9HffFx+qrCIsqVKLIv8Sk
zNX9PDDR6Z8xdOzGONvJCsqY/TYxVfa6D9cSX/tnzkSTiurWJS67CV8ZTfBhowmUmuN/1VV5PTx6
G/HUkNM0uAN9On+w5U3V5qVKGqCOit/lC8DEXQoDW1jE/70+aND/dR75yL5Sx84Q5lhrGLXNZr6k
p9xROk1wC6U0dKaTjI1crEZmktHjjPH9WPsoH70W4+4xgULO/AebSpFiSNi7xCSSTvzYyys/B7rj
uCQ/TZxUw/WIdfrA6M5uRQ5LQWvEMLNtwYQygJBEDsZrg4H0fYV5V4FnUpDRCLIgsFYemKBGoQ+x
coNMeA74vL/0FvuZq+Lb7TDcPTCWTTVzwYB0x7jvmcf5llgfog0c3xx6SVdm7Cv9iOXfDS6L2ffP
u28BiAVguYd83O59d86XJv9Gl4Ou/QzNQLW4FTMbQfOSUhhYbdVFAq7ghBm5V6x4pWg2CKa+NSuo
ivaG6aNTm5fnwVsIR3zW16hapgskLMUtTb1zCrs3AonQ6AdAIH9rhXu5/bbIlJ4CL2DtAmrBNUjL
UaisfxZd/r5+K79gf72RKGJINUUc2ZWmt5nLQxgAK4Zf7BkPlUsTTqmaz1lVcGg9+Gi/b+ZmC7YL
7lQXuZ7FZewaKlgFUqzJQf2qmHhEE+WaytcF8jcO4BygAIT29Ov9YNskX0OO7X7jccZBKmoQ/G+s
i2RqSGJP72F+4ZQxhUMn72GiXyuF1EhuEgEMuhuFxyduEm//XifJXo4G85rkPtbBXeEQPkIXO8lE
gHKSYgsvk8aZuIvyLtvEhPBX7B+8x7bMgfmnEy8IJFM4xnt5CE4kxUIDVFkr/sMEWXsh7oQo5Q/E
jrHD/uyEQaIgMUbFETRJNT2GqGzAu54OHpHUUcxGDzecXd4s8GSHoR5blYpFaOhM/u1yTS3nUSSy
+vEoa/wCGmxtli5qmrjeKxsdWtO9xgRB+zLJEXjrTuj5C1mKTlv4DzxkHI83L33j99OlpiBzDqwL
D1uT8XnYediAj8h9wWn6ntJjUkZR6kK2tcTJkc/EF527URmCJK6Xmkp4HD6aCbpafwh2mPrpaHXK
BhLOl0y5C7AfBG0JKOxocn4DfZVx1fSI/jQF5T1l3BivJz7LqMFfgKYwRgys0TrSKfCSMx6ZrYxz
d0uuqM+SbVpWh+SLyUbzzM+auVUYdellxLnS5BO/4OPspFJAmrsmE51p6sGarlBe9PEw/8ri1Bgj
UPha0zhfVSjADttWPMmWKJKyjwiKBPz9Bp3KhuaMywCM3/PoX8s44x4O4A48KlO3PyQGgquyfENw
/5dwkGAS3Erm95BM2MvAli9NBRe+CfUcpSAah0+kXuSEJdK4O6inI0si9dQbBY4uAsPCtf6XdGp1
Qik5sXrmhH+sgolndWITXi/0fXBrL1QytgoxFmkue4XUWH4ESU5KTd/ENqO30lINH2hEaMSBghyw
jahJJdc3bQfpaeskGXDzgJUC9pBBgYHy8EyaLenuAzeQjtxC44f/KQBx5Q7495oJebWWpUR3n2fm
szmxq2XaWI8uz0WfXbXRfCjUS/U/Jq2cI8Je5N0HGWzCTEVwDtlgbIrFGSin8BbzFIipkZklOr+x
ygVG7/f4oESHLhD9I5uvOMK5rnE4dai3QJPkWTvc3xU3lrAGQgHRGTKLtpinX+VDBtHd1+58DGLc
5LWsg9O2QCNog8XJ7mk3PobfXpI1jVaPEbXzoq6Hc+jKnTYYn1/qY4cWHF0nYhSXinSE/WpkLAKR
HyragntD0kcMEQJP2DIv1y6zbm7Xih7Me0p+BzElykQPxWdkNZQAzPpBcawJnHcqtSdyQEPXcLYL
UkTh8IJZyJAgz0oqmg2X9GQIspk3uwec1pV+KMMhrJjgxkfvwx+l09YHLDu2dgpT4ppYuyPi1Bow
Qh1QfDT9b+K3sn8qZM8FZC7K9OpPt5WzH3yel7otVcHukB5hLN5azwLX6vtrOpZvEYvcPKxVFs1k
B4PEWLcYTXJ/wvBa1Dn+0fAud3m/hIB0ZMk0M68dPsO6jgKBkKcKsTkVr6VFrAp9he+SlVHwNHiF
+aAMz7FxviWeU2r5q4T0CxA9qxH8AgUru1qtK2MRGJbEqQDSQPnxXbNHrtxVlQvywMXk/pxhEtqj
huVm9krLKA9GR2mS67IZh/yDyMcu3KFWsa5nQhONuMdpYrqkA81qVhXhsdXY0G//zXWsHlrC/2ck
O1ievIhHrqohe2GJvIVsXXA4cQWN9NsZ95/ltr1IRGM8Wor9ss6YUon3+AECu11qgacLmFZACnMl
W+laMNl/xb/LDObP8tNKWdZoKUFSUebo00OdEvRPOO/RNmeGw0laNj7gwIPDSBdG1xcPLTXZP8/y
GzaQiYQPdx1vZurNe4g3w+ogjFYlryHhenjEouwS8zo1KXvpuIkbnSgtxoaWBHFvaI6bV3bldVRg
gPfSFXwGpa5oR/8UiUGzej+BhDXj8O6+jKi0XTAtmFk+0YDDCYN0omkNxXAZ0y6obBV0zdfQd0No
S5dZCxYsbX1YCQfb/tmNTJP6KJhSHUsiPZRqutE5TUM3kZZByBc92o5oRnjjLrzoSo4hDJFP63/R
ImTJ3OrOfDknYyY0ZTSWIt4tKIxjsvcjZCSjN1V0bAXWReitm96Duda9fRb7sCY8UfVDfFG+Js4F
ps77EBqC8gq/kdsujCpYuKvr+cO13qISORoP6pplWO8bG7wm6VXPDnntQ0c9V8Q+rdNw19lkjCJF
QG7qQcyifB1Dt0DmNiiW9hZRtGlXYsFA3pnsTsiJMuV2O9qaxkD6Q/Ndgg0uYpg6Dz1hOf0KdXxt
NJc/wRAU8W5Efc5pHbb88xceQFmshyrfXeEDgKm7SdcqEYx502Ah+2c34vYrVegPyI0862fg9r1+
4CcDgCcPcQe/Wg25IGw/n+vwXPeTGZLIt4DZXm0g986a36tapxoj72uee5x4e55DN2I9rc769UiC
LZsumQniDwDiMmUwq6Nof2FuRMn1pcBiPtsczFYb1lxsgle3S851ObeZDYrF9PtTFMsEmsVoATQM
aZ/5kiVo0NeU/YjMD2Z4b6LlN40KIpQjg3iQuu/PFOvmd2q9mViGUG+WCBNzHO5YgmU4BJrhz/d9
XKhZUSdpDLe+lfjO9Xt3hJXW1LpGUJicx+56nz9qd6m+/LjTXH+iZDEI9UrrVloC/ztO+3U6mZoj
TnpyNo3UO8N0WMcAEtFkJBjHESnagsV+0TcBbGz65lkMu2g2kPZkmJ3IG1AXvQI8aDioisOiz54I
MDwp/DnpLol8GMH4g5xTzT9GQcos0NhAycWwt4E2LzL8wp9w5vvNZOVccYt4bJPoysY6oJKuf4eT
HgC5e+LAGrVxImXgsqjsWoN7kFJuC7zt1EbskUWqfBCMo1gpyKeUkFNVdm3vzjxjZ76DwCKdrCyU
CHHDnRioSPyFfWK7jL7HDixudZNHZhkBUiNd5wAFClKIXVem5hz2Wuowoc/9mXvskImoMQTXJyg1
xWYzL2GVsRw2Dd1VCsizs7RJpx9lEN9o2FDl8/deuP/YHoNKLFofFWn+WKqzIhVu3MRwSfGy/qH9
0ax120MmPq6upqtAYR9YfXy4/IaOlURXkIKr0DY3rzO5Y/5IoS//gBsEL/RnuX01zgjWXk9bHiCy
KxCJz2QB1+QlI1VyTHTcPzzs+vCT8FMUe5iRBxaBo4ExEsStuJrVzfJhKgMAgiUL2suwgUo/Xe0a
kV2NfCXTuJUt0QEYzTt+8MKtpgmOSLFdLJG1P/jOlGU3kQIUUL3FbTIo8toimMOe7TGOW/5BPp6a
Zr00XS88xvAwlyTLGAJ3XLExWSW+VNWPluJBwZ1W4tp8vaTHtOweslFLMVLFt0l+ac3Oga1955kn
f7X4ufSLOwnGc0TOqi1OcJKrjI7i+TFErSGmj3xjrdwP05/MYcOHypBSjnS4lCOO3yGv48pTCj3Z
jt5x0gT6VNGQ2iCp3zbHIASv6tjsRk8SHVUrqB3oVkE3T0gxpE7MNk8Q1CT9dNzLLsekfUZoM9j9
B8Cd/9bl4jHBuQJmtjFl08bAAQt/3IaSlArF5IlZ5tzMQ+3JBGPjV+NColzDKHzKtgqhT7/GtHg8
cRZCEKqT61ui+f4T7XR45c4ZHGS1hm0EKeyv6q8hKASbb13TnVXsX44tGTU+wLzuwipiJxuSq7VG
7Wz2QmJMVfFx3HDL0g3wQGyZl8bjk93HfmhYxGyTHeTPp+Xty/IILL2toB5d720ppYfPmEOuLv6M
C2xMpRRQBtiFBXarr36uSZ0Mv34qIiNWAAdhKGzxeImnGoHWRqFNCZ/6D3Q86uL2vw9I68PMT1IF
WUU46rModU/Do4+8uK43piOhSqfbyDAm8j8tDWV2ZMH0wa3xqKrko3UMoG1Naw/dLuoFIsm6ICQk
q20iywKMQHHv7a4hoTRyCFLQqskPg6/w7Roe1y5btG6DhnT8nh/3O6aMleOEYtIHWN0TCMPxhWq8
Wej+rLMW4soqInzDFKvBvE80GDUCYDeJ3NZa4+wsdD7LJXOlyWh4EZi8x4bzOeNuRrblp5fuYpiB
aLbN3aPnRboHbFuvIwA+VvPE1dbdKZ3F/mEnXtkxPU0gxnS9fZB2RMCsQObhbf4jlhet9d/b9ncx
ZGy/GizU/IanIMNeOIJuJlJW9sybXQ9NEBMbTkIwOiND5sRy9Xk0pKWAJ+J2qNwCe0TDvveFkeS+
mF3DNxkfV+bofZ/jmYoacyIoRlkhhjZ5RlHZSt3K3qowVEINFItaajn0ns4S1sryX9cTJpw1IH3Y
ztGyZlxIzqBgLpQqA1BMPOJwUfqdgAV/CPJyDSEEtwszjD9fvEARwD74+n3ZeIJxxzs4QTovArwD
HspwRvhpyLZKVTJ2XmObR42bvTzkfEF+VcMfBlcYTNf/GwMc+4RBc5hZsOtdDlvQgi0w9fm3CnkH
2eNfnBQ9IpydZnylMgIGveHHfb65mxSw4My/cJ/KltpazF20tW7s/SS7gga+NTSi6DIkb6xXlSON
3cj6BDgUQvk+aNXImjTKXauGEymuywRH1/6EBNOkRoU1cQpfu7swYDnUTxZ7DakiZNEcl305V0J6
x2REHOP+iMiS7q2R3r29Df92DRevU86SABoCCkNXbgg8DFpknOcgJ2V0KxPzltHFuDU8wXqqDDso
bnxKgkN29CrXLvYr1wi2JyckyyOLSHKDPMdXsFXoTTPzPD53jAXcx37sHEf8dl6cGyI2b9P5hI9g
E18mLuAo1Tu0GNnxYF5TzXosrptHorsby8+0HQXe9DdlD6PHdlLVpgVLWCIp+aySzXYMultk7keA
jGhZ/ccSCoD6eKHfePPZr4CoocMsIt7qdkvd9uFsz/7TcGbTRnyJu2eAfFh/YkT5gmKb8tS7j0FO
uMSPQj8gBdYhwvHEh++bIVCI016u0jAXnVc/5FqnOfSO7mQ/UfRsAmWuh5ERV9JlgRv81LXCktdK
tzkp7CWcqF9J/UlaNwFykZw+gAELVlhQDgGI59fbpVbCxkSJoFzQo4OBSJyoxhzhzuwXCimwyK1g
IB2copNGA6yxlsE9xuQMdLITrFznvxbgZSKfxD5bvlkDMfyH62KUGH/dftJCYQIFmUP+rzl0shV1
igGRzRiZ/cteSAw/bkcWKywWS9EewxdqsBGuuZdt/KUXDx3o01Ul2R0IuR8kvJnfYlCpPJSCRQiK
2GcJ1YagOAwy4hdUKwpRbOQDZ5fJL1aYRLTnK0c2z4YBALg1S6rLAhRpf8BD9VEj7N1izo7S4Xvu
jQeIooYZhPL6BhK13JupjQg+dw1Kg5mQLv0ExIapHzPtHKO8ntQu+O99yxlrlu71tG5lGkKGuRw7
zNfXNYhsgGKxeIrF8qfTCGnqLu+2V5VPDPW9tC5UTklLvh/lbjZFto0bkg81i9Hk90Rph8vBrQ0e
XMKRBJ7YrueLLcnYibJHwG6a8qG8j1RZNDOFojWGgbtAFsspLqwQgkqRLJMYODFkNtgoSnK2mngN
J+p8LDyqzpIZLqmgoIYR3bHKJkhF5oFUo1Su9RvWMfOgFAbTVbBCX59mkK132Gi6edEo+hRTboxB
UdJyCCb/CS2wI6pPfzKFJNYj2qCmLp6L8u3ZvnPzb8MR+GWOeZjlk1VXWeZo2+GllWKC+i1Wxqy8
g9XTSjEyXxluws+bYe5Z3h8okSTRacAd33+Ph2oBekVVREh5t/C+V1uYIRPUHHmFetk1szQMYNG4
7o8qfLarJqX4FxR616Iw4YSDWvs9UIRLzyypBdhQTHg0EbaJwjygML+6f9gQYlp9QgeCdKka5+C/
7mrij9c5iDaLVdJOvXL2xSA9Gri6hGdPBqImVlUWjJ0qgXTuhht5uXX+DM0lzQLrdAux/CmKmlM3
Bq94o1SxUCqWC4XgthjEXYmJH0nh+5cr7Z03yGT+KUEch8G3sWfD4rv+2XfBwQ3PIWsYMkwBpJ1T
nD9iEEdx0WHmVsj9jzcYV6btI6lXBeYwi0We03Iyi8xCTUQQ4VyV9klZsGh/dW7hZ/2r5CatMLR6
8rpY8NlZgAVb3k/j8k2i5+P/4jJ2MiXoJX0f7qAHCjT4YZtAI4D8VJ3263P72kR/aRPIU45KyDV+
6qRtMvCZDLfjAlgwzVEiP6Dm3LSF611Dc4wwxPyTurOesDWlOtMGjEkU8K8Un0RbsSJnBV4QFU7e
tU326hjVW+ITw7QqIrDDu+RhAUIWrEmdvI4EcBpnXuiiI0vQ+J6jUQjbj0+Ra3y5/UYWiXyIH2oL
G8mWSS+m4iVFxI5Otg5obYHzThMvtKwyMP8nAZzg54fh6WOWdb+c3ZkT643gcShaUx8J4lkEtjd6
bG6PfgLukzpnHPpEK9mOPaj5vr9rW88Ca6REmi/ygN4rFvPw51RbBgDoxdy5VF2SvsPG9Fdlqcu5
WVkrOnQkSkJaSVQermKB9C0ruhJWdQ+W42VQ6PO4UCbcu5cebU37npy5IBNXfLOqjG6ihGuB0Seb
cb9vOZBSY6TuP++uJwKc5BCEqULyQ68Q1ZHPWPZ7JFMCS1jSTZomUixPHRw/f8ugL0WgdiiIa8EP
KFedHiBKvQsEfk3STxpY++FGdPtlfnSfjehurjQhdP8UilRNCXCeuCgJ+sDPuBLgU6sBn8Ls7E+A
wJPQZMs47HMzL/d50z+NzzX0yNH/Y32S/iycvtYBiIJGEia/zB8J7pDysCQsDEcS20YJVRHQonqi
DkCwKRGNWnpU1MhayrpSQv4A4EyuSdGbUq86oHI4jREY39cYxhet/vf46dHuov3qf31OLJbM5iCo
cxM8hb3hVX41H6Fyn3OhL+2DR7bcEHPU7Fooo+IhcZ1s6R14z0VpyPni2nwIt1mL2AGlfaLMWEEt
YxVyy8y0fY2cYNxmN22ekYslkJH2ViYfDPSAJajxmyVM96cvkTYG/SLYodNeBqMdlpULcCBFC6Xj
DLNZJiipJ9FEcb8ExFz6nW5F1fyRwFO9v2HkqS7QdYEpWACtQ3QHTBIucbLfST95bFruVp6lMeQl
piGcU65X3XB6mYbhRtxEV5tVSsV05dG1dYFwLrigwlvDYLXIPVX5w2nrzx0p26mg/p8PhYuV7JY1
Id1hN9nLp/tMbfCvbBV32aKRndoHOF1JzvTEIb0FTdhBUpnO/72BJGZ7JzdYs9mAu748dXZ+xoSo
Ma2K4vDFJP1b9aWdV0+yLmtGxx+s/q9+BkPAN95bXs/U3aD+fzKhHn+Yuim+Bl1czdjT7sb1eCxx
WoUrpcaEqk0o+hAW8SWiuCTJSpoUHLlVyUsuzpZo2yPxH63L2P14A0orGXnWVE4UVyMqSc6O/Q/B
gv/iy5kgHk0NbyAJmMLLyXE3bI9sgQAjXoxQI8SSzAEH+p6ADfDHC5srGWV4pyAfytkt/zKdsT+L
4DSSLy6SmSkFbK1eGdProLHjjVE3RiUE1oGMpUM0M7Vv6waZBnHNrMMVXO99gYT7xt20voKzR63F
JKa7VA7saMDyMRzdDjEJP4FaXIS+G2WO0bF/bzIRt0PKSLFW8027fRDRImx01q0TbwgcK/fwMJ8a
4SAUapM8od4hPyup941ktgN5dYlqmNhUL28vWUpMJFwG0/Vefpf+ZNiRy0BMeefAInTp9H5FGMCc
Mkuh0Hntowg9qfQwbA5u9O2wvxBkXtvBSP5aend4wp1jAlaOBPucefahSrW4FFG3HmW6aKAwN7Pk
P8i5aKmXTfVGFRa66uY+dDcxMMtas13WN84TenJVLTWpXpEF6tr+YJs6vgnCsgRiWFcyPVM2zrsI
Odx/vLV4EUiUOMwQSCJpNbjzvQUX3IrxvzB7JVLXDAXdQztrh78m1ba5cWpva02qTDZN8+u9KXob
PW4RYQU+iCNZDNinRhH/hSsSgvw0yMb284q21Y6/TonEvNso9zxwPkb62roeDN9FuhUGd5GadFP3
EwIustxHVrecOYdCI1vEfk3ZFqK3/kkiPco4bYDhV6g0lP8ntYHadorvFtIH0pjN2w79SRv9VOZ9
VrVvKzTYPqXjwjP44UL9oGpyEMQF1av+ON68kIop9bsqHHfbIrPkin6jk4e162wxUcNH5l2PChGu
UE9jW7EsLz8wt40jdeZpAVwHPxY1D5+AlwL9UdNvly1vHq7lu4YZvrfvwRA9qQzLyK8/rucY4Vlc
Xzu4eWL85xtQL1hEedIW7HiswPe4iWANGXSmO+eXaf7WCSvNhwmhWD4+2kKJGOMTaoJMZsEBaPvr
oSis7CbOwVIjPO/W+utZdxCipLQ91pH498dNICyTEKqyBkXEOJKpYSP+ehdUuVKcL1FdmzTIHJSc
XDlRxr+NdHpuIAqbQbZnlIT+MQ2/bKcQk3tazML3zWWntD6cqDTB8vsTTQnNWsOYz8d2tl2Y4445
POU9OriIPX6wy0hRnvWvkshJSIpvIViB9tOWuyrnfLoG0rXRBEBABL6dZaWAcia+0j1R+KFjrE16
ACxpbrnN7p+l1G2ZdsMB3/AE/KwiPGgE8BAP/DuN8Umg3qHPFRYP8rwspnaHiKqE/XL6OROW8uwD
X8EfteR8zyRfGyx9g1N6IvjiBPANywFI2xJLsglE6LmTIwCmv0ZGlTP3oUFCMg0Qsd273/vxIg0I
IPafrMLBTGCL8AteQYY/00SUpaT5S3+SSMEJxGSipYNU4Rriy2zSg5xV5izPSmq6r/lySc/7Zq/Z
CNLRPyUYhEVfCs+SJFHqlv8L5EWesxasfl+NuGdD9O3L+H78flkw0YbWTVPGgbCRPjtr+hlwGY/T
70+MhmSpFovziyNTWqIJjXWdG8vjLimT81eE8SbuvF/7nhlzczE25jnujcrcQxV3ppMPg1rIsykW
SDPz234vgeC1i8WnqG59swxNJdS/XJmUBhAzd9upfFFLtCvuaVicSt1AWE3sBSKITq8Gaa79vd6j
q5Tmr9Y8dafYgoj2zYRvmFcOo9/5VUr7m2BgVACK4Z7QtAzUmszlTs6B2PmZyUF1KFbPsbzmlF1e
yLLMyw0LV5NkemSNbuJt3F/lxHsgHxPNmrdsQQ+G2dc2plFO7TuvIR1UJTuc2gD9F/WWAj+Pxp+I
SUfYKZZ//Fw1q1ZRKvORbHAkWmevl52MnQGTS/+SCCcROXcP8Whx6szQCWCuosNKJT+u5AA06aCY
Ot9p2xg7mGkPR/Ch2CaSchfYBo5gOfe1sJLWvyqoTrKWiucz5mjX1gBnZhIzLwajw2tYToQejMek
ZN+vtR8du7a8KICRL6r/AgOeMNszpdG3RGA5V1BMSOrUXRHkYck2+DMzUPXGlLC+L+c0RaKHfmw3
ISCThbn9+xps+6cV7pEymTd7OhxJaIuKuG3VOCgTZT4KzJmJQ1Pd7wWH0eb+9GS5ppmJX8ugF7Nr
d5XGIX8g3UUEQux39VqlJbw3Cg/ow4nQp6tuu/ai+AmPkIXpsu+hjavjRTolTX0rWI1KqwCnUNTB
lcgjWeJR1qxiroB8MSfXL2NMG3d7pmev718SrECA30OLdqvUIPKBVnGSjiKbapbzZwRhAuTDxMXA
9UW1E+S/Q2HcAh5cwbORqbimXYZruXesQxtHTWtxnXO1chzoTWMTrNIoVlnuuM+AqdvT3/bcRxxM
9d8b5etULzy/gmX9J1ltVUC7C96aL5pcZYiP60fkCKDddYB9hsbAZ1z32e4sEZckb71dWylR42iT
lGJ6QrLb7RJDr/bn206sUbecO+HOHvzQLkQkPHZHmPdNcRRvtPcECBASdLVeXDMeSUNQGVPTldaH
iL3fel0nqUdd5TGwoWe1odz8R6ACNHuTWhKiuP2/fAzgtroGs7cMefs0VeFJdfFw5opA8dSHx3GF
J2bRCH93qdq7b8axvnp7IWfrVmmaHOQ5OKxDjT7yI/YvcUR9/Q8OlEJllELHe7JAs2GWom1E5o9W
4x9rUFsfW9e7B0+280XBTDFmhV1OxWp59QZAi5G6irqAg5QQWAaSAI7i5TCyVJ47OMuobOrk6EZC
54Sju5b1Qqg8eTpcDEO1nU7JKdBHiPIJOmTj1H2ePb6QzbyeQ7FukR/Jk8dvvZthdZxacIJRG9b1
N0dkAO/tx6k375vcnfYuaTrKsWT3BgrOgOwEBGmRKZ3go62WmZGSsDNuO46Dc725Xxi9rnkRpMiy
v5xk1XFLk9idFVAURfWyGAsPN+eYVKkXDOG2Vq0kVdsLByicyBBLZ6039W/8OluHFQTuYwYMA0pG
OKJPYBpjZnow3QYhCfuMEVsMDC0IMjEQqUvxLat3jRo0jW+pnhQPe6C5TizL0nG3xCoUDxjR6XUB
ZY282N7jW0XYwN1hb9HIDi0erH2sIW4d0vFci3fGuXxWT4dgM+flI2xuxM/c6iaE/qpteXdKMHyQ
RlErdz2PZQ1KK6oYolU2T6LPZZfH96jJJwGf1VVkBt4nV04+vz3v5xkE6zPRYdKsJYuPuGSOvL9b
1alSh2iKxoy1iqwIMNaoN+Dk7WNOywoWM6j+UZMGPBfkNf6v4A4P10yodDczrO6Dj3yoLym+/bf/
8irtul1Eyqg2rFPeeMgfhUNQaNtBYen+bpWOhwlsECpYb0nrKRVYKzmiEhy1eZTHQarG4s/WvZZ6
mEKKZ8lLN2a1idjBM1mIMQavOKxq/g+WQpLpn7jLvQIR66uCsGpzdpnlnXV9yYjCCZlQmBgfC08F
NeTo8DXxmJBqviJNW2y1FCo/XqafBHMZToNDnt4OwpNbco5fWkiLYK0jUnvxSX2IarJh6VNe4J6+
DBaP03G2/pk3F+Zejii6dPyzA85E/mfBHgbaNvpxOIj6BmeroZSOvz1w/XGPaMvR3cEN1EvCHh6k
W4yrvCiWAQYcQ23FMSiZRNXQNOT+TKhYjj5+Z04K/A4Nd01grsCmS6mVipfOIGFuffafyIY/zZ5+
Q9OFE6Wvpwyqtl6/q2AI/F+L2cWlMhWtPa+jxHg2r/9s9WvMpbpYQqr90M0SJCTx+L5311fFf0J3
Yz6tB5MPmtBz4QvpeWcFXdp4IJSI3ElrWjbD88t4dwWxdT2U6UzdL5LTnRdbwUncSr54+te+KE9n
lOCNVcL1tE44IMaHnIUvlaDkRBRx/CrKzDRY0SudeBwnjK05vcrPMM8NnkD+iiy3mZg+Kui8ivWW
ajPCx/Q48embtSnDD8b8EX9tkEpTzrSZsohRJNIj2wQahjdcFzGReRCVocRLTBTGCb4PQnt0J368
TCtUMHjv/Uimj67KPMaZkGLDFPAwKw+k32uGWsPMYY+OJJR58P7TIyLN6/HJC1wh1BAaLfWe9ij+
CxunmHxyvAgiq81ruSUkUF4EjL2GznjGcnLP9o1MwAR8zqhuR1S4UCMLYXSUi1BaY4P3LvcbN+qm
U7wsW1sPAaQsSnG5GSnoX9UdiTllx6YSymdVhF9vpbDPGEdzs319Mepx7m5VN59mSBZSPLF7N8bg
tX+jMePDBPTQr7n4m9hwmBsonSGDKDykL0FEGsUXKU/VTKmd9Xhg0EFNihUpAdmeg/VcbbRgusuq
EJ4+jgFGBdFBUMGaM6ae/MMSJU0/cvYxUi1a3whOSPX0kJhXO4B25UKOUNqYXo2S/AF8OEhSf/Jp
FTi3/DHCEGEzw0Js/Rji0TQkn3IRzLVLkn9Aq+NGjlC9mCgCVCd//n8VO0CxO7Kb3KlXoF2I8Da4
cH3vn9PN6bQEUsL+lEsFcAV3Ppa8cKUEiQQk6l6WhOio0ZVUVPdOKPqdsAOLxdDy4+XXXJ+zYX39
8i5TvrKX4CFNqY03kbEE0qg4JG8UWJ6avLA1BIq98wdpRHrRiDRLu6QFhvldnKoGAptO+a6SzxJB
pn7FeNnVBBdDD8GPvA17M8iEnplZXzbhagYGTePi7LC7xSTjusuwb2gqgpDqsBxE1s0jXm0+ju5X
ZSOuLX/Hd6UYQJRUVKrdE90rUJ3KRkbe+AfW19cljWPGe4CnuD43EC7s6htyVEZKloZYwQzW8iCO
w7PwWYZkLldqPRralhSU4mTt3XGfb6w67glgL8nCMsgxrdR55w3oKNI4+6DfkNOCbjYF3LXIA+BZ
tnLRyd494p6kTd6k9Hrhfa4pDLnFaNXXR4w1QCp9RvHotv8ioq/sD+1GbdaISKYbzbA0DcvHksrI
AvvGNXShKzmXfIMQmO81g1cD+KkuAOnvbaxcmL7ohF9WZWDi4qtFZjzi9+s0p9gSF4esSHgK94Ym
s8rcNh8k4JKZEOoN7E2r6T72cTC75DeVB5bOdjGneGJkEEMbjgR2bLff0yQ8W23lpolonVumbbf8
U5bQ/x0TQRJ2Twxfl9R/CVh5ue3u9PexDnEvAo0Q+Q3vy7vFcip7ltQoWFLs2J+9rLkN71NR6PeU
7Empe6dgH4rD2qFtOYHiCof6d7lmpr61oId86cAKHzDxr+OYaKUksUIgNCcUdtlILHuzcboYbxuz
3TyyBd4go/7cR5qFyXoCfdUgdBbo4uivBmDPNiphSKODqb0TaklRgRS1m3irdtn9xYB7coY3gdfT
NYWgbbRqHmOnXClPEmBM2vjl4vOCf4Bz0WriMyLsESN12HBuX6CGjWikvLc1mzisYiFCo5CP6vg4
LEdavPc7sfiEQ9YABXKrzL7tFtAN2zyBO531ly++YVPI+FHFVBHmqsYSUFGZmkiTDQby6gXowFQB
XsV3hP9m7QpmsBn1ybTiqVJjK+ea112wVw+zgLZYQJVOhLf5uMNRS6wErzBzSBk08NruvK95sc/g
o0I1+piXVo4A/JRG8kf4zMZSB3I+mOAHhMkjpEfEuwv1KEkgkgwAT3komtEtQ43PAd0TCBbi5ahI
L46Od0qna9Zg8/uf4U2eljVl9UxmvkBXUBsP0vYJ+rJa4iTfHCZQlM9+7EXnAinLlXJPWsbASorm
4Ob2T/Y+qay5DaBOV7XOorpVNf1xOUNYe+F9GDq9gVSGq5hq4PutyT0VhJWsZ3r6H0PcrpVg/J1l
DW42xR8Tc6y6Ega9vsdEkM+rDsEKOAKDcbVn57flPR+y0Te78bcIzi2sGRUgEQvBjeZt0BxdlLY6
4Zpbx57NN+i4sQ0qFmXZDEHAxI8mbA89xG73RUl6VXkEvZndAMCwrae0hz2Nm+mvpZhDKcfwOvzz
hAbdTs/GwNje//2CIX1m3T3j+6wHVihkSIC2v8vQDsWKH8g4x5IJrM/+v6AcBH6OQlm8lwqRL3d1
yZRMkLpVbNunTm6V+JF58cEBw400vF7NBj8dytIyj+se+wzRg10Z1MTCXe25Kv7ZOmDcY0zoFke/
DXmK04EBSNv1K09VfHdaQBIO/sykNrB93WuviY/aw4W0idKcCCATTJGMpuRyG/7raoXjTnfxINX7
lxzyrtotXSgHbNAggyOhrrs+iMT+4mwxTeQhIJgzp7gXI8ajm5v8KjqUm3TkbLBG/AMSTzdaYmzI
JdImZqFmWtiZqiQjf4VVIHupHC3derSd7UNXO/CggnTvKF4/4k8/x0SjfnFGcMcy9bnxNL7R1fmN
Mv5aWfR+PrronFPUQBdwNNffFdCMQiRv8Gfpna3SUZclOvkPMRsRxNfn1wzwGTPey9h4dl/6TPjK
geZaUJT3m8ivtorf9BMvVylDA4A145+gXWUzEKNRjtT/yAHsdzBMj3pzAr/F9VSmF+TtGbV+/Jx2
u8kTGhICocxZzjTfbi3vO8/WHb3gg9Pnn9IOjJUWuSiwfxKhxMMCqjyIKQyj7KsRehL5C/zl9vK4
UwWZmuK8oy6fd4fWNTsnKjnOwKb0WTI316/Srr3yo3A10pEEIvOETE9sOsjP2FeTBCpfGni7+/JD
wtIqoVzz5wDJzoacDCFQ7gCYxb05PsxizWW8P3eYkRZ4DkPk9SPYy92yJMFylbY7w0L0G+Dq8P6E
4o2tA5LZP5O1CzgqIgLg0A3wo5WOkMooC/G0ui8GPJ5AOg8IIr3FwxXLD3qS7hCqkVZtQNZo88RD
XAX29bm6thuBQnVrXJDJrx5aJwKa7+OpFSx0N4yyaGofSdmonzUaq5LqTq3wSlG96BCA00ELLnfx
4GaUvMFktIHTMk1fpTppgiN8k2nWsecLQKi9pEz0cp4PlPUBrjCbPbXToHyQYd4E5Th6cUxPPsPZ
0fI5DbXsl7cl1aXLJX+ryc1CgWVTmwsWCdUTqLnVTAvF/ll4YNUvAqTATpPidiHaUjHyE4Fl4z3r
qK1vW+5XRb26rrBop3ewZNS60b2C8NbNMHAk9+B3Ce03csdPq6o6/rc61+Z8GUJmRMkqj0S0srsi
I5laAF0PxNTZ6mjckNOSobaubGUMbSJ2mr/xAJydM+RmRPr+4XVs21UPwexcBMUDJiiUG5hecaPE
VqcRqdhjVY3m4UiLdLquqf0dh4eM1/+76liG97Hy2Y4sC1zU5nA//S0oFoMlVjg8WuQG/ZiKl4Bx
p73D9AtPMLzihgsOugnvBkzPZLk6EhLH3ogYxj5tO5PJXj4XB43y+5ndBwYVHPuOhpbxpRl9dZO7
ASWPokvIO5qVyOuM3XIIzpq/L+nqpD77X7pr8kO4dquhKi9M7L1ukcywGjRqX41VAI59Z1uLgIGr
1Er8MvTC3g7FoVoIa9uOtB40Dkjy9qWxZwUpZSQLxSTesBqO+qtLTQJW5ZWzUYsKOnSkg66BoCFU
ghbefhSLpQKcIE4LHSiZxB7jepHGJibo8Sxqh5mx1a8CIGqgxDqgA8JmuynYSQxbtdt4QueLzREk
RnTSOa6JStoo8LaPlIEBOYGhq6UJYtlB8a2kz4FXDcjsp5cGo6MBKcW4+OUgp3ZpUwZ5Dr54teVF
aQOWC8k3ralIHdBrLFz2KQ5PEMNUExAOu1WtzJYrJFGFR1QAFtt7pVYTcBJH43DAVJYgAnkKtLXR
QV2TlLDT8EBM1hza6hvv9E08ElM/WJOOD0ioR6NrYlrEEprWRqwRvLPmOW9TlcW4Wp+VaH59erxs
X1gA5USysOgIH836fo72Q1FCpFYN7n28hU3V9w82P77paaTwNiMdIp4AlSX0w6Qti5YX0qRJZ+rm
e1qv9O/KmembzC+gnZiGltgIcjERhCAH+Iw9dJEbvJuMT2EsNMqayHEKqJAUieN4iUc5RlyzIOoJ
n2gDoVcCJG0fFwqKUUgsEEyuZOLZEazmk8BWDP6u33Qe93Xo9ASs56J/RhJykDG41iyIs7mCUHDW
j9bbdR5zgIrHtgbVQ/hXMFMaPW2BPGe82GF/mT1XUQ0nu2cc7ywzA0dLOWVYewU9l3gqfEkdxvSN
Qi98rgoimiJZkBNO+pN44L0kjTwb1E4GM42Xr4h67qFFkvnbTNAEbPUwlK4fm4wlDpnjTywMwk1+
yxXwLYq2QiG1LcKRByUpUSkyOwqGBv6hjlbYGzMea3TISDdv0WjIlZalHaLLRZFFPytAalxQdNpo
J12yGw4K7XWSqqD+5RoSi3yqfqYC5XFrDQDsyuwFxGOnxZMQmvI4gxyV+J95nY8/o/hIbklEe9+k
tRAjrA3oJkhvNoLdZmSGZK3is4qGS025optGxiX4iGZMCMMd57k0iWLb0veHT0FGezLHiEo5T1cC
be1nTocLskxFT+rlecgGZXG50BpkGdiFzN/SGStiLswtJRmLK626ftR1usIHeA1RC+cOctgp+ZnU
cuPTEPh6/PuVLTYATj1C5MkIwNQgdaSHD6UPSsAJhEuu5Jud46mfWw0YSGVUKb1wv7zSRZyVmfZp
Xp0x+KPznNoT/3ls68bvxnkFaU1GyvzBt7vcV0F5dVx2jLXer7N8y+ypfeF9kDMby+3Y5CquFEvD
iu388anCVMWf2zPUjo0yU0EU7IgUzDJTtQgQDhAQkqnSjeYQhMT+noV+HUEa/Pwj6Bp+Dvzc/DTk
bFmELZosZzxxVYAez4gllbo3QvaAMmOFGpv4k6+pG2BhzO3NPs3+s3ahGAlzvOQBMNpOX7vgI71B
/zHWm+vUENEO+dODAO5D073lW5RttS1YurtyzN4wCMz8Jq+FoAwCWxIfhUjKwphdgQvV9yPL0fOt
he7BIu4s7kxYq41RpIxD4B2iJwIEVBZdEGvwm90dY5DI5aexSnJYuFJlzdZeLAiHSQoQyqhz2LZw
XE2elPVrhO+VFU72YP8ETNvJ2y2s8HDXldfYtSFsAeFwYVfRIFqpgl87AV3z+o5I9v/I2j6mmZFd
nIzG9CQuGd6bimlLYoV6lLwCSE76rY81la4bMA6ySRmKlqF/6RZTRVilRURggQFxJXmcpPJv/USp
ptQKHCgvuaECJwAGCIhdBqpNfVgM5C0EuOl9vyRg9p0Zkrdicozd7zQJwDM9FqIbcc5zSH1eJ5UB
8e89KTT8iwh7He4zxO3nHECJxTfNDfztVY9eJY0TFPPHsAscOLaf1c1aW2s8aCbCL2PjmInOimDu
QyziLTby5dE4HR6nMMfOQK+sI8cqe1q8OuF2G+qvujP9la/TGfbWimlNsHXCA5RnaowxhlwU0fHD
KYD8PzqXul6ab+1r02NPvwxGSQgWke3Wyo/lL6fsvdrxQnvfjdjKOEKihgCkXmwiyooh8ZlhEIVK
ZAsg3IsxNo+XgqDsmHhxVKOc5AFXNJYKUeq6w4L9DRJ5PkDTFD8PvubZa1Jot123eoeD6K5+FySX
ceWC9mn95ax0VdSkI3KqlrwOJJaIKGNZu3hNa+pv3l2esJ8CpHYw58R5hcNBFo7AMgYGLATf0Bha
9IYFBB4KFxpEmmuq8/vqlfqvrxvapYokz+b1rZtm4xVq5jRnTi0fwvLiqG4coQ5DrO7PphyNvCOd
5RJ//bipwgRQL2jcYDTcDVjnQGmZHP9WEiFvFaLi4izKF2c5aCfJOO05uFBwijJYxcj0LBPDQx+7
t3pegCCsszeuH1YqVF28harBxyTvjBiVuGYvkOeqe3dp5/v2l9JS7qASSOBcKSJFqfyyGtAw5O1h
8prjYtx/d868lek6Zx2ySQL/7RuV13lup79hnEr1LfJkpSBSy01YkwLNrkcbxJSxyxSpc6LzFPbF
wLCFdLJy5K33QPlxiAc7rWU5HSeTHPyqqc/H50RwlIjRrVgZle7K0cMMrcqs2LaN7yCdYda7BoVe
dR4/dA9SnDNVxp1RX31EF703dYkjUIf567NAhG1lTtGsYbXsLPT4f61vXevEF0M5eycXJEseZ8x3
1ug+a1T/N2st+f/tWyUSOCJh5mKMfeDzNxypvVeoq/iAKKwQ7/yhDM0uIx6U8NSq4wXDoBJOzPyG
mRwcnBBauP2nF+AHHMKTTae+fKsGQilvzNTpA2XKv6SzM3Xc7Bf72XyougjdDTGlLSBvUFd3IdJb
qye0KYXw9QuLM6pmqQGLsJEnj01K3e561iupWcFIgB8v65A5+XE6DkjPax2r4GmPcd8uhPSPSPBo
PnmOYzDgA8ZMQXtFMUk0GG7a15gQFWR0fRRd9jpNoP73AeW1TGb/BKPDuD8LXbjC5i+4qczDbLPs
4cdBA50LrvDdrZTOV7lgrXeLbTGk2PSh4elbap+Oj1zUzZsLV5Lhix2JIO5uJuQBNy822h9quXPK
6+W6FsRL00Chyk3z6qW34di0FYDE3ptQYMi0+ofKFI7qUhDScwkd2xrnon5IocefkLKAoFGhbIwY
X56ECmbjIz6E/OblIUXOeSHZHlAC3kMEhy2/QukoH3X9PTZSBb0/3Q5VyZ8Ecq6ZrEqMwaX1EXuH
KAStVsFoionRhmJJCGmoGUbJLA7O3BBH5cuEbsphecD/ttgsjqkzgv/9RxOwr3isuD+sFM1x9qQI
R4MvS0IjpuK8MZvqdxz3T37BPWzo8SSNJ+v0ctAkso/qwTExHKMsYNnfTT1Ea25PNMoqMj5WgdkW
snRY+v+xT+hNRz6dKITu6hujl9251EkKHzW+SESHRW4k3vpwAlPu6MRhQBnxTwe2pfWTRhQ8WQjW
dRfFYkgmuVG31/zwsTLjayyROTc95WlKiGEvHTf2V1MP5/39wilkwHox4GX2OzXIfGYLUZVYRRSZ
+hBGPnHPVwqDHX05hLiOFfeNkqcbYwHBU/NRPvA1fW6vlyJmMFaxupGFWQqLMrV002bViYN8KQf8
Lkl/+3jqmDEPtAsIP5ZfGPrNnbG9bez/4gna8tEz+CQRx3Z2c5tkpiXHnF5CPVPRUzVh7WcyoFor
ZX8CAIZry6FpgErrkXxrg3krl0gnh5wvS8MGrqJQICeS25F0WfUbka963DI6lZnWJojxpCRwfqx+
l3PCzOaCl39bryQrzDYVovI9x5A8XqthiHua3CI/C73YMMb6+Rc/ADSIyMx8MVtZc5A24FOyPrvj
1748SdK24Qo+H4pjF59gYd7iVmCezR2up4cxQnG7iG+ozQLQkdYKRu3/h7Bvxk9p8QGdnrltk4HE
JYj7tX60BpFqwD17SXJrm0FzQQEcwcSqn/LcAKguXEnMiaPRWTEO1jxjWo54GhPFPftGgc7ARVSN
axuZry0XF4LEezlH8hHOsaBLsCQVSXoSb6m8pKu0tqhsIUVL+apyVoRfVrQzfbs3FACHZkI52mzp
XtmnZVAEmvxyD1wckkHwvmIR7qbrdyi/yl2Ux+8Hgljr2/xEgWKqLfOyEpIiblDBnhoHvXCQb4FV
J8VkRfarorKdyNRYD56Ic7GrnKu0FXtfBqeRo6/4OWPzzDaG1GQ1hx0WQBjXp7r2QVLdjsML51Ke
jM6nSa1W/ydhYhKOIcG9m+HbgaIp2h8dby2Dg8jKWilh60Y4FjID5R463G/M/ZYXCTNZPv6uIAcs
U0020HRp81zzL9Ui0NDcxe+5Wswi8L6gNrE0XuUktAmSwNyeXrPpCg8hIN5jAZbZnJv3j8cusjmE
MJfD4tIO+CXFhodPCRW8AwQgWOak/9QLOKdwRefOP5OE302ATeCFwbGrvIxEVFjYVnmzMt1FAG6Z
tr6eAhV43GP7KCZwifEKkX9iYMrr5bBwKVg/ioj36jjvWnmEZuWzmjFBCdwb32h9drifUj3xCjbl
y/6+nlwtjcWXploC0jb8mQPhvsRSvMhvdIP9WP3EWzkrpPT4if2VFLBsxwWDj5R7+GKNmWkQzGE+
1TGmwEfRu7W9qyPn6xWmazUPxY+HmcfnoT38XlaHUSJAvFE4bn8e28icq1OKBbFD8uEcANnjcOOV
CX/BrPZkaoddPHu7m/IkBFR0fD1jFdHnf86ja2meUmNou1XchM4hIpWEtmUWf1hcmVF6w5aHoMfg
9CGXCH3AUbPM4N2F+zL2JvxclbYBoUGiA7qxfZCPPoVN0ZSX3k13UkJO9/P7ZO/3KexhkCbVqGIk
B2zduRLFJ0UwNu72SC18ra7m5Z01Wid4NXTP6LmV+eT/JG4OGzsU1Riqih7nQgyb8IqyNaHWQ93y
ujGt29xO1R0fS0qgV0vdlWPzkwNpE4d9lmi7fY4j3XyXoPPll5nSLyMdv5jJhcdj2napCfgBq7xs
EokURC4kDU96Wh/U8SFRyVcbaOGBa9BLbghNmqP6k8D8M9z8WpeFNFq7XX6WJALY0VxrRSz3U59a
2pJyBgFEVhYKgP7l9kLZZNy6N5NZn7ljrAs138KPVemMXmmXq9yDtuBDf+60V/pZedvhsN8E/oh4
Ws2kR7bC3LCi5DXNc3pgXb679l3zd8vMhVJn6bx4ee9IpoMPR5lXteAJXjOisMvkaWDxuFdWnk1w
vh6tvPrGUJyp05PISUv3lYlFF76teDZwHRNhrVuBu4s2vjzSXWe8Adn/z07AIIKLULLTROjz6ROd
6DwYPKTZf4HedEVESHhFBEuiA+tl+84EEQG20vch+VG++JoqPWA0GG0dQXaDewidy5oCej5g78U/
64a8Aqto86UQ13FIAdCLX1t1W6h8mi6NQyhJrbRUWejlSRlqh5HjlSs+jz9anfsGCyuEoAjQEs+N
lgigQsbo+WhpeXF+CYyDyyIRpw+tVon2C9w0e0U/eU0mJ9cu+yDNfrtT8q2Fyo30+YWeskYSsp8j
+8/1Df8UJpPfll9zpGj8D8xwBb72kMrDf/M+rktu0Sm/G9Wl6fITWia63trFGFDcnyC9pQHiVHsV
MvTvamirsdCB3/1DEyJFbNe/MVCxTOhWSkZa7U8/OKHVcF8pTE6K6r+nj2nCCkJ26a/JsRueLH+7
7vc//SzOTcLQHBoRHZ1c4yAXuCXdYiG7qsednsViLvUa0Vk+iRP6u/Rtjf2oOS9gDexFBw8k4BDX
OmJqj7NZ6Nyo1lpwOkQ5PCkAj2SbsgorK1Z4lvJBdF17w49sTcDZa5GCqgXUc7JtWLShDwTr+V+j
BahbzKysW7z2LyRNCkozZJ1M0Yea3iNHJ8elKaNfoalwAsfU4XI6CR3qmmup/QaQLl/deRYav0Uh
OzxFoM41bMCk+921hSayuA1agl76s3G2V+DECujX0yNAVKCoJwnR2mN7IqmB+PEN07rb0UBSbFFg
rWJRqkVVrKQ4UA7g0IoStF1M3v/5qommTKgb82pQ+cBXEuzp6RJR2/tLsDiiyKOnWUUxwYa8lKL7
G3ixF2ilQl0NDg+L68j3yUDGaBPNQrweERheEUqRp8s8krBG7oozYhnpHcNbLtnbWmbdRMRWa4DJ
JOVcmpcRrhnztWB6WXpWtHyfBdnr0BMZw8oior7vILtxmpG6D2D4Kp6IxUtpq8HpjOv1JYCabgJU
QgLgWCuEP3JwgtrebFHcWdlOmwkmp7SgCk3J8JjTPLqzdRBj4cxFIUrvJfuNiU04f0xJRrYgFLoF
6p0z5G0UF8zdExj3mm3qBALmYiv60eNcIIF3ey9wdzH8X0FVWgd/PYfIHenaxqP1eD13BMAx/Isn
/kpWLaxLscPi09yj4O+V4XLpBSHi8xsO5j6vM0cV9acy97uuxpMSf/x0AuW8gRCn4hRy9aa2Ne4R
YF0ALZWr4ewjNafgCyRSHf/zPV8h8T49EFK/MUmtMB9rU2vY+jDzKoi0YqQOkcx3RrovJb21helz
c4XHIhQ6UqtAAtHjLdEmNVSynrksMhnsfjdg/Dyc5sj2x7UEdRqtowtyTl8nQm7eqNn3Ye8UOAY6
lvMGggKgEKoGhTobDNJOroDrBOysmlCzr+RszbbKU4aG5opzADmfNUpIWV9inVrYDRH/bO13/rr1
CFOZdGbXfKGGW4+2pTtsAam1/Ai5qg2BhyrtP9/HxpGNenxbp7q2/TOnUamo6T6KtVqh3vOgY0rj
lCpiP/66akgkBYH9xptX/x1C2l8NJWm/wQzeU3ARZoLsVQS6udq3aUgLpjPFEKQHSBfdA+aIjhKA
t0biwOceNZlJcWISnn+Lt+Y/OiNHKdk2shnVFY5wW/b6QDEu2oQBATpuILslk3rc3SL7GaWfbqYA
V8DcNGEZgqeJp+JrkF84TeKjluVuB6goqPWSyjDTGylvmARMHGnWSf05mZGpFH0IU1kv6z9EyKfH
4s4tUqUDA9LU7Hw6ux++KGcuQMqkifofTXKxxZrdkiV0Frua8I7YBUPNq265sOSKe0seaxxMdJEE
VViQvTLJDVtnEj2hbJ5C+E0Zi9Xwo9jQz+eiwx6kciNc0eGXq6WG3JsB+bpAS545YfAheBIK7okB
FDTO4zV9Oqhsh+WldDgs1EQzMd6LZKKCxO01qjmh1NXqh56J7Oh64uYG5ZtO4qcJ1wBDtZoTBynQ
/lNXYPpsA0FjUmL5uVq7BlghFPfeUf9GPwg0pw1KDY47G6JX6sTu3qKInAoK7Uwy0RuOYGxvlu35
+JKav0KHf8A/Q85xVt6FRoGIcB/dNbCrOoMhDKPRyQXvtj0b8K7anskcviI0CoXrFcFiyeDBUf/M
WKepwwUM36ymX7URDLSSXhU3g3XuoatZCh9ABRiafO24EBtjS9FeJ5QNqF45TueDARMJBYt6+ExI
7TH+uAV5+cu/H6Upjv4qIdi6PEl/WBMCk9pUqr0XYcJ5vNzG65Cw7g15U/LSE+kCnnTkAmt1x1Ew
5TQXOh6dU0v029LDDMeygSmX+Hc6auPGViUrejsKnx7StZDO7cI9jdd+p9Hrp8wPxjR9nRjBs7Rr
FoYgWkgJ7EpgSe0xdcUTIMab0aWGJeMhzx3kKpVZcGnKUU/kQx3R3joQ1mgikbopoQszGDJKdxI6
OI6lJa4k6qM5tndaJHJOmZCIO4i5bVzMub1QVYw9ZbhCsgMAW+456YLrBz2IHe90dNP7JCj4M9v9
Nf/jNgpvOnL49D3nWIJOuiCJAA++aJY6GD1GRcif7aP25iY6plPiRmMreu5JGANGKSwsigidiJsQ
PuWK/yvV/5LFBucN/WHVEDEOgTvsDRcJK6Eme1ggFBTsVkesbcJvGDfDWr6C/E49r6+f48ivOB6M
wHOjJ1RF3z7K9wrvr4jHaMOwtUY1DokaqvCHrsnNc/c44jksqNjP3lFWDoayXjoADdPoNO6pJ2B8
CPw62gyqn7n9KXtlWfLnbOpPZhrDaXe+aNt2EDe7aVM0SJXZi/HRdpyBrG45rYpidk2MEmmAphwX
5044YgVMTCKeqaPvcJbB08XcMcNIfeDfkRsr2BkDYrMeEL4oNf+lJFtZw12jhigxtAE4l/nkDRL0
cf90IzxIE9GFwITh9/AXxzmt/rFBV56tc8g9aQ8bQ53W8oZ1/Bjq0vItGtOD7dsy7ZtPDkMC+0NA
nAnw2nT3A8BcaABIL66eru5GmPGB/tMQs8Izxkhfz+hr+HgmA0D5etEmV6/apoAmFflbDgVoLGol
kTftNvkRqyebn2scPd3T090nCOfEnZil7S5kmxKSphs5E6lsxq2nAEwNbwdPyKGaYNplhbS/TUQg
1N9h0Wfr609AgZHjD5HKNLXilWZiSZIzk69b0BM4h+oU9GwaZddCKN9fFRda3Gd5nA77kT4PipfS
/IYDdGui+P4mKJC0ttjKqlxDP0dTYEGFuUjow5MTrDezSqb1AEPP5mVuroBpxuv+CMwp6IPevEEr
foEn/oePR68ZoHLlpXADWDd6pnLq/JoV5ZNJek14HTypjRdYOPMwLztlhKPxaLS7gUW+JO3XjfVo
jzRteatqaET2zFj5+D7cn5zb4NMy3Hs2CZQTpG6BQWrHqKP4h4SHMusgLYSBptljylzwp4MLEJ4X
KueiezxGofWofn5xqZdiIgHvYFHxJhAruwZKmAd/9GO0864h5nsUKRMllGeEJz3rYAZqpAvy40FG
HiVeYVYexy/52tWrsSNQ+JBjgkg4t2lND6Hz24hm+nCbjlfFMF9AYJ8z7sCNtGfkbVszXVIM5397
EnZxtjRtE1Mw3nL+mUuIAv8QCZj2Xa1iA58sGTuUCKJosL3/j5n7GEobHlmIQpzvrrlIag3Vh+jq
pDKOAFrICRFJ2WvJIY3487qlWcWwlpC196SByeNKVKyosuFr+Gt+tACU48ftNPYdHNmlpwdjuksa
eGFw00rcRkwQXDEHTBUBmaPI5qCtQFujpTIYAcEay6AslUHAXu8vL6mCEmLfJmJo2orFJXHYvifE
fkgE86SqZujDa6VCm6oaAlKdN4W+qPGUZZIIYjVBjO5wKn1V99ZT2+BFprm37rvOxJYHfmlwusWN
S44OxCHIO/X7oolXTpj64OB8pHt39PPYurXUqjOlDFnc+fKVfkZ53p+H3L0gIQTuINTsJn5qI6Bd
hFfT4MB3kainMZIGFpgk/84HPs9hTD3gupatZsIJEFTXQcF4TnLCBHyvZH6SZ/Uysy5RmdQjz9+b
uQyvs9UnP3h0E4V2JzfaGNWHf30/BS4bSs8Qe2HAOMRza0BY6vvMRZEmi5Tlcn6Gf+9UZLG4HRUo
kZIA/9zGAOJ62PXN9IFjSuyGPQHU4SZRkSA4IknqM/OHt7H1CV2EaKa7KZAh3ioGkIYuWWMJSGRb
yOrDyBXST8kjGC/pq2CqxyYnpure4gR7V9Ha1J7iNHOS4u4dcdnIGeMNgreNuXf6j4aFfuNdKXmU
2YVxZuisq+iBDp74bDSgk6QsL+riEv14h1uInloh0EfNrEn4AHADq1Sz6Eis7Mf4FJhl6zffweoL
xXr+damcmDjhi6UsrdQcpI+Rs9jxQJGad03s8HV8dTwRI6fsF7vTzVG8WMgCmO+m7pDzvwXRFIX7
Us/t7cd8xdYPDH3GM3QEbj69yVlNA9Rw0VKbYqa85lPBZe25rsf00i8I8agh5UYoUV3zqJTK7L6s
mljuQJqpJdVDu7Xx0P+Mb1qDIN1ioKT3PIOCOGKgWwcp5KrqRZcc8Qlk9aPZFdyB+mOmm9vre2vH
tRKxZf+P+8a7kJjOuyQLaOpqgRS5FDYuTVqwAapbeK5XG+4osP5oeF8Ap0+ZAL1bkBiX5HGVdskK
+jv64+PzJIW0S6CBdFYZednRqzGO2+mTRQh6MQ+mR4c1zWiVhRx1E0K9tpb4zs9u7c3GIFIbAlkx
2iS6QqDvwra/sJykMPEvWmgwgXERRqfjana7+GAVkBrN2tjTdCYB9ObT+Xd7MBWnU63vpQ34QlLn
ZJV03ajYavy6H0/K64Z+iOOZ0qqdzwxb1rcP2TCH2yiGgQhYluI5HbeyTHZXAzwywpTelalDho/W
itTSKdl7oqxxMvWyh5CVu2ZIwYgeykpyCcUIrvnpx5qczhn3Hx0lb56OOfgcuELa0Z4ygMQSgB0N
2whtgO3iWbL8OT3th0XHZXJGD054W/j5fYbatf7lJMzwmmZMxTwbTmb9+n1n9zSSOzFVfCEeKtU3
Hh54SCi3eNIszO4R1REM7LFV2uf8Nh4qmWwubixlaSJ2g/14ydATAanbKpXbS000uOnRwKu/Do3b
n4a3k1wtQ0T9PFJfCjUNw4GNKO2yfXJxKnKvekjlHklj0psBEJz730UbPYVC9d4DBfawms2wLqXQ
k6X0r2UkGR51vRgWCJi7Y7KS08CYWt4cR5lOU4XGuVc8uc3es1bDwLdgPiUBYbffNjxAjKSJ1n87
NSPxNcF8dK87JbBcJhlZ23Bd5wM31v9upIKoFzR8kJL2VP5imqaSF6VIotYl6n4DuaaWJM+Mk7Xq
8vOC6rWkSOJcsnZ47bGRpP3OeU4hGinfxc7K+K9wNzcGAyWdHtXwW/9gvOAwf6IPv0xZckQq7aQS
n323YDx4uGsX3ODEKQZBh6nHnyUGCR4BqqK+cNgP9vvZr4R4Gdk+FaIcJtJm10xsa6gKgHjZM1P8
4R4HSwkxBmSEfC18hNSKTsZx3XEJHPgynoWcSCtIWFKsrlIwft9HuoWpcVPDxxkHhpRTPqkqyvoU
WEeXQcG5Bu9dyyiPox7CyyGoGahAoY374ZzqjMFJG6qNSOPdg+0Qo7pCVFfLeW1Ub59vbZOHb/MT
1TRoWS5XvDZAM8oFk85XoB/bpUiL1XtSCfvvMSinqmkNYsZWct7cZm+amGIsRHq+iev08qSiL9uL
1GEXRzJhl6AKXpx5xWKz+bUnhbS2y3k/fwyllj5xtBjpfyS5z1flcqQbTnZdaH2ysaQsLW0tbYga
725O/O75CztdovYKMo1HIdGdq+aQdl9isqtths5t9AUgrSV7oX+m/15i4IcanBa+gZHh7QrJUymb
hDY6wDohZJSvveH5kBwrgLwWB2p5K3yKq9dO9ANVOSFBuOW32JCX5C+5KOG3qqRDWUnz8YP9qnmJ
C1tNWsbCLXIkC1pO0X0IfT8zIuYQ1Y8pY+QYNSFoI8Rggdgx1WQ9SQiulF2FgPqhifygzKxcfbjI
CWbc8u1oJ4ESKBJ5MROguDdgOYgbuRU1OcEdeQ1XaaHNdoV9573+DRn7o0ntN0aznoDaVrpG1DIU
CRKHW8MQrcbp+IsKd0P8ayNDtJ9g1yvwmAvzozeKeODPkFA0QH5RmRPTVFRlxcN6CDhpwAuBoIUU
K1E4DoKovlIlRvn34NfIJwQTnU+EjO4pBFeHkaK8ya6kQOJozLDKMrll5yC2CT+hSH1sHjcj2dzu
92/luaJ3Z1aCJk9ZG2JU0M1iQRNjONqfvcjz614MC7XKNUYmybEc0txAPyRBRDxrRcyouG1fpBv4
yGwG5worCIf77mingCIQJbzh65HehggZe3VFbO1r+qp5puXEu1h1IPqoolm04qK2Wgv0q80HLqCV
9Lj1v1J1fGUMylv6uWdwS7HyZdYRAHIqZwXdMao/Ieel840pq28WbCyagztu39W6BxDULaUYAdUD
lt8cP6USx3Yejl6aLd9d9YVfh5onTEG+mB5oF8rNdgBZcPFwHKc2XGjWT7QmddLeCz6QaPdEjsj7
ZE4pQxMeMuUs+9ggZH8uH55fFJKd+5LEKq9idezsqIJw5FEecMzD4XVtK+o9/nVq/OzBFZ02ns2E
NQBcAg3cjy7GJPLz2Eu9HmCWVV5vC+e23G5WekNk2b4pRo1pjw9330UHYZ5x36K24T7HvHYptKZ2
1uVtfgJjoFQnIXzRI9GAoIpTPA0em9+//rGTZhj2p771j1TUvMD1S5ky4ZhDDT8F3NJ+TOS4tUqv
rE2RCkQUyC9+CNQToyLDMIBJWpAUl0nqWEBWx+lMjb1dlC15CuNZ8ibEjLQbRZ/22Jn6jQmZtD3Y
ib1mOSQ8B00Nb1Rlls6ImFntQYb3RVDh/aDk5ALRSYYgaHGoet2AL4PDyhxcss2Y9bFQ4QnPAUhD
fdR7czHKLJRChQlR8Xpk5T9NHwxjbScKj2wAt3PxA1uMfuTe7tNBv+IDHIYcobaHu8G3C/lYnn/p
sOJU8mRAlzgRK/mK0zDZ4pdIcn8ue9xc2fJY1idY5EeNUr5nEZ3BmdlusVyzZc260Y8XpIOe9Mzu
G4FtC+kTntsBP3fxL7OggLwluaEChTvZ32T8QnFUe3mL/svE139ExVyr41bfIwA2dS+sfUzH3Mak
HXdiw1kRspC81sLTNq12ETKlVrb84X8KiuHTQ0kb12wuf5QEK5ZRQPxPGHXO0mR2BO5Ot3GbDys1
QH1AT+n93XpW4oyBHF/3qTbQ81e8/eNn7mXmm9rVq9PF3wmSNq4FjOCzM2ClUpZs122iTqEJJEj8
lUDgumjtDwO1afS0/pYijB0PXz9bbxy7kVQgVDPbC1Mv9/mjlB/7FRCUyxPSk33pUXL4/mNQ8rfT
KiAc0Nvfh9szViLOXiK+skBvidZ0B0bDlTPLmMWyFVdDxd+xQ4V1OFSk246H8qolAUb6yBdCdQAC
jZKMt26rkQCxGcak7XF1w7ZQNbvVjClRpVPPS73NhgIgkb5hZqjLEF9DjKWrut6vLrPvMPNh0h3i
O2EbGtZ9yWgqp9/YVP3OrHZLoOEFJH4QEndISCaOWfYI0vjYC75wEUsUVnq71izMVwbhMhn6PfBg
6ZgMsl/lBsyobL50OwcsqU7rFJDKf12dcCfwP9AQujrBt9ggPIrfwyfvvdOheOQf86ijgZkzJVQd
Y4muSWZt8V63pdX9eF6w1yfS+70guYZ0kxe61fgFZkmxP/B1CuOHAmigNllxcxVqiH+EMtJN3W+b
rzTm5AQNBciTV7ChVBIaoV0vRBh2x8/KWOwwySZgxavUP+TDNy5h/j3TF3+CxYT1xmSyOByryZ04
fxIgPK5cP+lnxn25Fg1fBZeYrSyOcpt9dSCIAzgsi+2X4X0zvx51JaA85v7T6HYdrlKg54X8DgIx
NWCvUITUtimhEuTTDStuDBb4z7y7GccxXb7j8/ZA1xn8XWUWhrw/ZDalCO1YJ8O9tW2YO7Ax4vnb
4TeHEY4yiUVHflGm4fvT6p5onI8FthbEHk/JkD9OOK2XiN9vOZPvrAR6YhD7IlWHiYMvmRFq8qY9
3YLh+T5lYfjWl7y4K+pVqfZ815HZmCS3xThhP2paYtKRmh8HUDaC2qllU0BUwjek/Q1toZtoi86y
DwfS296lMV6gMFaqSju/lBb1+AXx0nMsLGOlW02Np+Ms5qEDonYIG6C6oSLgQXyVBReLq5KuTKbg
CrzDlkdxIkfprPV0AKffDSEgv48t6gZMJ02mOM9e1vDhhA4fu+BX8ZGeEud0hqlpkKkpywmU/kEk
YFb1/8BogaFj7Gz+ep328O6hfYM42ED/ymGxIq750k+UV6Y01n22aqtkFGBRXJiRtuZu2UPihHuL
RySWKu99OMqDZrUU3CQG1U05Gue3KoOPAWIsHiWe21AuNOpwUec+B5hNpW17cOX94z3TFukh5xBx
ssliPa0TmFP5pNEbxCph33X9STdvWeVfPmjwYYBk6GjeiIraSdlav1aTWdktCe+dAr5myhe7EifU
AokisSA0cWCT7h25bFpK90IptnpzTM3UD3UIATaNMFJOSsZMAQ9IqGbBW2Hdm/5o4A5kaLc+NReB
EWyZyKoEOoon1u20KR2D+imHCTzgkxZ/wNBimKPAz/IJ4Zv16V/YVNZMreZBoG+eUh6rXDYIHAXL
w8iQpE2XPAI0mDzPtWrP6yKPug6sdM51eTDIFLS2ICn/jI8gd6pFYVVNTZQfiC7anA0gIst0OuFF
NwOileCyV04fJobSdJ174bwKgmUeK5W067KmXrWK6usN698C7su+6k0zLKopiIzKeCfoNtvigKkG
Ul2py8l6PCJmjCE8G6lKdVlFGu7ZgS3+b9HsbGSQR+9RNn5jyu/I6lcKYJ1TWqJDUea/y8ihYPuw
lhPJGVTKZfQnN3uHIhF3G9TY+sM7IEaYX7ezqgLb+E7A4x3zP1dUVNM0VfK0VlRcmCzpYTzwZf1H
6GyBVAepjSxo6C0ZGrHO9U+xfySM7aLMIk8qz4MiWCsSqSny5/yMditeLr3Tj+soS++NgmF8xiin
4dCMP1cIXYZRhOIDsM1YPFH19WkVcFMABnwKewhcw+A45DU/JOA0d7PMWtLrIfvTkZedUfBmsesI
WVyMl4lLbEXrO4bByny2MipfM9qHdFIGtS2crErvW85FwtjPDdp5ItvGzlVblAwhx81l/AXOYfc+
KTKt1jT0xGmBNv+aoi0ydeUicHQzwP89hiyHPtW/UNu4T/h7B9Ta7ejpHlRs1Yz3SElspz7RRn11
r54KQ45dzL7cGsMNYZn9KRi7IH01ecSWpl/v/eSEUlQ9tqd6o4Q+SpBUlGbKNc1yGkKYIjAMPfqe
JSbkFn/N84EH/f+IxfHEJR/mlYrYIY7gb/4fAZb36qj7iLmMYb0Lsr8QiENzmqqLMSsgjme7DMG0
zrLkJM5fw87txzdFGkoMd2bNofDaFow2cNGtoqQpb4QwcWVUflSfxH4QiKoJO/H6ES7KOZk/DNCZ
/sRX1ZrFuc0960HbUdW0jdogmBx1IQPJLyW6Kchd4O9z6gKi0NFuYXTq7O9u0f8a3Ha7p5TflN3s
flHL1YxChgpqo7+sIrHOh0TBPATrRFEujS4J/9cIml3j93E9inxucgoLJUVWEbwz8CLsAs6JZd+J
OBZ9kJR4Uk6lR2feTL82nquLvHM5nNtqFfBia85efRTfLu1u/DmApkox/cYQ/SnXg7JESEd01D8J
7jyFvSZrSY0VuMQVlMsMJpV5C+Qp0lsU5qTwecAPoCRQr66xLOXLEzoz6OJQMYB50UjiZJE2Kycf
xCNt3BG4KE/rRX1yNgd6LE8nrieIUZcmhhDKmfxEWnC9EKNNz/nuis0E0o6ca+WiXm+y0c+UNsyG
YL1y8woAOk3OlEMw1ynkgBDi001E5pUag4EvU/10NmNVRQtyvDs1LX6a7qH99JzyzLx//lAyT9KW
XPQmW5aDQztCE+HFanKeW7i0jO3EO++BuxIydV8MCFPIyNqtIiqfmGV47hK4B5MMRbwrKiyDek2M
3o7LLAFQnU/RZRgZAxXGAdFCMhPT2cFuy6QtMORnVznp1mAojdndXqP9LBJ7OekmfpK4otvQWJH7
F7Sn1cN2CwTLCTx9MBNlIWafqKOvQN6nOR2+az3fwkKRWQKA0z6VAd7aGQ4Pan1obSxDk8gU7Ezi
g6KLOfsuuOGHcmOnG/GJusDUA44hq9KKsVHIhT5rmNUWuTePWxsqOT3bUrDAXWI9Vhr3juyDbaCk
fbK1Q4oMq+cpmV/JtDsblTW/H+xuWbNdMuMblnTAj5CywyF7IudhTC9oXbj8QgI2oqE1dRGvdop7
/w/lc0pF1OBHdI6TA4OarUAgnoEAXlKN3WL4jhoLk9LgnLytho8ZYZZIZ/2CS6sxzaeLX/FhKjwy
G3+IAn4X2OsN1DeNuxK6WdxwfjtOtMLb5953vegyeiNpQ/yATnshXKvbHSAWK9TozOsyCBRwOHvL
4LV7MMlte2OvrNyy+86lm7br/60UcvAnFVmt3v6FmE0k3e0eKCJJO0Id6QLaspixac2P3vDLN2FG
O54SUbGzxmH/zwQJksigl3c+qy6QZi/ZcoSOqwJ6cT4PU6vSJ7NaA6v190sKCGcHN8WTxzh8BQ7K
cJQVCQl81SWTHz/wFRpqE9uiBQFsVeWLPc86owwuXt2J6lpOPyN7EtccMROMW1KjnmGn8cg8XWbP
/BaI72nE3SoH5RuRbHoM8wZDsxRorPsOw63i6H2RsCJohY5PFhELSJ5J1IMagm63DsitQ33AEr2H
qfurSHJtMxsRSRVfKPxsPAhgZQSh58dxXFv/zSNfjqRG+h7LlZeuquZxMh/sCG2JyCewj0O9PX5G
kgOjqcmUq8np5KDruUnVFMcdKW2BXUJ3HAsu34l5PJUU2gTedVAaBsZC5rSNzDbhe2iUrUiik/ex
SYS5jvLL+CB6FdxOBz7XGG8THvxQWOWHM6bYh6ORFDGrX1TClZxFflBjYO6goFhw7nPCR7GvMHpr
Yk94uxS0LmAM7TVzUqRkIsUan3xVcdnV6w4ynUV1ShuQrbJIT2jlEQN5VvTXaMQS8uTEd2s9lGtT
21MyAkW01fBHLvuX7IzupSXLVk6yZccdaZ7tB+6JksAeQJbhn0JvW80mikt1f31HJN7i3ZE8bTb+
Lq9MFqqkVGoB5X918zoWK3RPX+p3ZUq62HXhk8lKngdTu7gNsKx6QOVzVCmQy3idFDAFFq2Hhm93
OyiBVsI13HWdTSiObPVChWAkxZGtlmhBgRde/AjLx7FGOUvtlHzUIbFFDR+r20CTNCqLokMrGVeI
pFo5nQldfKWYYkZI6DxPMcYoQG1yZpMCkwv6pPXJ73PW49l8UIzzAP1RVu7J/gYjvriEZ8n9la9i
zHqoPob2+V+19ltsB8BPX2umIr1AVS+edWUUO2lcrVowE0f+SvHzSEyo+WQhGK6tEHkJnXMlZNYe
sFv8xUn0U1IKpQgR7eXP0evjZhsNGAC3NIQG4pwfIzZTvCDQVmRWWh1fsgeDAwfS7S23nqxIx5fz
fWLZGC3hT8bd0yfiEDiJ6ez0KSRLt3nTwysE1VRdsa6MMvxgjftVJJWDw/iJA0NE6+yDrYi5OWlv
mXWb9rQP0H80YF4SFNowHESo0i+SK2YOMx7zYTCAtfbrOzRvtnZC1kfQXj+0GJEE9Vw+73Apf6lh
c0bpqkKnaCAjKftcXN9sQh3rNJL4ldzbfRsq+YeToqTi2t1eX7N8HI8BYYifIkp6ialwUfREASNo
dNlTnGnJhT97blnYo5Yx2/SpCuExXXPeJ7fTWckHKplms836FOcXHjMaQ24nNESItHjw8+cVq1PT
SqSZ8uLPb67rbQkSqGZXHWw+ItUbghLygTdxp/OmnqUIEajBOlv1w3u0OX5Tb4+BUQq7YbB4Li+P
lLyP5CSLzGAYbAWfjF7Gd7z0Ug9IBfcPaQs/hTdlv9zlzHse/j5zM9NUH7h68Us82lSd5rsYJWvo
lCTylk8BSHoT3se6w9j6gbQBg9z+9kFHAuSbEeNCaeFZ0YTB5gzGkBxIWObDJw29zKGK4hdanJwM
qe4xnAjDveYQ0jZPkmyAmsSQPDs+BpbCFbjCho+LFXb3UpdXRf/hcSITIczivCHpDLSVus9U2Tpi
dskBbevQI4dZMiLBjSK1gqdP7MXBE3BUuTzyD29UKYeTmHiYXPOSbkWxrQZc+uMqBumcnamnwmvK
m5TVq7ooOpP1g2wAIOImFy/882Z0sJ55IguSYuqtqV8RMWPs+ufwLtP/skc3hM2mkizO7ss/WtO7
4tF9nFZdqw6Y7kFIKMT3H/ztuEA2igyZ9slnT5iQVLb94YuwhPBuCguYNcNk7wDE1X8u46wkRE0y
r4WYv7sbeTieHfzW83Xxxi3Dm4Ip/JLR2PtKD2S9GbS9EkP5lmgH514uGfmNTsYgcWBwiYW3pevA
0mAMM+5M3onp9Ostuxq/dcuKZKnJe9RONPyC4W96sEQU5eyvC56xBofIXX3I65tCWvtnn/2r7LUF
cfH1Fav9J/EJ/dW5n45kqtNn+rV9UpGSwQr6lZ2VfnjFwzdX9k2iokip4Qt7Ftku148cAgIghdGH
/v6EiS522r52c9fpyB0AlsSS8pKUm7/7/Qhvs8yCjgC6lctNYArRg1W6Rxq98WU3zY851XE8MSkP
Z/EEQYQEyl4EuBuiXkwc9T2x4UpQ9CE+j/+N8b0Co7mTdbFy79ASSBFG6xyp5N3F7Mzab+frP4WC
hvuVk3XwbAjiBvtTAO4P1bfCk11STcyowo5mvXHwDKlWEaM00NgqVAosCVueTPbinT952Xe9ZumL
9167MCnnKjR/2bIk71a+Bx+lwzy86jwckcstAgHa/C2G/lvJVy4YhAzcLTDqmHhLkK6+XbAJ/9Xr
uGzmPZht91YU5J5S3uY8LBfKq+mdZ/xk5Dd4cp2oq8Gpv4BUH/tWliL6h6QbnHiFvC80VWKDO0SP
ufkIiwW9x1Bo/kQBePEq6XQEa8+Br3enZkY0Y59ahAfgYFRivq7Qp+ePWK+XFo+J16PcV3dq370R
sVwcBGB/oh/9nDnQ4e6ThaPztidcXUQJieo/N2t7pt32tUznAOI1SgxLZQ08R1wmUN77QDzek/Ay
R8LTpe/PISpca5G9WoJsSI0+qee01JJifzAmjwBFDhkQ1swt5LN/aKrZq5LBz3ZZyBbrJabs1rHa
oQqJs29rJhZ8DkLRi72JcLfn2EgCxCeTvrBSkp9pvvIAiS+HIXTL4CoI/amX3SrJN6SCbMs10g1h
4SA8zJmm9qe13rqesUWeNOV7TAQk/kTyG6dahWUzBAlGbMjO6+vPbq6z73hLcswZJVscDfUFB8Qm
x/j4HJX1uTtZdRiEpBjwvAX/VvFAI8xOQ2f6Wsh0o3133mjztZwQtEfN6zqeCyWZZrGoUBmaD+TH
AMoPND+9OicpkVXMEOIKDahVjf0tdyctgRUXkzLPeRzTyWrV8GU0X0btXc5+ePzgb78b2hJTgOPM
1HRyLagMJZ/Vh7lWbnJcqxvamWHR/j+t57QOX4lOqFxo8ap8npGWWMbZiwwpZRbNqK6eKgiv6AkD
eCLO9E6gyl/9v7w5pJjhWco0QCzV4OtEcWAnvc7uvtkffrfxl7aw/wfxajkAbH6tNWJcxpXmtTkB
xaDVRa5y762oFPg7PbIqpfKXtAW3tOzbSdOK9QI9kWMad87S1DFjDidRWFq+BfBbN/Maag5TQq2w
Zv5iZMbHaElLpEPOWZGgwBORr5xPlTchUYAFfhmys88D+i/0CEEAJHRlORTi0H6tOFgo88qVex78
WtcOJRc5otc8Y+VJNw/Pnop7o9egsk79HRESACAVQiUVbUamBadzG1Kuk4jyFqY70xzSgca35a6f
01LWivZdtHQLuGJ0n1Vc6mDeq6cuGt4G8nBk6Ab1PwuJolLoLC+9h4C/aLAUjFlZYZg0LFMqF48c
C8wGI+7JRTGkDrLXI+gzyQmAZUb1RbvALvB1agt1lK6789853kJXKVbDjyWNgIj7S74O7ErxgpKD
VgicyoAXHqu5wKj94dPnqUT5gpBQBYBdPyCwkyucCeTc86NNrN8I/pVW5xf3p220lLnSk6BNuiJD
6BpueI2Myk/Y2HhL9S5+aRJh/EWCDZF65JVA9mKcAg2JZ19UUmggEx1yQrioyRRdcczJpcr7ihRB
RB1IgwojT46r1kTEt8aju5HbjocBCI+CR0sW1mhCQoq7AdVLX1HOd3LX1ET/JylSWosCR4ADadUt
B4adJyrt92eqoBMUGWH+6lKfLqog7Zso7wgi05Tk7EbEZeLd03btpD4tgo7BW0vcXEAVYmnC4JYU
57ElYgtQbJ+kXjhU+nCdshUktN/bQDZ2tBPwySVIpfzBdReQ9ItBDfwxR+bM2vcQa3gMoc9HyyAR
HD0W/dl4Dypn9huuVONs3Q08azDknTHQ8AWWnKMjHZmLiXDKIgJTBGQywVhfudwS/lRFR5uQo4Gn
Lh41knSHJKUjJKDoYqOb8BCT1Zjwix31dZle6cDX63tdZxbVF6zA61ZU5Lzfon/z6rWs9i6YbChi
NK03hiOX8o1lVsPnqH/O6hLbe7ggrSbamFy4ospiPJKN3fvOUn3W38PHRpYk/7zZxpPrllR0Y+rg
akItcwTpRFgsPRy163/knaWGdfSW8VmFoF+AaoALx59ebOXrc7h23NS+8cMXjlicuyci+OkG0otq
tZrBJc2Txwj0x6lOu/3p/xO9JeIpbXZHMNrE0Uax8LCyNkC8nEuSCL/JcPH3pfg/oncNkQ2wyBk+
hZw40eRKGBnyZWgeRLku3XaSpnjnP96DT6WwWku3z0inwi/65m2/XeO8gbr0GuBzo+kRi2Tjao3G
n42mvXCoYZNlj0MrnCimuKl2FMgkvDAlddDU1qPXIkzuA+G1QX/Nic/Z6VvhCbuXi5+m4d2R8rHj
t3yjQhXcUCnNKECWPJeWnoLP/vxVu46j3jhaOhhMyQ6qDZ4pfg9Jhy/JjvPJ3e09zISy2xOBF5rh
QHGE8j3ZB+MLN7W/HV2j7P7LEKSRQVCkDvS9eahpy9DHwmUvyROM0T0iNP4VyJTNh9p90Q8xOAbK
J9thg7pw7Jec7SFqf80TsHag76/A7qJ5dUAsZQ+pP6OAhNzR2/mZfwMwWM/La7J3PLJMeFab4Wi1
5XMvaljFNOKiyGw4ZQuqQJwpklMkzNn6tY1p+LrN4Qf4B/wjCM9mz9HefYIX9pqGuanaGk+ht4WK
0xRwS2R7CHdD21WZfPWp2z6toep6/DfCMaBZSqI3y05xg5dqFoPmwf7M62/LXzrNZr/3geic6ApX
5S2A3DIQp488MO1gih7NIFHeubLZPJFWPBCxQaEirQ9kgfqs66Dp8fspiBXduTtmCz2+5BA0faQS
/rkLJ/IKqsHLKcvDsAuULOFTOZnXZO0W7sm4yw2nuwkNbshespCD+QKWbI7wjh+pcj6R/U/dxH47
SRoE7H3FT4/inCmrxv7vOp9+X7utGICr2mEtWS0rZ5bO3dhrr9ySaC3LputiNzEuwuHqhQlrIygK
88pksZcLVwFqxo6a41/NcBMkO92R5+bJYj74wQkwm+HjUGg2UD1iy+3u2sTyTtawcnBaiIy5zDdD
LYGNFPs40JC7pMrlVyXQpJq49yap+xjkdUfrXjeaf4JcECZcXPjl9s3GSVMAQFNUaOzxbjAhnuXv
fftnsdBOS2cTZw+NaSU0WhwkUp+YAurKfKLftvJfE43Mq2SXzfJV5hxi5BY0xb+PKijXeHBPVOgc
Ywj4UfTYbMK8Vud/qMIB5LG/zGkjcFZKRuFCIHgcMH74g6vXgaVLuPgpsl/xJJoOq18SsXX7+dEj
CjnwWY1E178R4Nh0lGL4tpudutph4c8tgKqL/lT5JJ8fkcmr6doN/UoT9vCkE14V02QDYXhLbrKg
97o0tXtj9Lafjfq97owhOiwom7yFzuUqWDVfyRiVv7IALmfVshQ1Smzqb4zd06DkCs+To2+2cGsY
Q745kWG+L0XTtyF37BHwjZwrIMEio+N7BwKvLE8DxQ7jVvGeCDGijVebbVMUE/NQgWoFv7DTPPwW
Z6Imc69IEdk741TAuL4eKBvmoebyI+Gv7z4ml+BY7jiPQEfH/NUoAcLdlJ7AZ1uGt9CgV10HKU61
nBEH8Er+9jryoY7Gz8hMOoOjRy//BKrNr4ggzMSZxmWOFH+Wc2pHO+1QeelgEqMRDqvA8dGCdE40
qK87y9FJSNOYTpxP1ebz63tzEAjvckbDo7K190PeJA9KDHQucbYcb7Re3aL8Y5FH6zDwXfJbDekq
ZaYOS12K9uiTyKIi5CNM/v3INgWNy/l1Gs4XKDMAa0/UbjaeOGkLoG9k8B1CzHT5tXCIJ9SkCJim
BiMtoCXcHrsClwLEywE9rM0rExsHikaRTGeuPaJu4mB6SI9y3C/mhHzB6aM3JBkQ12LcxOpY0LLm
e3/5jOWHMDlI03RWCTKEX4Uw1C9mwR0bVwqN40OxGAUqWxtongrJJ8mNEuurqB00CrWcKAOCNGR6
R9vC9BwCToABXlVjYoS8t8u9l88RcVKFY78T0z1zRyI1rsFty/j0MwHejrCRKeqJmRnxtUpOOiEx
VagNfwfpi+fSBRlfcC71eC2qzwAPZuy/gS8QIrH5x9oT++qy+YJp38XWbZMO+53T4hlBDvVAcMVt
62GxGR1V1fibVomfOcjzbvxvIqhj6vzDH4hvMw6Dlf9g4i6G1RESOeBZ7iq4paoQFqxExCcZcqSl
gLgR6XscCA/vsl5iBzT479IT3PbiDqIP9yn3fbeMCIiQoj13JfniTEUXPqUIiaPEhXBVsq+slpbz
4YGiZVnwEMHD8eN6sJPqQ8QjtVxMR6eh+uW7o8GltgUbh1/mjWel9gWPvh+YJIsclncoDSdN9vn8
8Dicch8PtPxoxDseSY6apSqBVASU/hBFlbI5+9rtMzfI7SUiOEpVjuc8n14z9mbh2Kut/6hZVrcd
8SRVz4znwv5F0nOuVBa1AT9FvqnKO5RsU3yXBdWuiAkDSmq3V2cslo3RYuYvfsoKlZV5so8NsuNk
jNdBJ2BJI0dU4qDEx4N3tFLSJJrnUztz/p0eqq9fGjWqq3g4MHV6rqjmaV6bYxdmR+sbonFbkuc4
qKl1rnJLL2sXnywbhLfkTD4b4J8dcc9iT0NB7XTEKp1telMbpHkZlW1W37WaXpw5ut0LBrT2utHj
5UvJ1bPRJ+esoWFC6VhP3NwbAEwE/QsEdzV8KQRbqgLid5BllyHKyqR8OktuQt7WCwlKf4tsFZWo
doU2tdDLS6UupMUdRTpfUl93YZkgSSSEywNFblvyTAbORfAW42LO5/8iuwh7LqhAWcSsmBflShWT
lMgYrFH6yA2BlobW64GK0L4VS2Q1Ri4m/1ttwYse6Jz7s8rYgzZlTDMHzroQR+DweWLGf/l+cw4c
BmWltA7Fw+h3BhIYAYsNZw5UYquj8BAPmttbvXOLhc5xvFYEi2dybvm/IkKzaxb+0I/qvtRu6+M2
Y7w3ggvmkO8jWfJ79bOj5qTiGndJfUfXHfcb3ngwtiB9R7yDM+6UrQeg5BxLc43p8w3jLDPExWNd
qRE3SHGNyYo9mcpLb3lpNMVhPRIBVEEaZ+IrDRK4TF8l3MbrSPPv0lPyK+o2ixsW89mnPxma5rw8
77511hsa6Rzf1qkejx0vRql3GkGii+qH3T0LEDDRrLq0qxPn5JPcn6ac1Ek45zHTrqt2tqf9zFdX
os/JqoRBwDWMUU+A5JG6Zb8mbcTiukDuv1pjrek9oj1rbf0IbGQELz27u4uOElUuTYqRUupN836i
BZtHQbZpdq6UGo+pZZrrrAs6P/qCgyb6FIINYCjCPpynuHhfWGT6EUyN3kuEqLbb4q9KY+QClARw
QESzkb6ogYeyTyYYIbCgvmEChlw2+DZDm9W8KvB0NbuxoEFIPOBqiVVe+3wht7cfSgGPDD1oRnM7
Jix1XW4FNOQlyQP77XHEh82DmebxcskDOXvXF9e02uu2RcTPH2Ep/SFWSG+sdd5MDPFb5PiRxqiG
BCskcee5igD44Haz4FNxhCTpZa+b74WuZ+tjXhlHGymgowsbDmYafItl1lp9kC133O/lNP+AjsXe
qp2EsIddiPIahJXwXG6TI8gfqXsKMmHyhesL02UdJxHe0/i2uVW4erl8Ak08v9L7ywsydpCWAxnH
u9lldvwu0mpX6X2DwP1KQLWwN6rsCdiQsU12yQ0hSpVe5Kx5dydhJON3jWzCnUkqynjw+eqMs4mK
GHVgFSEI/YMdAMVA5PN8h/eKYVcNeZJW6Brn1VD9prQZ0cOzMzSIqkAqhaQdSx91re4t5aly/wT+
pPjRmqgiFe7BVb8/IoXcE0vH0OhNFr1dLy8b0vYz1ai4cPgdfrLz57w7lyx1FO+zZuMeBgepvBCc
yuGaD0LBMNvnuYo7RNlh78wNBWq3hGGmvjevQcgTcQ5ze+rKi0hgojg6C6hWLzw/eBcNajaCcI/p
KGk2Vny7h98jabC6VFOVymnBDywLjTobZwfO+O99czEgZAGlRnyyVN7L74qFRn8ksyp/t7qEgk6l
k+v2Yf9RjJw9bB9sAJQ1jy8kLkd2r3Tim8oIYkZiL0HYHiLywVPFKwbJ4gHuj/GTsLrxTVhADM7s
SDxr2BtzY6CPq/qnJb9FhywTJomWW+zSiRv3MeugCAs45i6Cmj4Rhmp0YeDwXOgtCAYXZPYDaNZd
7KOdpoW7YQZRNEbHdAHZbLCfWitgMOW88WaqNiQa1SACTOhBTMaFpV/wX5+7+SV9MFnxtNPsf+Uh
1yqqHDijqo031CuGYQLb4keVddg00cNqZjdts2rVF1g/Im9m3TFdiPXjyTi9ahUjAGqnMLe/vfKZ
78vvBtvwoAUSaOLB0TiecnEnGP6Bye6AdwsNXFBq53N6aj4XmOLrZtEtBeyTd2E4xsqlh4l7FTLt
eS+a7/uJh9Y4Urn3g3d/yb/uqNrm77p5RnSH+kzdzs1NHt/1rBIreVYMRNHnhElMFOIQSBAgPWb2
I0fn4gP2hqSJXGVTbrjxadP7GfzoL4WSOWYCH+zzuxgVf9e1cQr2nct2n3BKrecj3H3cnHvb2zZm
xW+8EZfbVy+3HI9A2nwH3aWJo/i6zC9Huhd9tEk9YJfuSA/H163/kp8+uEQfLeqpdySSKzEZeqzV
qNkYKc/PrT89fC2xMHdoUnKBvb8gU8Q6xrcskgjCV5D40k3LjqBLf38gG5eVVfyP6zZadB6cBkhN
oHPC9anZJWrYMpJFvvMBrPCuSEdTpGW09eDZZe/0J+fXip44ubNO8NM7IuLlwbYw1qR0EduafQ3m
G3NWCtkn4ynI9Y0TlfWBUeJKcqbB+H7xYsA/OSkqMUCF6AuviUgAjcyxyzWePnc2YZaW+UyDC69R
bWHjuRBelQ3AjX715MG4/btWtnm6xn8dZ/qidODIfEWZRhCJz4FzC1bvkoTDWysMVPV5BfKiyXpw
dtD6IPrenNFt8163iAbmdfmb28LAJ5+jpaqoks1ENxR1sP/3PfULSh8QgxgrTX9v8igsGDOTjCxD
l1Yvke8QdxzyWg3PZsjmsPa/ApSVVvP13C6NQMwzZIXT+mpwy2R/lcW8717r06E8Sz/3PGfqplQC
8ZUWyP97AVsQtZ+dFPM4CSWZOVxmn3ajQL+3m/OQ715f7zxljBgl3gGNb3nGzCOfxM7cDXlXohZt
CIE1l4JsH4OEpW3Q1DehI62BE353iXYeRA9n20UNyP+3Kp20Bb4SMsVEV5Fk2Bknw+LfUM460yhS
KqeQ6yU+cjORbtgWmTHg6bPbBtALQ1ty8Rr01jM4EUwgDM2TUVo55lv8XxZB/PEn4cIDCIyPgM+D
yfMKTTGXZLLtkD4V9Fay53BBd47FO/1Bv6CuxBjPHuJ8MJRq02V6ueBQ+RVK16N7tisW3PWGQ1LM
LI7kWpIFV57odxmgmiXP5KfFg78felyZ7OD1slRhj+u9+qdiIIjybEZOMWIGiUwr4S3PB+Qm3Ezu
h7Az6oUnlew9pctEMQ8Iu56FuokSa6Y56lMVrkKKme4fuu0/qK8hzW0KYBJeTFY/kviwrqizzoEG
HEYnWL8hveWMxY7mXq8YiHWV4GoFAISqK08dUxvI0n+xRPaJPp7g4+Snkd7v5gd1DEnxAy8cu/k8
ZCQniWfafiR7W4+zrfT7OyaaZ0GbSoS0TGLcCSbtskqHJae9X4J4WdqvMBaUJxPl9C0Ae0fffHnd
vdtg5tuara+e/+8USinBcFlroayrMm+CMd31yiL0lx9/iGjBiJ5T4aTp94Hvl6pUBnvP/QXVi7HJ
Jf6olTKrBlZhfxjKyoRaNdrWrk9FYPUk0EIXqTk0VAU2z6L2Hpt+TnRxUNwp66dZsaKGxCZ3Ol12
niOlTtlQVW7idQmLb1F9Sann8+6uYMDqZewekmL1I/l0x+5vCrwoDsBkicpr+qqt8HfvpDTOx0Ld
w3PJY3AAZcUNQqKOOQRbmHFyQKVTtwokove3nQ8Ac2/hNTJAyoyffy2Z82NjetkSl4sqQ+xsWddE
qlPjddNZCmHv3wCR94hCNfisX6o3Ch4DE4qtbRwIX8MrWe2IR0SGUeAZDjUfMVoc2zzKM8fk+8Uo
Kwe9p6LeZ67LKXPyUBEZHeOUdIFHutdjYb1NIzp+R+34KC0a/yaPchc+foF/Lw++KPffdl9FqOAM
7xeQgO0SQjWQ+N9Zgq3nHA5lLW2ZJGM2NETXzwReiCbaPZ4vFd9nERtxUclMtCEIualLFFy7TJYP
SrDU9BmwpL435kaUlPvCCTpMy0E7sX1Dkur29kiF5F3pWVUuwWzHoZBSZXOagO6uEqiF35LGwTZ2
Ou+ynIWZjCIZif9Lx5scwPv+h7ikzJO4mikBnw+fYkpA4Dsu8SFMUpq+bPFA+aQXn+ijKrYa9NGK
02xj4XsGIT8UPMXDGrkkQ6BK1NpaEmlujXE8wFTc9LMvdXK9g6rgF1sytNpK2TLBx1cLGAK6/lGe
sxYOj1V3lVG/HffdlXnTnZIHbzxn5o2sdQhKBC6a6xPACIZRlLN2865+xj0rLwJYeFMy3PsOyKkI
7D4dHPajsamnFyj0UTiW33QjX5ybll3zS0QaOxFH6WdowP7y43azK7l1JjXQu1Lx+sRayBa0tLV8
xBa3hP+pyPEKa740o7/x7qqXlVfiA6gl9cOqgflyegZMLRmEOg9Urtypiba8q1O3zwfwUd4YKwRG
Rt5MrsuK0z1PwFQdQzlVFgUD/Yiibv9OraCjqk3WOQAXzlDvaRy3cgQgS/2lSXFuWWT+L6I6KGeF
96JbzyOoE62f92Ondmhn7pN3y3ilOdINF3WhWe+yrKZW0OLR0fifDCgiyfT/M3drkAbGcRv3FTRY
4Ba/f1GH3k3A2E5JPHpQ/WDgjHVaJisLtwwIRF5SwnzkoRqI0SYsKfKiVhqpZkye+APMOuRgS3n6
eKP6nMo9gPS3ZBOToD9o7ZJcGgNadDFJV62zZyBRt3tmpzjuXW+YeHsp40UH2/GD+fA9FNsIXrlQ
NqwPm6ndo4TA32vF9TUNTEn+1wxnAb/LgNmUujwbl8zqyZKe5EgNNDO78G4JRQGTuTkq+ehCILJI
7nVeQ/W/1C3MsfPariFG9SAKL6RuB/eZ8E2wkEMRAzhhqGYb9TRkKZxt2A38ferD8rBrLlpmDE94
i9sSQ2J4Sy+l2ZyUhrdOtvAL0X9RubSO7LAmJr4XwwhSPJBS1+lc5xT8z1RjEMtPWLdTXrRIofol
yDo8mZ5m9y8ZsvFRwawG6P3a7KOKKQFWHScna8x4z0ssqE8+P+Aop95WcT/xD9p8PmmppWnrcIjn
zpYC9ANsYPy1Io1MZxTDFqKB01fYmMENJQyeX2ndpJPtCRLM9WfKUVqSzWJb/ew27NQ9/OtzbD/d
NqNYAtfPGapaUj133+Mn0PzADO5PEU9R7jc0JJP1aWvKKzUUAr4Se1gv0L2abHP77hXLGSZQVT9c
Wnrb+c1FYLRpTdF38xiC3NyhUUoZt9uG6ewO8Y4NPFLXuc/EXGO3ClhuNbJ0Rg8HYz8aHNGdwkFV
Iqj/HH3KwPBT/cMRSHyr6G24dxq6aqTXyBSToLJepCC9wDhlaMTPGIs6gfJUI/k8upoiPBTO84Pa
Fvpjylxqhd1Z4AZnh04e8C/dw+ecTjImurL8RwimGdDa2ePXLwATLDzdbNr6xVz2UsCGKh+cPlgL
5cHvGdOiQ5ZU5JFHq6J2g4cb2JGL9ulE8Xa/rowLwjYo6oMx9fjLAEop2b0pkygzyx7YRfdmJknq
oVIyPpXnzBbT074bE26lfTt46QVPXwsnh4DvTKsUxxkyQz699OziuOGTpPAFDVV3jZMWjvP9tnTZ
0lY9dpPSBVuWra3dwq0De/apmw7D+J8P5oyUFG/obsL8KuFLqUyydwqf1XxyTaFrYwvE/2acomHR
AMVTNfmGcau20rWM0iG0lXcyt1Tymsu/FWu2aANbGnR8mG19hjHCkokAcgN03nvgj4ctNY9EIAfm
/S0NVUliND7ZVR49O9L5nrIbNAWvbm77YrwhDvQK2BX0rsAXns6KobgHbOEp26mf1u0bw0RjtRuF
sYn1aLMgnnlPxEsFmUGMjtBmtlKfRsV9t7+Lsu8WXEydKan8r3gsxFTrzogUgRsCxN2dSwxG0P/o
iwB+wJSsJ1UGneuz1tpH0WxjwfrnyBhP9oCJ+diIVx89tesrn5CcDxJm3zjs6W17wOJUVvei899n
22xWrn4XMlB466swqxB8aM0Vb5VsK91yVXgTu7wak2EUue9ppDylqYrtDEZQh/pinPwZeqNyz70g
7m5BkWpDBtuoMHv2AIdwJ4OvCOzATg49vahDmhrGnFQ2Sl9NUeQcGQVVBWf9xE6BWos1YJjpGGN1
0PR8gEllFXS5NCZtmFHPn8tE8js1Twhp37wA7FCgj+W8amsxW3w32rh7vA7AYgeQ24CS6A4c2KjW
c3p1H0Y0F78km7t6gL3s2ac3FjctePTVdAGPaXUDpNjaV/ycp6qTUyoSAyf9+2VCENMB8zNDpE/z
WGPp1tdHMVWJc7blg4XNbnmtg20RJ0G0hpdwI7a51+3bSGdULcprnPOSW/0UQmKpoRf2PKoxF3Al
DMcSsCWI/m2Pbov9r96ofDKs2oIKIgCS3uVb6RLEQNOr6n8h62IIRBbrgYzW0N5O+6mGhjTrLgij
GMrV3039WPl/uV+DUT/EXDNKU7XnNjTELmQhJn4Po0zlYPjpa29XQjvSxu/UZIghl2wPecG7Krmk
aEKHeG+LoNPT2bnSASJfwwHWawlcbE1o2om1ZhHLSHw2C5PXNEt6oDQ3Ot9w2zqkYDCalzx5bLtZ
OoXRugI1iiP57LzviCLEAP46c7EFDg2J81B56rc54ZmRnWLUKLF7ba5KkaYkYjUD6YpUDF4XD0hj
XgBUC3ZJbRhcNzzyz2wDxg58ENU4BQTWIAzeQAm1DASAc/61JejxDmzFTvIn1v8rKBjv5F0pQY+O
hmIvYeUBGRLWDlfyjnM/wGv/viFQ5YVfnM277/L8KEhtF2NMhmV5x2pkuxAU/dnwcoCQ6mHY8t6E
Ujkwv/tMKEF/OwOOouaA1yhsQhp//ouhIRr4WZoYdjawbPkmC3PbSOIPidgsmc7v9DsFLedqYc1j
9epGsF1DCseDRZR3KalYNJxK3ZCyFnDC/5Vg7aPAbXypZIF0agPYVwGR/FLPo6tJ0IZf1bc0WTzM
8Q2DbMv3kBhn+xPELDBPl32HwGsiDuKI2haRBXnpy6kaBu8J4eBtk55gawEYZoYwpQmHzDE0e/8U
fDyIQQP9kuzldHO/1pul6Bwy/ztfWuPu+xMa0xC/pEc5p81oWQFKgVR+IIDizopBTNR5BP0JAnkI
eo0p/ONQ2VM/Xnm3BB4AVUqXvCjtHG5PtXoUYXJwIeNfob03X1MHXoCj3E9+U3qf71mQW1x8F73W
TuiK2q7hYaykpkfh0uEjGGNTSvjvk6MlO4i+fifA+eqo4kZRv2jeKkCIGlS3SvXkgDsijxTLUVBJ
oBh53c37AMlwtQfISoWcBfw9FfeVBsnGP53bBM1qjaAdkePu02eVjKvHJJXpxp8sgu1LsJCri2Ge
FoPifJTDLjV0HM8i9AiohA7hp93uHONtO1jLYXMw7b9M3bH9bndsCtLQ9rBYFAwMk4tFLmYH7gvH
uy30ya+YERTe/Q0szR2rW/ifbaSphsmExichH2whtyd3A9+GyikXLBQUHNR0eaEZ5gwvpc1WhtZa
Bz+j1Wc3eTESX+4LFUs1l5+kuMX4vEMptEBhROImQAzPO3B/DTa+mC4OxG+3A6PYn4oquuHFj5zT
OmquAqTY4fxMp20lbP0a1FlGzlABGXmugYKgPhCUvTXkqUx6JfR5L1GeLtt0PEmTRuYkG9hhLOia
3QzKKMmAREAXWDKfKunrSdW1iQarP9ONwS2a0pKNK4wyHhUsROYCPO/l3bFZULfA7apRyILpTh3x
82+32S0XpCtpUQElYJTEu4IuUyilL/raKoh42pu4Ldf4BIuawPF+W8LJwKDwmvsjgw1NfYbIZ7hF
nVjfNUNFVoIv7on4/pP1FREdgVyUJ8fRqO09sjF1DKJ8CM0puhR0LvW0zhTgSkpXnRkXodXp00ji
wmIdDpAD+/+yj47xwEKSXaqfWGdYyDv6WVGk0jWClEV8YZzIzrHmbR3be4La60IXk5ZhGTV5SL+K
D+npCXg8awGLFmVTOEdquHR5YKhBStbjhxIEDjyxYJKU4dIYGGbd1TRo5YA1m7ts7xRzwGFkBnNn
r28buxQ5KDzg56YfjGn3xej+PWYwKhTcNAxmoXIIN+a2q3YDv5gjdzhm0+SSulCs1RFnTJbNwSbH
DnxuApGngqtoaolqrYvK3IQZWyaCtxUu/nPFPRUDSI7mWJALqR0rrme50SAMep0+5THTfDEclytb
tDaUHjU7ISp/GtuZL9jxIe9a0TsG7ZPcpmkkN1iO01hgPiZhLym57Wl6jgIL5XIBbFgZZvF7gFYK
hDpkYfFOQxjq4tkJxlUAMingNh71vhclXhyIdgq+Q8+Age04B7XE+5QyZqK2k2xORrInlUagaS+q
YNJt9c3PRuPd2NSWbKqDUYf8YZdoPgq6ozBWxrQIy1KWdn2GKFqNHnx1ARVbTJsNo2ePc4wHBjP5
/4nFpHb7uA6pnWKOvDvyGChQu6g0gBQT8FfYgVw7eJRcaREtLvCZ8G8NNR1XXrLeMZr/2kgxXGfW
zhuFIfSwFzgJrgi9XqL2wtgkFjUMm5IqgnsKBV5Jmrt8/cfQL5dTCRNioQQmcvRSE6o3CcAn//QA
y6zTjjXoultkkPj5MQP3MCc4oZzx+f0WDvZjuErlVXf9JjPJf/VuBtNgQ3ULYXm/9bX3ZxFZ7cKS
/7lwulawLMOyXqK5pHEg5T030auv+WRljCnVtsTG51X0zh1OKBFDmpK0RdTPZFqHeTRy2xl6l39Y
B3d6MLDINU50mAfbsFh5OdARwDfHNT+iFUGO9gM0/od/gLgkTRXiyNw+LVkq0rDtZDj+CWB75tar
6Wa7NUrI+6hvIITn3Vft3BqlLenwcVgESH+RaM7cGJDeWC8WjZFgilqrtWcnc/RdJl2CzsXWNe/M
DaLYTQzr9pjvtpUI/TpNNmiL+R/Ic4UfGQtDFBg7e1g3i/kAtfARin85GpbNjZOzjNAs/Bco8aZX
BWoczML2GjYEBljDVb/MBnli+6WDtvqNDHpQ9brvjJeQvbZaD47OnXAH13gyY+B6q6dOKuy7cnm0
SOXCbEy/RX/Jd5z+XCxUdDkrojnxqKcxyiX4V4uBwluAxnv4+kjdUZmIxOD9YUXPtX+VNQj8WjaC
bSwtCRwq9fQ8k2Qwh/5agLsLoVkwbkQ8/XlwismsetD0mkB+2a3bGkg33xyPcDxY9u/5u3nO+HrD
AFzB4uw01fLEI8VYmQIKOSqrr4a45MF/0Trh59nKEwtcX4Y4EO1jMSw6isvjQ/sL8JZP0ivC1UJQ
LG9lLYE/R0s4WoUNYByaBz8qOd3vELMXND7egbNZNuyRSOwTAqW8b8cgULbGqlU+FtreglGrOe3e
qTXoMfYufxuIFgaZbZz+VbUEiMiL2cYy8QCTKLmX9xZ4sCBms+JFTCFP8c0KJ9fqk9MCK6ZX88TD
0fmg9ourgyMKRZihVbDsKpwOt1dcpLDfsfCZs4K//iiCRhdUk+9Al1kul9mrJqCr0XE//unL8JWw
GQAO9RY1N+TXe7heOZKwiM2x4buyzcZhKVxlQTrN8f007Ef/NDYR3YYAMQzeo3nd2GsCju0ItSjm
WSrRDufr+9SU0zWFPeaYu2TuKHBHjM4ZbESXrukK1X2w5y6wvwd5OWfw/mehZjeUAyVFR+tQ0iY1
KZeQAa05szZYf9E07MajXIUoyO9Bh+vgVSS9dBTdifjl2Pq5dL5vX+B+n9qtehJ8xRLswU4gagK+
2pCfCWPyyDuLAZHUsnjO/gTKb+EXEmK0u7m5gJ8hsiuVSFkGw3ufSPt2hgpAMV4Ko7LPEqBirdlb
2M/9C8lrNH7vSgTwCedaz18QDVUcu1nJEObXwpa4c5tGzSYJhYXkwvgdYhoZe/qqD27hAYJ9PdG4
TTssr4zbJqzkhefBdVPj78RfDSYOIZ7Kccrt+1N4Mowem8MyWZB7aEu9ldQs1447eXupkR/3Pr5f
lIbGLbDX90gUSwy27nOobhJ6As8zFWuUQ4ObOz3TgdcBDtOEwx1GQK1Kl/wL7z3/rls4UyucYs3f
lqMYfrqkBGGWIjbuf4ocav+fVuC/h5pzQKS/vKyG9yOffKMgkUr+RZunVl1btL2lARy84or0cts9
Qk1Iz/QAWbBt8kjTaWoDPZy6M6f9Hxyh1xuwlt9HjIe595AFiUA3bEmD6UBozA8AHbZOFYAShGzF
LBfLan6X3yzszzptiW+SqYlAMRYTJUEJJEAw0Cz9GFh1nxHu2aC7+ya7FZewCZuvU469VV9pJpSj
qfEME/x2NvvN5wRgxzC/Zzdn9ipOOYSt4I94VQX185D4rXcs4SnfmCKMF+FkNyFB6sr9nv0qTIMY
148WNRtznFKC2GcLUTi2rmrcK6qNO01voLMiF8agMbXNpu3gpeEeRzORXK5/Zdeyt2f0oINRndnV
vFO58MFAnXrneUOgspABgr3ioKW2BCI5gU7yTeHYjY6AiFR0JnDPC86xTiUVOzeQFSHBNmwIFVo/
BU1OBdsPGXxutz4YDK0xIE8uMJUyQW4XKnvAVSWQR9UWYLvf02n9Sz93qvwE4zpfCPEU5h0H1whz
HKNMMIP/MgpKF2CKHisEdoFx/RHEfqk8QGdW7QPZV+uBMoWDxa06HDmygox4ylR7J6VbERpSglLv
ozMAKjlQ1juE+bMtvEtBCwnPbMITDS5c9+ihIUbF/EoTPWLWPrRevk3pbG/HZwgtHZMhmc6+CruQ
CbzzrqqX2UC1CYuk2BvARsBHOo6lIk7SW7Lf1EI1Opoi6XOKK6mhOKtOevD9AlipB9k+9ckriM9K
wYmtWd+VR0chXPVXuD8oCHk8nIRkZ2xaQCz8tnyt1YnHVdDWE7FkUrKMLhk2HFb3xFcJSXdZO1SR
Lvyty6js5yX2gJu85fHzzVKxkbMIobM+1hBcf8Gc9wgZ5ySN02n/h78qFB74emuCsbTvpSRsIUWs
2VVCvIsuEjU97xhZfnD9xXGDRBG8mkOd/TA60GRjYQaqhVPXD6ueTMQg/JMPlfS+msm1Yff2x+Q6
JU4fAGIgiDYV4drqayi2Ch+HXMJ45CRgvCE4tV4fvIWJEKVVvv+VfVmNYLxtMv0JRy6GpHXV32P3
7SjtaytRe62t+DkuKRoosKKeL237pApPWu1htIdgaEP0HA3jvxrL6h/xZDJKOfq3EYAnwybaQWoO
s0a2RvLrBXDcEN9O99sG8EypCPthMrOQzMPJFBh65zZgXUZ1L1gAkGcGHFTce5RfIWeFvQZkNuez
BLSeAyazP52cgpqc3VhSLaYNDbBe+z+Saovh3XoXkFXY22nFuhyl4/DgLBjZSagz8syszdNQR+zc
e61k0cTDfvegHZTxh62maRMWeN5nkKghQVjQiw+L20Ci97pSygUsqkWZN5qRiVfi1Bm2Cux3FGIR
3m1qWxVvTrPuD2/9HdRZGpOS2CoS+DBxyqrS7yVeE4Ro5OOavxquQ2TevYR1FhqaJwuEi5C1ZuS7
a3Nz/rVkHyYIRHFbpMlSJhacS0T5/9HW92C6WDvoBsKFCsCsudB+nRifyMDfh4L4671aMonhVMCO
hSBP4teSgsckLpx7E0ifJKQgx7KvI8bd+E4fvUGDuqnz4HjqXTM5LYH9BUuTufJhokbq57J0q1+I
5FCmX8f1IhkURlFTW4AjjSjN6p9LCNSpqGuxs5VBQEZrBj7FHiZr1qAOBB2sbqq+Z8YehzhL9iwG
B6xG1A2nBOL/Iq4nIOQ4P80moHCLE3wJUZhwur8PAgDV2OCG6hVrCYdXEBFoJ2KuT1O2j8p2B/8E
7QCmWdb/AmNq3zQrFp4SUbTxpB/U4j5yLDgqexqMJAdzS4AA7pOMdU4Fx9jumvaOr6RMxrb8ngmQ
AtnDB+XwrJqxfrgqtSozUxi4VSFAhNyfwSmIhIMS+qAoWCSzLmL/iXUQ6sYsrQl9brBbOO7EQT8T
wTfa9aZsm4OKZLIzhiOJrRa7oHG1ARaxonSq5CnMy/GXxU+yfPfao2U7GsboiWD3tCbc7vKBTbLZ
pV4tdD7PKXWbHqlAFKzuJYWFlyy7EpOCaUQutGmumqFLD19jZujQiq09sunSPiJ9DZ/zvhDmHS5L
3JLL1uGSS17+Xu0CIevDXzrprHaG3VnZb8J8gM69aceOoi23QoI9g44nKElS8fWG2vsCpB7V6mNk
C9I2QYvwvFbqSkD+LpmJIpDCogpLZRsZOQuvCcXRqn+NqWLo5z5x0B6yMOGZTfjvzy8x2mqj2rH3
B3MX/p2x2pWtbUHKNFmoK+wsYIlSuRm5Cf32agh1NXonK5c+QSP4SyZbBcc8yiBbND+3RT0bSamx
qm3GN9/ELCtJKa2ojkW8fYxB/zJSHQK7pj8QI95+Yo3OFIWveF1ImrHfp+aBlOVd+nL5PhbWlNd8
GxUR2fy/HAlEV+oDHlWjwNT+p71C0h2AMOy1vr1N2MozbGqnRU3aQyvN3/prN/Q9vKXZRaIpwEw+
4rLQJuVixGcEOOsAmoXzZcGrW9qEI4ri3N38XKTFhhE1fTMkXWMF4uaHy9ASuWzkPGC1yNtg4Mq3
gcNJ1wEAGYvPAp73heaeTALtmAJPFC+qy1WFG1fXHxzeZEq/9zWxu51I7QX3mqTGWh8Ryd6ql24i
eNINiQrVMk3QJcaru6yaHX5kQJ6tI6IyIuf7dgfRSkkTi6ni6Iis7V9P+a86V+oC7Xv8zLT46+lD
ufSne+w2B5cTNwCWg+pq5lKDd3qp6q6t3rzMXy0XcvYiNVq3Rj4cBXOk5+wcJnFT8SJA+fqzYAU3
6ylo9NOvQMszaK66L6g8P2T9XuSHr9pOF83JFIwxGBZ3rKL3bcJaCycI9pmDkGQevqG4szaF9jAG
zOQEjAfp+aygx1CxOA3V/YmGfas0k34pau66WPUewaA0JEgwUGrdjaCPx55c7miuV8nY/YwEC3t4
lrYC7SO+AXoTvAam8oqUAOuZtGZDnH+GigytXP/BtdNRAX2OToZ+cVps8sDhac1rIXz1Dr9pTmws
YAjYafsHS4m2njRtx+bPyztDo5naFn7XlZJaTD1NHWMSlOWl+JbzxKZWydLJEoLpXRTy02p5GZJb
X0vGZq3p2JQJpPrsVSB45T3pE+oKEshObMs/CdMzgCjYTRJTd4k2OHHrphhbGbaP+pbO9mYB5OMa
yglwQCZnCfYRBi+CcHdcptEedX6OJ5/GQgMNnVut2j/rZBGWhadQTqLulH078zykekvb+NrJrxCP
A7xFvMWMpHQjMnFYQhpt/xna1o7mRTwyCjHEm+LlWmikiG7Hb6CY7YBHFNjWzGRPj8cWoY4kjUsu
keH8LFGG1DXzKBiv7AR7+fS7siSnEFEHuCw5CxWMYkWLTbpHPlVeI8hFg5UYLkyeEAAvSjsB+bir
+k37yvB5yVmSsqpo+e6B/zzTzEFCO2C2Fw2Tfr0Br3+YyMypztAdflVdh73ImPkNflyUkhPcIBsK
ZV+o3Gxm7/IfBT8mv/uDDBp8uyIjHvOmjz2jTI6qYi4r6XzcdCqxZf5/P+hH/g1monWwg6cvTNNK
Vw/Y2IwUb/qjUTxy7ItfzjuuDCwH5BP/OysfSPhGNsoNEf8DdsC9wVgKCMetlkk0LLfH+l0u6rb+
bIOOJaFgmDiuNRkqoX7nrjX0BOAGD1MwNoJxG4EUdix568MxTGDnxp2yR8phrgA4GBHldwvmUmUg
T9xtV28YmEBhcIxGpXsWqxabSTRQ2GnvnqIkGX9NciltwU81HBAiV2K7i0OfDcWO4E9AN4e8xgrJ
6SWM0L8QFhFp8t9iuqh/qQ24w+6L8pHB+kwoe6A2iCXtw86pZzeC/X0xMMqzvVWIRTzN8oMZmJ9Q
b6iAutJitwLxcG4iMzef+/5+Nh+cvuwhJaau4wD1wFTDq/FgMrmCIWpNFzZhKXKF5aDRnjGHf0tp
y3/YWJKbtViIgLvDd8eLJPFitctC9VqRCr4ndokPhItjCKKlEWHW6y8PKN5m9zv6sCT905kPjK4G
36OEpFY0gU1jP/w1DXtue2ua5Rww1+Ya46uY7rUUQiHIzjr51yKCIdVz8kqb/ynrl6/6NdtyASv1
g4EYfWkbkzdUZZyZLDcBXF2qdHbylDS92YYzL547lkh7LHbJQ6Xw7UyR1vjANqClQZFeUzTjsHvL
9qYmZTQPELSU6zw5Sjfp8MqgNPW9RkJmZp1G7U9UUOkXDydoXjdnYVdsJDq7MgcCUr2H2GuwTSDL
u8H9n6LEINHsEoz9PvAXdhNfknp4kUSEtoUYn8uyY2KieYUO8PT9gGYNbzE2QOu2A1tIV6LMKI2o
jfW8+Wg5RIooJsA+yOxOTocY+iLNmXlS7YMjNkkrkMhNK6qRYPTARKnSTmXEpB53drG+a7SFrSlX
OUX6js2YZLvRwDzxPBPoJM8/kUv7FG+wQdsHyRBjadVKMhLUKcUlOczpqKhZs3FI32ODvIqcgB94
PaDtsq0jBV0Ma2Pi7Lp7tamf4JqSk3OxnbqctHs2tBV+xNskk9buC40Kd51xNrE5aRKDOSrQYS1K
RC9rfJ3XEUwA9zg+e92NPoM4WCkjWPjK+UcgI+fFP5iytXs1oQTWpNtUFRPQkljZn6pwjHXuemLW
Q0YByW61vJurdGeejFnM+CUQyZplO6ASyaY1SZfhwd+mkC/FTZOGywOJdwOYPHEkRiD9A2/NKB0n
Pl+X+u7jabMYNNAwCYQyUYq+uWcz4R4whSFZm55iWem5gScLjMaDtuotLmpw1HTwpauF2W1MCDxe
qQ/avgv+HHPeIcTtDn1qIBCzwWInNXVsb9trJY+c5fGB/PIssBgyae4FScEZ9vqFTy+32GMIQDv8
x0I16f6c7kn/JF7ybiQ18B7NsX7SoQi5qfZyfpc5p2rdyQm4qO7x3c6M7R9WU+ISXVrPDdM89Ucq
8OE1q2OertaI1uHFsk0FF0D7MWKc8qTNNcgVhllW3DGS+qu+bozPQf24inX795AIQhc8juvUSB1l
hVqop4y7s4bWW3oYbaX81/AxYwoot0jbWhkezU5425fhStyuTMGH/glNf88NnRSV13V1A8y8SVQc
s2PzcHfZrw6WC8qvoQLvi9eKyFKe0WLtP/PuXICjiVbL8J2laIBS26Q61bPLY681nCS5jtr8DmBr
VNxbzQlUk8EO8tP0RvYtDvQJOyAVX3TJPpgnA5rNvkG06AKd4kp+tH3lWWI8axgChu/0sSvcP7rL
wMsKIxaiRO3q+Ck0Fm2+Qb3wMKratzN6lhTbw+BfPptAWh2g9EzLmvZCdL6KN+vGN0zT3gsQbN5J
nAyeCVOOqxqcH3dmbmqosYqec3iHQp47OxkAUNTi05EqHWJVS3dz44V9qZtpXhHDOPP8EFWhFOwk
0gvuWw+zrYkG6KECAUcilxHIQf5zcrMp3IGQAdGJKu5Ydj4v2892WzHq5Uhqnt7BS/N8tToYx2dr
cjgCqgpOkbnn9AjRDK0eIqrPfg69mJe1fU9e2CWGOpWvUyVMu285xCl5/TS1SPbQoCk0JpEkuxIN
JhAKWB1AmN+jhTGI8GgM/CljFl/Zjbv/XUqIUyMZ6myxRqcslSprr4/2TnUgInhQAeaCYeOSlnip
Zx2FtnNuSHAOFqaGk/Ew7mxO6GbSe2TDYBdSjNSUubCbckDvUw2wrHq7MvkX2VTE0sOlFsgc9TfK
jz0rzvzo4SX+6vjQEc+2ERtgiZ+TyrI3lhZOvEsCmmc7bUrhnlNjGO7IuT99cGTe6FSx4ALCN8iE
WF2/PGiauyRg05qymYaBHUFmycN/SjW8RUTVFUVFj3bd57vSI3+so8FuOqt2BqW7nMNLBXc6vsaq
OIPs8MaR02pdhvOsgT4/wB96YBslPAwMUK20RTL4Muc97ZQN5SzS3h6LgvFIhu0HWsjyW7PL46DL
y3zjHdIaVEMaied9SMUNuU4IMQ8YkYv+FLIFF+78a177wQeNO5sgIWNIB3JotQb3rdq2Jn2uMYcd
gdmqxxQiJDJtSnli7+YKpEfjdSjN+N4BrOdN7bnnkBzlW/syQHZdw89dDEELA4CWEcxMnVZKoK+j
jaN5MLPYA+ZvjLdDJd5N47BItRWSZiCvYPpsgo2aYneBmxDtn1PO8ee5VHkxRYIdPfdUcr0uESor
TXa1jrehmuungDzn3oXCbwn/3zzfutBSnHU/5f+FlPWsME37Tq7v5/evjQdXKMl19xE0RXXAYHAg
JcE40sfdR4YLDp7+FwyJHgj8ABlj55ax56OaznL9HuFFbZiI+d0PWWoNhWyEENFMjAeD76CqsAHa
KUmDjDaRJML0EzO6140Z1qKEtBWPPlrvuNmA1RemBMabDQbOdktHpwoT5IOpA7NCRx62HeT/ULgm
i6upP6dgmPjV3BURS3zhqCkl4pTrzwBMMZDqaWX27K1WiOK1sgNXMyB4I6Q5Bg2Kl0XW60zML0tO
ouLR/70rXUx4r+MIFUY8V4IqZNtON3XzKtwTAPy19z51Aj/eOdJaZHBAs+SCgzl0uQzW4PtPi3i7
Mx7tu4RV6VZu+1frgpaXebjDxR3fJAive5qI1qTe6ljN2k0EFnvWr7A+AXDo+YQU06rXaPz/97W1
nAL3BC19pSS12wqDCd2hWFQ+5Vtq1f8+McGzM2H5Gf+MZHsPFR87JTYFV28f31iw0jDTkotvrT7A
IYfCNE9WZ69Nq5xRLubLI3BE04zBdtq8sufAeuCWmxYV2lKf8mp4aSEq3WBkHilf5IAg/xkG0jaH
1LGT7qRyHeyCiIwf/1D3wCzJiNfbdXZfdJyM7U1kA1SfJSt8UvZJxLHA2HsSEIIzWCSY+l5/HNsE
9leZWNTdOEQdgc2srNfySQQdfgamUiQBc8XenKFk4XCYaensjouG6xnfVAHz5c+nNjXJOoHQMoDM
OHdUKDoL3goFwDLdxOZGOOqmRimfM1pPGPzi9kl15xB6sFuAaGKGbQjXuV0rpiSg/PxaKi7+IHms
nhTkZ0CjDJ5CwYvDl6e2TWjD+Q4ttBEBqNZSvdaQrNhxd3ZIhuqnEiVQA+stH65DsblyelbIa8e1
78xziqwNpWTg/0eYMQoGlnUThrYG7LuLtr2t1FmtOaDo3nXkRAODFrvbDxTQyEsIPkBFNxb9/2ww
Of4IGqn0BjXmK5w9cA5G25eaNrPrCBhIt6u3fNQvHeqLMhfntkLVF2Kn2Np9R7joX9fDsBkGoPM/
7O1D8irEb0VErpknvMQOGQkvR368/mFyCY6VApJbdf4QzyTk7GLnHjbeaugBCU7UX9eGE0BzqR6z
BUOEH4iTsr7h0iPLUP4n65YlMB3bS07iGUIz9brGrbtWqvmw5mrH53TieOewdk955b9w34XLnHA+
kEsFXClR5qNtBJ8JKHj1DIjESaBX/0Z/lwwePZU53wyjdN/MSVIQj4WDFi70xbd2/f3QXrJs4dF/
Y932oNXd6u5dNNYYV2BPktLXFvIHZHUT9v2ETWyx16fFseug6KQ9fWWeGx2iF7qNqjzyBra45r0T
uX64AwomjcvYgdwtoD8phT9PdUoQ54ZnrKVMD0tmcmYFM6685jmo7Sr45dIPn6Uqg77L7mPPJ49N
78I0XaL2J49wXoJGKeGvbgbwNe6Bh2AJObplFWtAXTjwYAE4a1Kh1ge1FzvA7uyJO0bR4OVguUNb
tQYU6TRUF9+j06yxF/WE1wfh9duqVjV+gzebwdVJiCBL8OgfUunqTygegurn0A7KPLNaedrnTSlc
sf7pUOzP8JGZvWgRvuHC/zwd/9IUhIzvDqMb2W9dLNWHoXxDQAlAl1mFAdsyLhRqx+WkM2QgLL4A
jKWmojvliAI23Ddu/zA+1TuWvN5oZgHOfTWlpQezkfJTi8rX7+iwwAWZNXSFJEaX3sWJp9ED8kC8
/w5dxmg20f1MixdegyEnVv4NXzLpLhT2nBeJesh+s//ggYKgs2a+pcdxEbYU183LepCxqy/CZceb
i96AbGDvqrXyB1lyl3JALKqYrOJKUorMkPHWm/s2EjSN4/v9xBaQmOLX/cxVhuPBjMnJDioZ1ORe
6XPYnPsx5z9k4Y7bxl6yzNoyUZQyT9MAzZyPDVxzOZx/FiVnoiNN3YJ7CSd8gcwb03BUhsOkpp2k
pbdERXGYi4kFw/vjREFGxBUT1PI4pJXDxSnc0jDt68i6qcrAUxPjCrWznAy0F/H1qZxTh3FB6Dxj
78jXQJskj89O/iV+kJW9yvpXGrwbQtBrciKYgkM6x2zPwGECqpXjvijtd1uzy1oZEUABBkqcO41y
l+mVxmGjat3GyhamcKY5BtxsWAJRxdd5XC6nur3Ul8Lbr6jUZgAy83AvNpDI6HntgEPM7N2o1Ttm
m8UdDYkSrGkTLOIE7ydNmTPddxhLEav6pPJeToBnIUY0BG11DPY7JXSZwg+3C+tLNFwWe1RUr4Eu
9jXHUufx/Hb6kMeEZiMFxQKnRvDMiuQlaBT79ggv4C//voQgFbgksIpmPvygvtKmgz2+pPtktYdQ
k1tdOfw6oBQF+qEEDw/4EoYg1wxclkH/9OCTWstLOpOz6Ky5quYmUdpw2/1n38GTv0KjkwVoU6lB
kAT/UGJTBC3UUKqqsQxCMQ0reFwJ9XWrJMHynTep2ve4aNLFa5nAVAxzIKIA9c+Nd3+Ngl1lBXxz
7ogyZYb72JdCd+sfUEzXr/icbPpPJXvA1wCyIK4MV+TjPfnzsXyuQAhqjebEez+xF7gocFdKKJUF
NXuYEWgMLPXUgHbOjK88W9AuivAMTOH7xweABxz4DbcL5ThpORBepl1GshS18zvZPKHcgtEAp/kr
r3Zp73qEbd71OeivJWbEf2XdyJlPr2BwCFwSQgqR1zkk0cDgtgTx3mDC6vWsryMqm+tAI24VgltY
iDSecqdkMXJqIxpG5LkI4k1dBxQnK9GNdSaLKbvz/GtnXECk4CcEFltkHe72jS5O76lmGagIDAqX
D/DhyUoiGq7bEJoyi26/1V96Fxsy7NO8CzcecAG/HWhhT1PoF7gusteAGTkHEv1bpv2fjPhRpF+C
vVx7xbBUzl/L8DNBSSwCvjn5EoESZlUiXo5tV3HBJ4UsQHKTZFQhTkJnkLJkxCvq16fLl5r92mXc
1ua789Wohsky7XbOUeqsoBBRIjVy4ccS0QWivy/jiMgxZBcTOAyFFADrx1EF8pATYvuezU0xaYS4
nlGPeM1DjZ13XvqxAekIlsiFO8iJJGjp1ACVbmCbt+iLypLKNlOibOzWThC249vSMDCuj1fR4fuP
aCkArB261OXgj/wj8axgW2UN2R0NVlSGZB/9zfwXmWMCo5y+iJ5HunwUObAl7IWrdXJlehzji9tQ
J18D7cokRCCCGc0wKQjpC8e3ciP3HjJFh5y9WcnUjIZDqUBdW6sFonYH6SgqGllYbKoCg8oLOfbT
32/THcCFoakb5Lu4VCYmNPmL1uuwhoNvFR+U0t6OeI6DIpgSqpwWMXCTH+0+byj2v+Xv43gX8H2o
QaYDgSeQjEkvmCdYCWzb2BKrFKuYsRt+9gkJ8jZ8VW3ec0el6808LsZoWCTaMh2aSF98hs/3XUQ1
REHNBG41dWtWwbzJ8GLr79MpAarc6e9fxIGJ5IMMR2yRA/5oWmeESmYfG9efXjXBMoamjnG8+1LT
0NB1VtYLDRA0wrT/q9ZzSVRgB3whJ8SVFuhKGRGhNJgI2x8m+3zCpwuuIPBWMp0LZXHyGvN+jkWg
6xY4ZbDlyITljfYgZdYA57z82hvMn5zyRZLmZeO+BntIivniNElAR3F71NPaXKG8lz7LeE/oTJU3
0WJ1OK6m8ptMq3aiAwCb5oBdwtGyZ/xL00gXi5ftCnX0myElESdfZt5LNygUHYWP83sOHQSD2m3F
9VA5Yo4qxvU9ZDaR7ZMMv+1VS6Jp5/LMQXVF8HNQwhqYOlNoYgkd05SaqCQEBLT6YAHr8jvtG/A+
x/vtFj40yxQmmOlu+gSTebnPBBOCCCEcY+v8HNAGlDv5rvW0w9Ml+W5W7y1Pe9wFiUnvaj2Msj15
3otTFWxK3QSFs+66AAr/BSezCDsrOEGdg3aajAIb2skLwubJDzdtRAP9CexDer4Z7Yyse5UBYxVB
KCA2VMneLNo7YbnGn0TjxazDj/0RfrTyOzui2Am/H23LJ8PRqgNXximm5RCIXQSli1oLd9KZP+rA
YPKoLhJ4bnfczbfiWOQlbXK0Nm1woIFUkItyqXBuCEhqKrvU89tALUfeVhTQ5B4Nq5dqkU0obBfD
6EIEcHyNKwcjbuT0rCRB/ny8ePlu5ozh1yexpeN95BKnmtIE2B1p7HddcMxFjg/m/a52priw4Do0
mVC9TnLhrpUq4ZXIS57N4iwi5WjIPWOuMZRRR8wdMPcA6xitLGVgk4jPWGw/XCfaI1rngBTLdcwb
TnGSX5U/0XiUJHUaez9mstQX+7xnhMy5r4QCqiOE/w0U6khAJlmViWMO6twgr0oA6QHYzNWnlT9a
P5BTbqUB86zFzFrjo2Qks7gpJktlEP6dtq5HNkMOFFlHNVVGL6AtwvklbzZIfCSFJuMz7OjzjgGC
hJ6NIRRefpk1a+gpf5OWcMpb2M6LpfNDzRSr2VN+NEei4ioDtpe0fSRcv21rjP/OTd2FNkOM+XUy
iOrNEHGsS59u6DqWU9GCFOC33M8/v/JygL6/dMHKjm6ZL40k92Fh+8LNuShjt0JBl/vnEE/ossiO
WLA96HcSFXFTX85i53p2N8W+xGfr4fT8xZM8nFZPIOMVCwE6XkcsuBrugPLr7o++Uwq3NmsHLntX
Z1w7yhd1lC7mjPpE9ke0Wu0gZc39VW80h4jgNkHuN+m4aNoukWcgUO9N/G+HlJ6h0phAVU7i/qpy
ahHYWR+4li5kGDtFb6s5KmpSTwKTVWn8+zH/TRPSMbnfMrM7jlfSr/GAb/JmTW8Du7IvZFk2p9Yo
HLtArCM4akwaWfJSPSXfFoZGDmgV72Xi5+k1fwzdTF6FI7jaMmhHvZrZsOgk+2OdQaKqxl2ycDcM
O4f3SDR0SrWZsgV7Ydsg5PquHTlhKowuIEawKqZLcFoaS5J/llCR+EzUB3Bv1O5/nFIPLr49IXZD
EzPRvbO4FGaq7ihwpb+p3RbF6k7DY6UvyrzIwW0zkiQ7VbyuWX8kISy0sHRGxOZGTPoNfmVIYm5/
EqViHaQ9vQMthf3/3oWbaAcsLPWeqsL7+C7PYnjHmzz8bJ059cRBICXP95CtZlaP3X+9mnglLKEG
9laZy7+o/fHAI7RvnJOxkquQ9UIWQ/9IGKInc8zymXHlRuwM4Sd2W6BfGwG5/Zoquk2DduOzzCjE
XLV6mDKdQHgJfFw17t/3HzFQsGjbq2RZ44fEVPNVSFNuoOKU4tCTmUUPkdQrNjPPODDj/sWcFVc9
tR5aexcFe7ky91vhzCR/p2dOSaOb1azXcEvB1MkoDz5IZu6w3bDdm7W7fxRuKyVim5O8LGzd3Dup
f62gHj8nY6JkxlUuKO/f6tedlz2IM3Fk4rcHCXHPc+B7ENL+OtGO1tCD7CpKcvOGoRYnDxkZhrRR
0+nmyEpD0FicVUaL+F2TZX6pOJCSpYq1GNNi+eBwBpcXi1V+scH/emrgJy1U+x8hOzNc9nEEBmrP
hLMmcHsaQav6KMt7MgQrcsXONEn9nO+S15njRHV+5aMj6dOw9LKynij0wVTTRRaHvMB5f0zlvSjL
X8bqEjXhYqDVygaD6q+h9WRD66siPfZXtFMpdpA860o3y1ROmUZNpqB+JMG8RqvgO4hSo5ka8WX1
edkhSgbpAq5HG49+70IKX+2Ied4oz5d35kjZZHrjDaEiLv5MfxjhnEBydw8rRbeI9QddqdKsiIuS
okvIfnOcc4DvhyPuaaFzJsxXS7WXfV6nbxQYrFrJnlhr82tomN3ktg14eCaeFBPSJsgsQ1LA97Xt
wabuS9ItDuZTr77/OXiA51NhU6Ms67D5L4uWv5HjBJzZeaHmGUdbuDKfcg512FKVoaQTtXFBnZ78
4fHxdkoY57suqPaAwKGzaugjvZCcud7IVs3r2QsOn+74pC4A8j/tmsOvvAHSF+arzvdVf+13rxpe
kXHp99c1/AjLiZz0eh8jfmRUMWnphD8miB4Fm42BGgdJz2gN6C41sUbkXB51swzDZKhPjzRSeVSR
+vXL3rDp+zlj1HAhd6FPuhKn5zIH+6eSsWaxs79mH5z26JuFcSoQ+i6uCifTmOeFZVmBNgkchgR/
wMyAdlrQz+1NTJjGti+EtrM/SWQSb6gUYnbTVpHhkkVOl3sbP3/R0F6/JobLNr2QKY7w35CO64JR
18NLh1DyTNmxvAHi7Cgp7Vc/Fm/UmjsP5xKhchBtuRn0P0qcimMT8bsReSQ9E8ZFf6A75yBSd+nb
KzWaf16K5NQBtpPp7kgAD7PBPyM6azR13iCYEssfeZ1Q0mkn9vMPOfRxPGGETxOKn4OLfolTr+sx
YQa1GM2v+hBFPItXZKP5zW1esZ0Kscjp3PTcvYvH+kEaKFVGmFvhRQAunWDnYA6Nz49fz8l3hKTQ
y7/M9jrihtzv5KhAEPXdgAlgrA920yZn0y/rjRP0GZIwJDZbtMbLrIlTdSwRs/+chEao4+ySKeT7
uR9hz103gbgmezS0LS3xsvwdkOihJDINLmAYmh5czAYEj2grrlnfsz5PUHUmUERTnOwxVy+JWvla
M/f63cM4zvkg6QzMZEtafnaf4/aJaULfwm1lHvYGNSxMbCawhpTHmEHro5ttp9n26oOzSQu5HsY/
E/aWfzxI99n4GeLaMwpjc2vU0t7rn1YY4B/OI3t8mqvb+NQqGq+7pB5Ezu0kBtMsizn4c78yeRva
OBGzRik2/NaR+JlO0H3z0Tl35vQ5Jn0fhpOFMZLXw0vkRBxGl0sV3EXTGnS758j/fs8eoUuMIqEA
2q1BMgKcumJHgtBbNsC/+dO4ZtXWaIq+DLlFnEw2Rd4gb3pRPPQF2dHJeO049xSItzNnI2teZCDa
QJm26hh9bgQt4/d+FFO5Z84AFd2CTchynyF0VZEvN0DfYXIs9VrUF/rF2hOjrVbUiere/7FJVJpR
3+qDBwNEhok1+mbNwSNIOSB4uxbHkt+XQS9RfI6bXrpL5M+PQ7w8iSwVQZMo98dZIY4pNUQ78m83
WwYDD4tSxuDOPJ6IQ2WJGyfHIvBUnCD1P7WzY6UTzrjUsgQyaz5g8MwOtluAJBZbS2f8AEmYCsvZ
FSW97qPB9lj5tCYQpHgctOwotbExAY14hTN6OZ4QHDz0apvHLWw6DKZizN5hjZcs56ByNwcmWUGO
lHZ2Idg7eyol7/0zVqv55bIt9smYF/ZbV3bjCloNaYwRIz9eRcLhcSCbukVpgU40jyrsbNi6hAXB
IlU1OarMgOZSl8o3y5nLyzozZ63P7dPTKllxUvsaYnbnhZiw1TYu7gHUgL3nuK5fVaKgFK8lu+Zo
yvX3uyK6c/1+ljR2ZGim9Qx9Z4at4GsKz1JvkNilQVem39HtkZaINNdBsV3DnEBfwFJsRqGTG4tZ
+oyBZzTgSd4T48Vz4OZ+6BIUyrIs7Z3W184bs2me5CB5+9Ih2565Kr30KfUbXzaL59vEurkAtxoI
7M+N+pUsyUMvXqP3FpkKoGchjIQkLsl1rsxsYDwlVSs+PzXLaOgPaX/qIJ/KntE4HViLrGSJ5BFq
Ob+6XzLPfDCuAfJx+2x5wMWXw+0y7z+1+V2YDn3OjP/mpfXXIIKMKvpUEESMKlJKklFL2omU7dVs
++Wtqrx1y3roKBTrdVCVTfeLQS/N+YvXPjRv0sLQnYpoUBp5G+8D8O6APHAtBB98r6UQDcOs+KQH
QGMYgGreg6TGzuze/hoTKoRedFIeeGBHhZOOPO1pGw8ve4y7eKW3E+XmwwgF0rt3kNruWBxEu0u9
/rM2/RrYfgyxFk1G/KRcbuQ2tIF9+YGQYkGbBwGVxj9LaIF7TT5lsKV+KYZjOMvGJl8YJz9HM7nT
9sug6a24eFL/pM42h9JXojIqdMGkprGr/L2hO9CvPG6fJZrNsK704rcB57utsu1yLUaoiCZadTu5
Qo9ZCUWIhXS8srSANerllNoK1uxeaQKtehbjvodOHZBT5IXbN9G8NFs7rqa1cn0cJEogKYc3cEmF
BYWeSlIrN3SyP9etjeR1zvBD/8WLwHuO2jpwqGyAiTtt8OB3R+y7i+mmGGWH5OtyAVbbjOHafFeV
e7+afhuRLvAC7ljs73VuY4v+kCC8M4A+geRed94ryC04/o7EAqmnd1T6tMaLIIw4AW3Yb65tWrwQ
x6WxKWal3w44jQMrKRJjZw67LfrZkS9WeYmfv0MTUmsfYeiV8m1FjE8DVm2xstsolWaKE5cH/Pa+
Dx1KJiRuszvZSZNsKGFtcGCOVbCb1U5zUaI9BSVQBh9ZHGICu+gwLEs1Qbz8QJMmKE/AOJREvIKp
991GNpklxTGaPLmtvx8GB8/l97KB/HIQipogyxdfqDKNNWVt1WFLFaL7WjXHeMXWKjjL1p5kBLws
276PmcSzHD+kuTZtyNC277OU7tOrMwKmQ1EYXQAksYkhmSOUNqJk5ouO22tbuq82EB1FaQXuQ8Xo
y6OiNN/d0BDYU5BLtq4X47GuauwXfYvRr548frUfnMldoxSjwHwW3Uufk+BL31JU3rzioo26PJyk
eyIre06DnP966tKAM9rZGsSCWITzhAH2kB0aXIzMUKNTM8hap2sGmJgtNtD05lWearVMfuWlV2d5
jmWeN/uDI30A922Y4uZByaiN5gIidxKXHn21kX54mTJl4rv4tUFarlBThsVKdjmokMcn0oV0eyWe
ziTVgI+71dYOBqsK5Vd7khEQwGB88LC9enwS+oVW576sjxaBtdusYzBfnRNafhY9SEA1m3ukFqwg
K519qPTN6VHfiKfkaZX+msPcWun8DAwpn49nCtQG8seHkO/Mqy6Bj/+CsuJB24ed9R9rXQpWuiGy
ZNnB9WtT+gc4c+Dvt1Aw4S3DlO9D5CiDmX/sOJPBk+VDahXraNz8cvmlLCaHn4FPfBUkM/ddfaX6
Wq4nx2mChudczSRJuzHHAviYHulYKZCMi8TNCSAnSaINFN2xoqCE+A/aZukH1cmmidN/+eyQtldg
mNFvAN2BMG9k5fLpArm/VAYBWTNfpm+5HyBtrU4EbsyAeXxageXKqMjJOLmv1+tCh89/bOFqR/GJ
GfgTYBwEhGInPhJOpxgM+ufe04C7Pf42n1Pog5Jwy4mU0EJdAeTHg2HlbdyT8f6xY0wC06rPb7x7
EcHFUpuRpDMg9GktHoxJmdtNuNlAlDTNp5WjQFp+os+dbVq6n/NzrOqufdrGJFGkhrie5XIXX5UD
gX20sAMkO6kqu2EHvLd2kUGEGAx0B20DIi8b3HCTFeW5Dnx/DpzwiKNprx+zk79PJ/NT3hp6eHEc
fqR7NysLKA5q81au+G4DpG8vKbRC4weL4Ny2h/199iespGsuWTjBu+cayUd5SAyXeMBhf+zRb0JU
ncR74zUzqc4oZCk+dEjGL5G6wRRkqC2H4any0uJ2UA+011RgQWYPmQzXItfe6F0uwKjvDPXwjzmG
tfE4SDJTghVMr9kIhmW3OdtbpCHAhkxUuHWpP6Yhsd/Ypk4W1mR0nnpERSoAa8DrEXmAe7znVsxR
FAuAfSUjBQwripP/3PkNPUh+5bmI1kNubtSaJo0jz2QlypRNClFssd4aPPVKRu6dW8EfgjyVcE1y
XR/5HG4v7f5K8SDTH2Qtsk8vwzGgt0f2ySMtSKLfeFvmkpjabJZ30Jk+wHSsudrIZiPk1/uhI7zw
+HSzK5NKaRvkzISEZqDPcbOAWI2eOlgvfCY8rhRZaduP0NU8TJM/Qba6f225JQYSbDAN0VYPcduD
DFGkfGnFoVf06IotWoQfKnpz/0MhZDnUg/rmD15l20rdHZ2XggXDZ0++5qtxBU8d2fZxe4C9Udyd
S4i3M+rxglgAkTyzguMxYcP2w2dZmJJN8VxJuKBd73nRCUHpLOX3hg2dFdPcTlYcIWVRzSnLWqH8
OgbEtU96DDRAVkKf32lgi09ZIrXVzof6QBpnVpGsuczm5kAXGC0Ll96sVu1FZn685meFjGa2yq4n
LqZLh7hWRrM+7irv+//nmLW+0jRRis7/6bgwlT8NJG0NNtwT6gXROpGMeIr4B7lH183jF63jZphv
324Z1VxTOtJSP+WAaHdEfe9III/t+IFXuMwuCAlx8Z9HbWOG0FenU5OcPPGHjtoo12vQKmDvQUwn
uLtGi2Z/xBMNtOThkOLXZYNz2tWX+a2/ayCjGeLJr0wJxwXVLwKu5PiNv+P5+HyX8NEJO4jb90pI
Cv+dHf8DsrTMsnDU6SmG68TMuztmZ5fxwd0wgWAX5pae/oeQAodFvSsHRxCuonLLD5ow0FpKoZC3
v3wHX6yrvcT57wMDD7KAxSHL9W+hmMeFS4+nhjZWwUOLtn1Tjghd9VYSMlbn1m21ciAwMkGVtaD3
JxzZyoT0tEYqG0J72fGZoP8kn57OAE1oKNoIy3szRdl/1Y3Ni3VFV/jKdXClBX0Un5idI+EaJPgW
Lu8I1peZjHyONPUHKX0RG6KTBFtvFJrhHqppqTM7HFmXkbM0JW+BYq9j6bbzE64nKuIqrPxIpli/
/xT2/xNfhRsYwyvUzVeQaKypSmgGhZ8X6jFZtkxXJgtCM4g9esiHhbmldlgG8jhIBq/7pdCpU6i+
/vOTYSpKDrh7bWQGRQWKzmzBWCvUz5XcARFEWx2Yx+HeXAb75mDJ/nkxD6gAU11QPYl+n+E7PGJt
9Ihd+thfqajp7vS7E9aJNFbfFIa0K9ArN7JsujdCG8xI/O5Oyv13Ic5iB52nX65Ofm0O7rZV+OBw
A7PWUrlxLMwkt+P0MDIbRqc5pzWFTQXUd/XmWgZhDqUvL8PHhvXqoV7lwD4dqilNtnZybMSylpnA
kuIZrmEIcIUElfWDmOgkrm6KhjiSo2u1cqzs+O7dmZt/2N/7aGEcCUO1MJmi897x386QrvsyrwI0
zh5ZhwN2/Ri3OxEayo35UgS3+Ybxo659ihzu+HQzDdemPIq4sknIUkludVaP2TduV98TKdPSOdie
gG+4TXT1bfm9s8Kcc7/4CDzIS8VT8V8E/KQOQOYj8xLof6kM8XudoQl6PkEbnCC/evj7hrqeYS/9
cssN0W6jBG4nxGtOj6f0Pt9DUTGYo6TcCgOi1KVfRHHwVwn9ntYRoTMX+In29NWN5YyegBPRIY3m
tJ+s5HCa3OhbuIUAD0qEdaFkX5/M50+O4hbTcPrRVNXgM62I0FfCVcTF+inbXaMYtGENyNxf+ffu
PCugRSeWdH5on/y33uUMU5VNOxb/XwQn2bZYeyKJmU46bl0/hAmANZmdG1Lapt21gbfzXvU8cKo0
flM27PeVegbXzgniJ2jUxjGjyzcFb1SVRWbxLKDtd6ULMF5ze/C1Ng7waRAhHaAuRd5EVzy4e96Y
RscXBt1acHP6VoeltB1/lpI+iHcEQJwDToOeHUM6VpAtMfSHEqHh3qNfglSEU+qMHRe8GLuyOj13
y1E3QBd9iNcfdocDfVsaHt3gv0V6jxTWq1DWjR/zdWnrO2dyqRhkjS/pQVh4vKRJFkZYMp6/nsz4
FD9nEXBhLG4xtGrp9jyBN19+gwHGx2Jf1Fp+OEzzVuqO+02wAiwkfdVSU/sZOHjXrr9bclM67CEh
HcbG+Eq/4q/fL5MWiU1ovnFgsM6kOpxksXhIpFPYT8ZogiSjS28NRARiNc2W5AuRwepNjuBTyC1P
Qjs3ecBp+RIuys+l/sIEUiVwTWZ9iEXlpyrhMY+jez5QCcGT0taOt2x6s46HE5fRFM0erh7cROcf
Tpz2UkTXsX+bMdDnni2JvUuftZjsrnaxyCWxZ7aewn1E0VhEN3GJtMPhAoqcm5g4yOeUXXJsw5BM
YhynHS9Ryjw3+NsczfBERuSHWnBUxRc3YXIvUuTQl8tg9d9u8guYZlZyua+UJl0kj2ElxdJAr+mD
UI9xi0m29wv/33XEGOAKPfP+ZBPmN9zp1vj+h/4SI051I6wSkvKIqhD0a0ORaxZI+LnosEg6YOTm
jlac5oWioOtA1IXZEwZ74nu3feomapwPxfAYPBHEvaTYTqAhVWK5lmz/aPIaZpQz8TsQKnh1n4Ci
/qjCnmhHyde9goRiT3cdTjLuBBVkmW117QOXfO+lIlCnD4zo1zMkU9ZfxczweHvcHZ5jg0Digtdd
19OO/c2qToNeY1t3WnR7hPwTkXeuj5PSzppdeDszZWG2nU/iaDnZVtmW+xWtPFkRB5TSld++1O2K
C28RPXkoSITA6IX3Ia3y4ozc5SuKFrQ5DQa6HwgoXXBWnOcNjD4QSQEaWZW3+avLsbgHF4YfZDRx
M+X/dXnsxnDJAZ0YLPuKGnTwwTEosflnkrd09ROEMu2qrdKtd/785Hqkm9rGYTg8LJ8mqNt7cbK2
SkGjZQwS2RpMvxSspXSQlhQTI8OE/uRLwpAr9Bn9Ss7+XzCRHLv7dXTFSiwk42BtfHaN2UreuPdz
5ySrzMh1cjrpidXPLJWZY8b4NVSt4s/hWLqMhAdjg91EM/o/lafXHPoKPk1FYbkNuZvfa5ld466E
taScHm+tkjx67IMCned4rueSLVpfBAax9ZsW5I/GbVMbtKlkSeKcpYgNYeZqY76A0ohM1jh7rFpR
iqkk6+v2D6/lu3TwHw0lq0QM6aKjsmRuakkYP7zTFi++WeuJgAdlYhAfRy8PkH8nwzWR43yxk1YQ
YUZiIK4074pzYN+gA2LBJh1kK47PF06GOnFrxNKSSuioH9PBWmEpY5EgIWkGj2Y0Mp0ZwxdUG/pX
XsbZcrgERP5nt4hN9WehjkwS3VgWzf2eX1Mdndo0yVerE20pTph4NiSHbbuiTCGFbkTJqyHBW5hv
JMGr6JzzyLlu5No4aU2U+YmIrDtQgC1Px4DP/QxMv6OCKNECXlJ2pBttzAY/l9zACb4Pdyrk/eUb
Qo5b9u1+vbeTws8zFLG9JrY0ThN2ovFdUCQskcmFXyLxJuj/I1TNT+abeynauaRaf27YtCv5QFAh
ws6FNCmr1d3RS2Ua8xt1N5UFBZ/P7Gy/8HYoZQ+Bn3ehaUjd8d8WKxxPcDD5sxFSYKFKjIIkCqQ/
vlwYFVzchkUTWNkNqggwb5wUgLGOK+gkpoDVlbTx+tSmiXKn9p9CRT/Da6XtmpPPpsc0grJUV5mL
WvHJGSN2R9rMqk98hBDjDiPem9WlN080KXxeKduqxtcv5HhOG/LHQ5kbOReviTmlrwgNsFuFFXDI
saB9p5zddKv0Y5P+S6J5aLQh7LBKR6jNYs7ZeyH/x1y47HpQQpXb1r7IjwZLxXeluKiXS+MlPQV0
qOicAP/wP3Fauld2px+oWYJpO0CTPfEBGtkFCHcix2b198YEKXLZChQtYJL/imxm+gzgDdUWpMif
msI5AxpxUz/ehaoebVoA0uHGa/XyzwKEfXn74/yZT/4QwGzZbggVIlgjZFtJAd2sM7MjYWXZHj6D
XtLObvdmZwVEQdAHhNTe4u0DK0DueoV2KvZU3H9Js4odhldgWG8ykjOynlkg/KfqBfbh2oPv7G/b
TveKCMFiKDnC+x9hdy1TK+JB2IaxLcaXRMRXcy9JB0Up0zb8bK8dHy/xFhCSGYYeRcbuEa4gZH/V
tS/IPEgEVn+bMrCKxaSzYqoSk2gd9gghiVI6+/lkCR8gbm3xybofsoWKOHLv0dpulO+sI6W2/fSs
dMj/1FimaLlxjapzyT3g2HTlf6f19wgnSDBb1HUgJ3oo40fHuq63lkjUdtgbF6k+hXY3v52O+Yeq
EXFveJZCURzDihSogv5jhXL7yxlPRwX78C7e8fukKBEBtDteOlRNI3UdLV0E9Ja8Qx+CV0VHWq2r
/AsG3WFCPKnmZ3AWlgWqUJa9J5SSE9LBKhsYGL5mWCM69I8yM6N6v1FezttuTs+tfzrye5RXuYCJ
kKQpI2gLwEknhB3TzIXKzIiM+UIdL92NKi3NbLflycZCUfB6H4XAqntqDzTV2Z2zelwB1+dIZJ56
V9GVxAErKtWEKja4JHMw0PNoRnecJZYFb7CH76gw08yJdCJGNFzkUV7UbXPiDhXGRvix2jChbkMV
PZ0pbcmfoXoqtG1eyP5hMj43PSjzZU3MwAI5NDYBKbOySeUXX/Uy4cdiVdDqCU/ExVx1k0aiQVDA
ELE9zW8K5H/sM5aqPR+Esay5VTAyl2MbvtUI2FZqlVblcUDW8IYmA7eFbA8diksMPb9+F/3fW14f
mKta6hynSgL6rmAeHFy8fsvtsW/0QP2wugMMjsY++fDjv0MOG69XyL0t7EZa2aEldwZAp1JSWBqX
ak8+q+bbt7ueM8ffeLWRY6P4z/829mJNQgGK+lPxq4amQcCt4y1w70n3kY0BjIiW5kiYLpU6v6rK
NFARA4PQaDt1tQb1P51pgnAiSiYwfHQ7UUq8ED5Ixc4zvka2/P99nLX8iyXOxXG8PrfuYZ0Hl+Ug
v6ZXB11y+G1yJRjv3r2Ah7tFREEP+Hkrpzx8aPHVirpJMHK/BcI5b002/IwSr2VjxFLWvX18Cs0H
uWBsyBeHGPi13IhucYMI5iNp2AZb57/bzqFMl+qy5Te4VKfaRseAcSd32qMrxsp+PCvQnr2WMrWL
o5+D9WG+/1zsy3/ZjAM4Z41OhcLfOaBzqadw+BJEYqQuNjxOlcBe1X38Xc6503Ilo/TMOq7H7dfJ
P1PGQ3Q1F4CK6T3NxUV1h64t3b4mOVHe+lciqGW8P1Hq0fyVStKjIWxL40Xu35/kfzPcdHAFy/qx
ChflJoeDe70eZFD8HfpqiIlHNqUoA20ZwaR9lz0LUMt4UgSUCQoYnN0i2tSfrtV/DYpODclHj8b8
82RXVbIrwK/wTDQp30oOTTun50d3TemGCMijyM7HCiG0y04nsQ3D7t+UouYIEZuKY03QQ+m+k6r3
qp30zXn4ObLASuCbBuxejdPwDauFjQ5G6eYP6D1FzdyoeLyGNBnymbaaBktzXy2x2m0GdUKGIoKH
OrWhid7/6UWVYymvX6cfb+3PB4KUqZMg+y6G5BCJIgTFFuLsySXcHnv9fC8pRiEXSVdwzkQ4tBJN
8FKk8CzUu80BOt24+YFoSkqqyKB2MApFEV4N6iT96U61gIenjT2r80C4fkW8Osm0BrvW6p3Y0tg5
ujT3QfoRra/Ye6AseFwBcmpslgGBgyau/4MQWZg5/lqqGPdX2zaAVPuFZsuwCMOMQO8cDU5miba5
4Pt4610lLZ8woHje9TstpOYDRQdHhhP2M/T3Tj1kgExh2kyzfdJbV3+m47ndr/BBrHeXSOo5oNFy
yMbj0FLk0l2GVbIXPkZuyrC2it77pS0rBcLBzE2Efvq28FfOWSZzdE2sjE3aLEYSUXdCk64jX9dm
SNMlkOpsYMCPcjCtKQuNhsY3Tl51dI9/NffG68ppkJdDDkTt617Q1DaFjttF+xMSMjtEeDaQpo86
BQ41psGDhNgm0D8GzHwqWCR+Xh0BvE4k0Z7+ZVQ5QLQF9EnGHcj1YQKmPUm4T/Mx5EmkhbJBqpW8
IkR2Suzt4etHDKd1KrkSpzk2mw39rcfqGEIPux4M15NLXkhNQMrLs82fDaIU2kdq2OOTl0QdW5OO
GW6maQqqFEDYe5HqIXBwT76Xp9rnpWNkM27yiugU0L3pFjTJo8zSLutb6TyhKJtUTc0cSHAN3aRm
7d59NsAW0KutUMsbJmJ8byDPubG5Ad7jz6J41bnuHUNf32MKqs8Y1c2Jq/rkoSr/riHF36RsNhTk
QuZTKEaXlbbXHRNqGozWPPDd3ZUp2id41Ron+kzTj2okAwZYb/6qZxXo6CJhSoqMcwIZrWTMXO/B
NHL1JnWU7fIF/HWTuAUuTfV3/lfI/7fKBN66+E+h0+hQjKS98lbz403/jIwi8rgjND8SYVrTNmKW
lk1MlHI6IeFUw4lyLF66Z2mPRbdyxch4Eoouzt89WG/OepSOS6SWCwmodzEM51lMFvpH1aS+e6QE
M5YUNjUHnOYhTy9N/aomFNv+0VGyuQRa/HwCHzI8mNgVLEubvC4KtkMMqB0c4QiD3y9J26/3z9DM
CJprNperApZ0/r//XzAL6JFVYRPzQQdryxCeVGYGcQU4I8UUhTEgitopQBcolvS04MZVONVMpuHf
esL+Z2GYNHkj92DodhOUAMOxqC+zxq3q1T4OEXHygLQHDKcVwpMjaCC0iTsHfpe472L5oOuQ3LhI
iZtjvh3niR01nvFxLhqHpJ6RbZI6inuzLEL2R7MX1eYY4YZXCpk21X0E9UZcRoo2GIzx4oga4JrD
8HRcF7D9QF1KUJHw0ZsDmm22PXz12+sqPjn7RFL4rIE75ktPbtyeBswSVu6lyOjD9HylqTtna6Vk
AEAeQCLwnPznY6cH6fnWftqx3+FBHuJVHIUwJEptMPj0mk11dRs1EpRavJm4+fgs+Syw0ByjtydU
E4q62oTI5TLUbebK1KHZOJeL8DbkctA8gXDCn07W9elLmvh/7GUN70yUMtmLua4Z5R1FveTpdZJh
v5B1IpbN+7tSP3Mh78xUqHFhyQrHCHlZZ/cIevsdW9leTUHeM8aCrbLsCAfa2pJfERywsehgrC5s
a9UpB6KZ9ATFH1r5MsIAiHokTxzg6uTgT8emQ01/RgCr8RaUDvh9rsmYUvQ/u3FGACsEzPsi5Xci
0F9DilkuhrqFIZKOHpQBquvrVwClP63N3P/RVgNCzU/obSqKnYPx55PC/pnGOOsv9Xrg/bMAWiCJ
U3SAUZkDem8Fo5iagbSLjGX9GfvErNyFV5/QcD6l9lGzmDzTqih9iBEJTKibnMylm0wtOPsZJcj7
/eIMltDO4bPEfwI/KLgI4LH3ex6JbJfKGiqiOZNxtVNQAyDq64TqZXYuvL81kM9Yrc29cpPdGTU4
It0Om+EsQM12jQMDInEWzNC9RFKrCV7iraHsRE+uFbaQWhaVX2P5FZ3EFmvthYBeVKArmRpXPxZP
xhH2OMIZma76E+5AGxshqlLuaeghmCujt73U4OOEG9avkMFDyeYLW/k8p3HYo5ChoqD96pneHpMw
UwQrOsDRCQf494tFfGuqZHynzDbDp92jP77PnTsHc632j0Rz/vrsu6M+VuVbuMw9quzMZwoHlbt+
WlDZO5/pGnfyULzER9D6b7HhtQTY8F6vvVwxxNKYyOnSDrXUMnZMVI0EaAzKaPjY0U9epkFW8sqs
CZzF0KltWVhFXJvs9TWyzBg6nrDUkYmiNM0PyYvF8ENntC0a+XNz1UJZcvI3U/DKe7Jt8yfMtwbK
Ow765qwRPObbkcYmARlJ/0urD9tUAOr65psU9pgqt1ni6PU/1EN8a4xLn1KPy821c9FTWIO+a7y1
iXnsncCkekgw+rOw+tqx5qqAyXpUyknod2a4cdAG//ToHeYnInW3riwwgETjYVOtaY6J/Gop7f2o
nxZAxFSbyi6ndxwtU07xR06OuPPv/0QBOxPtTJ/4+5Jrn6M4cP7cEODpnuPO0++6tQQeMmTRfIM8
Sq+dy/K0QV5TRBy1CUQVZmKN8NQwIa0HwoWARSnA+ptB7s9343mZBuKe4e99Z5Fe+2VyyouUkRa/
9VXWNO5NjL/H9LDYxuSMtIIKB7c52aokaw2ji7YcdIqpO5jfMa/HvwByFqaXrIluS8Iu41UUFaGO
4lZxwlFSDAEH3F5zJh9pGO369YlskYYKvVb4OoAKe74zXS0Gmz7p8UUvv0zeL8TjJMzRK2rgo/wh
jd0hWhQUjF0WNdshKyMdkL7cmQyTbuj/nf/jmAmLg10/vXmsz/5r8eYcxpjACvW1CA3JvUT1NzL7
9fSCmkOcEoGF5kk8y90ft8xjFCX6vyWAu2GAVCImcxgl9JaNN99QCmZWrL1G6zrbE73qvnbDYIyf
rLgoklUSrn37gMs4GccifJPJsamzpjC5QqszU1BtIkrmBKN8bK/VI2mjn/JtWaurSI/2ZlBP0sba
35tW7vatHf6OTKGJeqYa55Z4SpUXXWdq64TenJNa6x6EURZ+dWwXttXNnF2FFZmb5Vgyr/xStnGT
uN5q/t6jhzsaSXaXKaFy8eO5yEEzmk27N2VeTV3ZuxkXWd6NwO8mnGFwLKjaQ8oypCSFV9lbF7ua
8edtsz1Tv2WRO9Y3+Sfu6/EQPD0Z0bhQba3+CWMXg5p7FK06X2a+ktJi0vIGyF29cY5pZjQybEhI
pBtI6+TWaMOynOvTrrx30Oa7d887H9f1GeK0c0yKpVxVp7caQt631yMxYHFG4DJV5MorUMJ/ZAuj
AUaNfb8BFfwUki16kcFaXXYeP5vFIN4jbbjmBE01ugRbLgNnO4xudq1S3IvdNRMFnTBoFhQX4I+S
nfGHtT4wl+tArnLqMuUnyeIb0F03jshwsIZ5qkSJQH5Bhgem2bpM+Z2g3S6wkfD7fqXeN7lV/mZj
yJjWHtnzvGNloL5IfNG2eJ4c26YSHkmHdF7nNzjW8IdXvXr76YPyUFRvbXvZOkdTzwYpbiS3vxvT
eFzFiXbWGZ8V+/d09bft2zYNZg91MORWp8KhX+bqbqMzTrOX+ZFStfiseMcFxtvup9lvNeYV0ZKe
kNCWv35x3RifWeIlzqlk1ndPLQLhv9pCq3BiglihqQoLkEYQzjT1UWQfmr+u/T5SuuBF7khQYBuD
qACWUWSTWhHw+D228z9tqywD6acZqtNrKH2lIsZvplK2QWWNIenxehzd8mYyW7EfH229bdywmyAQ
tiPU6xujeVi47CqneNuVRWBSj9bPe9KhSF0qMjZGFgJRw3pXUYDg/0bkyvFkyiqGJmCV4c2wvxDS
jK0a8+78DY3PHTm6NRZkafDO1/jA/BaKtFBjpwVnckOtpvG5jcm00btbBXTV8Q6zqp0+9zSwmEVP
oeuaJDr1jvqALezhbyNdbQs5KS3kBX75K95O5Dh2d/LdrknH6FbyletSF3lxmXPg+SUuo2kk+Ref
BjB0elMCBLXtq289vUbJKb6s3O7iKrgM/fgXqkUw0KgxdZLm6EmatRrQeluTCzaMIy/aBY5NXVqj
QuEC97qJEkgX7NlhQG1fXDHEiUsjHAvP1VvsslPAtgBBiiqcVOyOLWEyHHZqGotvx1j8QTxsuG8p
v/8eXRVffMwAzk6Jvcn6WSzErQG1PDhdnCbwfcVT/oko9lz9swTxueAZUI5/EuCeoamoenYTHOzN
pJItv7EUxSFSJIF5NSCmgWj/KBH+qrYJFxUufWoIqrCw4cTnCLCISuy65Px+Lq7zLMyPncWiBsLi
P9JwTCBV3kXFvQdj50aO7Q8l+Udfs1sLsDPgGIkIe0Sk53S2Mm2EQ2Kzg9jht+vd1EtTB+WlKoja
VMhQWb7Ctqihkx7K3a9/FNTPu0kZsoDNH+/t3JOx3AmoWUeZrE8JdjNdI5ZiUN2j8DzunTyogGM/
Yipr2U55p67lm4tFAq3hYHyxc3i+eE1msfV9W5j+WW14J8crIgsLtowijR6Nm9N+G4/Xz5EMPrFh
Od2ryq+P5uKwzflFQTEBQFMSHe2wdVtevToWhwMYDlxdu5XZFR70gu1NqDomR+Bd7uHdRHSXp37E
yoSEGo3n3Hvp6aMmr89Amg5elOWqhcOxKY8SWcBaaZWVx/gnWbs3oIKYaFalXnyr8pnA0zewJj5S
Yw64m8Ejw6iCrMN0sKrpJ9Ffkm/ejxjQMD4+TPgFY3fEgLwipQYBjRHXpxVhFzxO5IXvxr+XKuKR
yb7ceZNW13pM/3S9v+CfkYCADIE/xAfyxjJzPvRaNmSy4aPWQA2cA7/JlDziBnSasVVbGW9A7YcB
X3AII8yAUglVkwY6WZqzQxnDQ+pBIHoIl2uEulAGO7+/g/Tn/7t+4MhQBoeyonTQjToo+VtW6kdV
N1YwCh7YKvV0hB1uXejnSQdesOHPvpZRkX+jHS+SQs4toS7Bubk5R5F/kQwobTP0SEMCnZePFA4J
8FRT980vT76QKCGghiipesv3uxa7drQrmjWh5VFURPUGzpvJLnoLY5hVfPy2gfK2pGao/J069ny8
X6gTcKbXuSD3bZ2x8G2QM9gUpI0tl6JhTnDCr7ZciP8EXKbkaiodEqlm7pchgD68cc2xiB/kEF5T
9b+xzTcBor9KQtt82dd5KEJEr8m0ZVZPesT4gXCOIxRmG1F7C5Uw5eRzRMeI+uxRCGrJ9k5Fw/uL
QmHTo4VkDHGTl5LVXc3bjSlD5HLlRntjrMPJ+/RVDhh+xAZusyOGfdXYl2toSFUIPRxcQjYoOxOo
ncPxQQSmCNpLH/+NEmg+hu2B1MdnzNb+xbcVoyJe+CFAANpYOF+rJM+oo6ayjK1rMO7wVV1HsaxL
E4bS3pzR8THGI/dawnRmbfd/PtwU9YuCPdEloGvvMQLztSboYRQtMCHeRlvNB42c0p4RccJjC5Am
s/QBwQ06Ek/adxcQ4UfcXX2prZjRu57wh9CLs9v++0aq6/DU2lwCVPkuGml/W7MQxHjGEsVOjLW0
h0+cZlTKOLCw2KzP0aLYhGu6rYtxQeTqeXUzxFT4y1M5mEbpOGZChv1c0+GwOcH8nrdKx3Idfj7l
NCUWCIicFF8Dopd9LFW7J4ioVV6V3h8eru6SCqjJAr5GDokxsX056/5ofYFJ1ijFf9UayWl7o7zd
xQrhqee8sBqcWodhU6SoDbY3kjsaglZd+U+fn+HTHZ+yCcnP7i3A9RoRVpssuFCZtLuw8YtLEZ9B
IZjmC60JXBm5MkollYTD8MLL9TLIJLjgER1jQVlII3f36WfjY2RYwwrtWLHqMbIx4E88w9Cxyvsw
49VSzXF2bxbijM649f10tqW/AsDXNlmnsbDJ/rcwR1uQlflqNONm2EljCsYM7WsW1WOUKJr0tyjK
VlN7LioUN62J0dQbDRZjK6DtYjS2KOyBJxZZJtm459aUtnX4qPFZP0WHvilBKiCi8rYPMFEXvNQ7
W1xrpTKsMsSQAujHzEZWWpjy+4yiXmg/59eZ3Wb1xsj2/knqc/srg4fcSW2vMEEnufTQ3FtTNG00
TZMbqc+E8Mswe37lOZT++1Vx9mFjcxa9+APbb4AV9FszGCB017qVge+Sa3B56VmYuaAgVDY/9fQ6
UJ8wIT4diaC8WHFqCstFPAtlI3m6UdBiuxE9v/eHoRAolR9byb9PMbLVJYNu4vCPRoUDErfJTlhW
dDjYuXb/FXTAb53rlJVC/cvwT4fvCnZOpSLpwnJ79Eum27Xl4EWUYL8fQkopCL5UTmyVdP8n+dCL
TT3iEOvTcLoqntbZ7IhZENU1YW1NSkQaKgXkserJCIMSLhWgAfkjML0HPrOBLikndlq41lVxzM0z
cQmJdOaN/ABLEaalN0XnTXi2d25BtENuE/XyDjIFhTZjsVjBhEpqcLAkoCYrv7zvrpG2GOdXj4qw
A4NGlEHdAqM6rJczjHYwOnerhVgQnBFgKa8bdMY6ed9ix8+AVA9c1OR++5CsWJyMFu1O+iMAljmE
WN5j6VTJqRmMUiMfpemiOhUNTnWoZDzqRrFkWqQv68LIpKfMFhBFeV7GxjNflO1J6QfIpmaTlOx7
tD5INaGgwsLBqJ5LDuvVFd4db9Ra1NSi8WvOnMo2CHsZFhrMT5mCGwofMIaQ+DeBZuWN32qz4/Xb
USjOzT5FG3At8v795dwooxOkxTBLMWoPBVGU9BM7Uwu1NqrkpxGkMOC9V/cRWL0J3EREgcCW3SsO
YNmeo01YX+DyK46OC4GK73+ZrsVqm12PCMM09G0LyAHbHhGAEdmCFq2SJF38HOSy/iYam23q8odN
GCCf4/ZRI6kkiCxmX15Fe4x6/59RQb4SXhJ+PgLyrEY1EFY+Pl5XRDpSTAk6mkyy+Qi8YBPR9wT4
/QYhQuhEsxPMkaHAxdaOSrGP+MucV4ErdHkRDYzCWR5BxLjHathgn/qWT3D5cVLqDZJhFoTmNOnm
UoEgXDipm84UL6NhtFHeaRc1Fir0tpqZALWurLtbY0UC4ROUKX4DToCpMD9GB4oPEuQBB98A/AEo
Fyhcgx4ATxC/doHytfjZgTMcLPMTc8oDRIJPNqHBe/UjvsHDlzQrHogvdqjneoodSvTQKTFCAMya
2CM4hK0gvoCqjk/UC2M+1ELG04CQ/6nE9Nqjjin/OXCOSRTiCdlVQ1OdgFSUX9Bhqtewot3e3JUH
Qh5g5+Js5Zpe8zU/JkII8MLQh0JnuzCFTEWOhJvyq6AIMVO0qU6vfV1pMDlKY3/TiHgyHBv/WA3z
cFk0O9Sf56FB4ZJpkICmK3BHsbUBG8oO6Mk6do/cTgwB1FQEKbBryMP8lLj5Fpy8n6apT4KQ05dO
2D4KgfIAGZ03cwM7CRIF0c9lmxfZ37V26u+prDtK/OPYR2k8h7g+2+8D73zwWgo8A67GAilwoJBd
DHEhnx4vwIIcjo9sTp9m3pJbVdD1KqITtHN7ZykQLKhAOe/ohKjT8LoHC8jWjmEp8P4wGFCb7m9A
DOT0rHmbLHE8qkErNmrKWSdO6vfj4dFzeLfgs/et0n2sZU5EIkfLieJSrCW9eLwHGBwHmh1IfzEP
o+QDY8TN/S6o1DgtcfSBh6UqLZjTnHetuAE4sIm0SlYkgtzBW33ZGzS+T5+eZ44ODQExxS/oBbRd
uI0iBiAm9zS9rtk82F1gUBazYC2B0nCZnZssNKiUcZzTzAb94XDIk2B5440VsA+NYpfSqHHbzuhN
qMxg8Tvbu3l0WktBH1N5nzuqMDjbqksR+fPrHlLudBEkjwB3yyWeb2MjbcedSX1MYMi2/M42sODu
nXSVXElEe2FiJ3xAab/aYaJPW1Ygh7T+sPim3UcUQgJZajqOqoWDoTxAlx0rpso6/zBcL+zA96xu
SZIK55XK/tcUL8cVr+Q0vOksHisMExzjtgB5ufKntIfnrMoemK1FxMM5KKgDiFNThGjsyzpvl5ga
EwnHOTGG1zxvWJ6lsg1YMmLSCx7gIt7wnItYFzbqzIJ3ddRW3cNA9YiDvVGRiW/2IMLUQirOF7c4
lGsv4sCYJ6RNOKXCjpEap18mKLGJmj6wofGmzpnQZDGsk0L+85txbZfhv1EypBExmgMe3fTxXJas
eyXO7CyhWDUAaXIi4/r0VQS0ywgtotK79ErTC66/ApBvsfZ2hARt4Jse/JQGWW9HqoADO3nFkIMf
Uji0khmIeJdN53bgkXIdbo2s/oUizRg4Emy5ozpLoaDH8/C3b+HpeCMMoPEqs2+AgXvF5yvWJYPW
HcxG0jj7fca6/GJmsRpc6qd+Fhi3ZArPgCXyM9LgKtuCRnNAHTGq9X+Ta2VLB9Dnimm6jHwJfplq
nBmNB9s4gmS6tQHAspQhhYoBrPC8yjWpfGJpaptDCwZnTlvjc7FjTKOUEjzWaPFZMORCE3axHUF3
u2KGDdF4oRU1nX3c/OdLk334pemDal07/Pdverlg9tfQMM2ahb7l/j1u//eLjbqvL8QcOjBRersk
uPHY4y+U/37fASt5+qepANa0TWkg2UVUlMYBRs1ZbRkZyU0b/v2qVGOfyxArgtMHOA43y/7pOv2T
eGIcZi9HS4tVPc1hTUW48K/6ScWPLmQbanoDwWRJ+6iUVxFUedcCAzh2Qp7vQrcvDQ4X0GuKppF3
cTsIYc5zZ3EpZyEQwdfVW1S0xOVWq1Pg9zt+xfa4FBzER6engWoThCSV+HD+CYofWu3od6yzushK
8RQrcmK7RkdNciIMcHwxJgdabPxHlphhPXMNE8l+yYyL4SI53fWxBNExs0z+TMieL3yzOuA9X/rU
UvzciYsNBby8A1ZNeO1r/dOekQ1jNTS9zb5uosLg5x14WS/sorVpeBjKCjpxrFcQaHXBy+vRTwpE
Du8Jmz4X095/8NjnZVl80wtosTNkjGoMNzB1O6pRloyPB8FANhY6YaFur43IWIZJ6bBVSQ/NsPdE
0ibkVx+tO2Fe6fbvNl+2Qz+1y920gflv+EXe5Zriuehe8HJ6WDK6VRPh+izrh+NJ3E4ze/7Y6aGR
5CrvKdkHvPReSmspyBJgcYPKXHG5YQcUl1DRgSisU54ibIlNSVNgFu+R03Ty0W+wx7x/QJV9lHXp
yQjR/zvdwhfDppCbeDx+gjPm0WC2+km+3J0g9/XVLAqli/a5LBq0WabYIe5UzBChDokEjSfLj/y1
RJ6fZxtYnllKIu+ge6r6Q8LEGarSlfgmMtNIg6LdRItGFK5VuQsymoMvcChCug7Ysgl294jJzn17
8DpgRazv+GtTVqhmAWVFnmhbkAy69/K77kQybw2aSWErgrwjG0FFcRjEloSAQp+vYJGBDXIaxp+c
1vYBBIWPx5DqTB6ciLVFJ7FmF0JqPoTXeaCq3ij7vqR14fQTV+5qj+u0gdjH071itQUbvyIY0Twa
IU7z1WCDL3NKFNiNuOYs4fRfAtQS4SyG1LEhpPPqWlMIXIZ9jTgCA5mFRVcMrKCSiCLqmXPg5AZI
HJNNcqggH1Spd6i7LGRVhAh6Twn7o36FREt/Qm7gGUH91YACz9npcvCRpPFZdrlyTlZKfV9hndwh
Fan6C/1+2sDBG2gPjAUU3aGuvRfuerY1a/ppLA5lVB1IlX+qMOkkv32qKq/4FgwWNQv4esuc4hBa
TrMc88jEUb2bYSq/E0u4kLm+4/cXckZi4YRAQYDrIyZpxQpqZKN1MacR5dm3AHYJjxIrDbHdtip9
wC26I8iCap+dyLfbHKQu02PyfZ2dRrSpPe8sLVZyOuIXbSOHPSg1J9T4cCzS52kM/oBpwdYFPGD9
0xEbsGrESDrbwmJ6PGsr6tXNV6chsqBgmUJ2tMGaG9G9hKegdJZ26zBmDTYq2fIMkGirsdBtkKj9
uEq1TVbcItjKJVRVoxcQVLMsPLELIUwKX0O8kIHwSEKnLTVZaOqdG988RRnvvGtOLOEcYwmwNJMq
Jx8bOztE4TjL5gmq54JQEsMqvbjBNW5MoNeKRvKJcuQdrBPw92GsFGcivWSm7V81otbggmhJb2mi
uKAdr56R5cBUTrhzGgIPbb0t8YSSy+HNKUOucwv1Saeo/usV+pClJvx1FqxIEGpqOccERnxWbhEW
xUAS9PEB67Akax2eiwHvaYTV1fO1rZs/mxXDK+NVNObXllrz3V1nzHz9JE9nUDCcdGgyBsDgVwh4
PaFlogKiOO1FU+5eEJ/xKBWyufyxfX9OQO4KsPYibsiDrkeXXW3YrwKxUKIQoGXbMPJQeOQhYjne
Kj5dN66+RryJPWomKkA3cHicZ9NxfEo/SqczSJ1/JfS7spKsowkHDjtDPjUrBwSMa1a+RWk+hiuf
gTlnDjbClLjAUsjttFP1NKwh7bcWVUALsbzkqgJxBxCopb9K/xXF7pmRANwIac6C0Qty+bdVB9Ln
1anzrjxOfumKrV8ZqOXLRutW8yCpmDtkrUOyHW6AopxDHKEqqnHurN6mgQN7VoaqYv/822hPM9bH
xNVvZ09Rvhy5ain8+Rf/TU4V4Ek5JYHDQq0Xu07YgZkn2rCfVpBofVHg5gUJrIEGweK4t7r6L+Tn
aRcmMIL1DyzAYgUKzSo8kGfi1HGuwAumt1kcmtpDL/EidHsRiq8UIRyqeoHyNXBTA+QEwXCNvE5O
lutJA6I8tfJrEx7SoZ+hE9JhkRi0MGLFgbc3OENs4IKtw5OvbOl/VLUYGlubjBoeyWKac8pHiKc2
6Oqhxy+LsdTiYVq2PHBbyz1RzrRwYutlV5K9qwWHTZ9+JS+FweQqriyaGtrm7iFG1EaV+qNudDu1
HpfrNYxgRdYmmafXg+K8ltYt39wRhfpITiUerSnA0w/2Ab+niOtgjA/AuPjN7NwX49QyIbqN+ZqJ
7Oh5oh9XnPoMlMAdGRy4tjJI7MjKk9m2HcAb01fO6yhodv08MMwdm1sOO3wx34HaxCDogMpvW8GG
KMw/1thu1uveTPWB+q5tLsKTUMVxMZo4YBNX3P8ayRpikxpPOOUc17NCPWGr+5Tum9nL9Y+COuNr
y/A3vHf2tAmZ3imb57ew4Y64tGfkyeA2Un8/yhoSMDn7KIlqKazCAk80cgGNUu0k33nIJGlFp/WD
n8tqn0A4dTX1/2qc/myOcbYZMBSH8vg6K3firEGBN8HqZdkT2Omfelh6AxA6/ixV2eaPfLLEXe6y
nRXwy0sSe6In6UKyBxjA7Rch2Ec00MEFlk+58h77iCvaMOmBsiPrYmm1t1itGIQpda04Exo0uG+X
hiOtCbYEOX7x9WjwKJm9VGjtTqslkkY5Y0/tTzkPRlCGxFv7urXYhkDz1TcjI3YH/3d388fIpqBB
ejBHrkGtAKOMOjZpIHqIswbv0L6GtUPhmqYZvhbAGqBOQIFhfjwTf9rKGDL98axHFY/4vwktlQii
VCJ/8h9+q0zD2KSnHKCgEXfgQVVOkUgGkB9jbnaTWfXok93aHq9Fnft+YAUmCqvhnmUqLiHBKBhU
hSTUY59x3+E1Oy9ZuFuzG7trm62uqJIkrJ+/VTL5cAJ/zDgWaz0lo5gxoPTPf42VvtTtq1nFtDa2
iQXdjrk/y4pQelql/Poi3FwB+8XaeFE2mBdDwJM4B3SJ7bX9QVmXDkCde4r8PNmE1EJywsl5BbEl
wUeI6TQQ9Ez0EZ6n0tjm12uggRaqgzw2z3HCh+chJ7d/ThXsRYNwA5e7qeYjI6VbA1e/jvsT/pGP
dOWxAwlN8jwMIWA4Hcm54JsAExhyRPmW7uLa0T3AwSDriV4S+3Ik0su3OB+XPxPLhfuRZq7ZA0NA
/P7QPOFGshXrWK3+TySS0g8SStl09rASST1aF2VG9nFr75Y/m0KoQEkLsk30FqIq25AAziT+74k1
ThGOaOKZdsWknDQId62tqkSPcIO2lCJDBGKkwyvqc7691JuI8kHPv9qbneWmT64GF/sLy0XpOBls
dcvheQeIB+5pGcCrcgpbEMC3pm6ltFHcVABjMtbaKqeiE/ReJLRq9YkPOqBbF89XzrfrdqjiKm4A
8UY7evqLS7jkivOKdwB9Q5UOgIIsoI1Jgl7d4uef4NIYCrv7P4Eq5BAlak3AEP+14n2hMDh3PkVO
yn06v9gNjlbOxYxJHWjwAtBGV+XXWVq5m+pywIkw7GtVU6LNaZ6tZDrKPC8i2mdIrjDtqI8FOrx8
PpHSVy36o06mUhfxfjyR93dmgFKzZpHSkIpqq6/ztK63+WDEv6Pf9eOkVOhTGj2xswSWxMerTd2c
epnE0VnsB9K4tKpKJEyrx0ZTszgyAL9sM0A6OKipzjw9IoPNJuxF/2/M64otC+RtcvjwHtFc42+u
zDm5vqGqeNHfl4ZdgCuNIjAkas2ukZs4e6WaR9JjTzdoa+kyRP7rVCPzOgnjWSrLZWxjK5MuEE7o
w8r7i2iPZfdM9YgpxN/B5L3GRt/QxMfsmDYjostC4cuATpFsjYCnZRko/hslaFdv9D8/5cI1qssF
4jElzFKrQ1rS2xhkWCduUeyCSlW0dGk7YcErOnKhIEf8PsQGSeFJeeTG+H4npNLYt07wa9iD3Agy
68AsC74927BtV3jH9gHToSALVHjwi2iKbU4Ct5F4TXrFSnavG5F5NYWeQRvR3KpSbhY7Q028v89Z
c0h9dJ9LeEKQT8KQaJFrjqi9ylN0jLsu7Gif7YXps1h0WjGXB0UygduDCr0arj4zP1b9RuTaIwDc
okHxe2cQ19M3XC3fAFn4OcLyg72s4S/82Nfmd58Pi9vhbq+ScGtQcPIwmCYciceBzbUkHS76Zzpr
DO93r7N+Gp4uqxLFXUevPlkHuALs8OOHOurMqP90lBT2ct2pX5zyjuaPiR5UQQ1L87oZgr1BUHoM
ab/Y/bb5u7GufmsWZTg0KAGDBD12RT3e/HPY3A5Y/YpTYXcikzspNoO/8lLSb+Ud3ak+9LvYMd9A
gpeVqYLgZyHanMitst7uboTQHCd9WUmyG7d3A6IwIPwb+KGhD8GuJe/SqZRQQMtaMR6Cy4pljCay
03GgE02vkIoXRsHTFIObA9cVDURgsYfArfRIOC7L6ci08akLTKGwFwPnRMlAqXn/o+U5HFRsxr8G
uIMZOnmQkJqrI0T3xkZwc5tKtZOcLWMXm0Lj+yWfcstC402M00gMcyS6BIqKjM72Z6cht8uA5vaj
LiJSFpCafXGjhuSfBPmyxWHl+sPtvk/HrqWlSVrZ2jc5VuJNDvYJm/6/Kh4ePgVaCQNgwK65LKye
hAhN2IfwgCXMdMtBaaoUurO4GP5MQg3eUJokBc2Q0TYU1k/cfd2G++wtgaZFAZ0scVzthuJnYOFr
ZNhViDPqI/d8gSecVNa61InTHlNVudyBoJpjekttUewTmXj9dnDkflygW56GUaJRHh9ry9apHY/K
0Lpeoq9jg9hkCUHWigPC8Id8hA03WuVCBagvsV7WCh/6CeVM0OVGnDliR/BR8TYBNJNSF/UkNwqn
PDKum2nhyrZ8UJjx9pPn1FHywqoS8KW50mpU7CZryJaGUMarrxtMAOOBjyAWf23VALmJYP/EbVa6
01aJKtCaA6MSzqytixICjsr13ZJYY3iaDPHLy11Mek08qWz2pusvDCW4/qwTaokWy6oijg6RdC0A
DlmgfFULa5J6OIw2QYRLwZSvzQb31IRLT6HwJlP5Ob5p/WV1zj6/qp61wDyYwuIOMNJiL0CLxdsz
N27vlepTthIYMPi2Uk9Gp8yIhXUgNJQAoLU++Cvc5uQkZFPb0cTBU6xKCifZ1UAmV8VQ/KfgsHHX
mRCVNjPJghVta4mZWO9Hakvi1WjVWoGlfhjppp+x0aRg9H/F8tVDaIyGgF8d3rCRBFIeVl+Vc/rW
ARR1bHJA/ZtwST6H2zNy8pOYBY3SUqkOT1tK9mWCZJRKsBJ9vLGOPiqnhc4EIcq8AxF52CGOk7gE
AxIhLen1Kiu9H4K0LyspcF0KRikTN1vZrtD1BBz8QiNg36D1uEAoApiYxhgOcOjK6oemnvonsYjV
nNJnZsvoY7WoAqMYK2do+/Z80+FWdKgVzTHh73a/YaspWXdb36WR6xv4iD+vo7nZrZWtDLBxOqP9
8n57ZcnbM+/Zyt7f4p3Stm0rcdecwgrI1yG9cRy70BCJh5RxqvGld7gRHa754cbYKSbUOdQkexOR
fD5FEyOm64BT+mFuR2GvuaOWC2KBWktEw3J3uWsfU1DhtwrVVFEnNf3xzr3Z47neVQIUwDhJHtYM
9az1LIkXmQf4P0WLEOD9GV/Bt+LDwXF1Vfuc8yKh7CKHQGRY8lZ6C062ItyGasuoVK6cVu6RFz0u
aKRHKlPnbAlrhea5ujpH7aOWaWtPLQl7JUrLoywf95mk9hTK1nylu5TQQMPsT4T3gxyenCF3zfIB
bIjfQA2Qla32NoHaU5nhDlUoYe+OP+ANOtDdcVM3zPRMF4vwxY7nXIjHd75O8mDxubCa99E7kdlP
cXfqzHu0gWSA3KOtOFH4156HJKzarNZAidP7Zv717tm4mtdnmULL4qeDbOzQbMvboKnpPSamISv2
Dp+LfypMQrJPAfwHRzZas6PLSxWtxkScwE9s5AJ5wFXF86N+LWWztzC/n6612X2T40PXHsNIIeZb
3NbDTmPd4xCHSk0Ay8rXey52bBpdAVKiHbTnIJoHjN5iJ5KQOAe6J4pZtQ7VuISobzCSh09ipJXi
5VMhUYy+Q0U6oc04sYjAQXHZwjjo9w778ix2kfA4PjYhvtV8O0JNPps3buOgQdnPbF37HcV9kOzG
MmNNiIX4i5OpHE6XqxsFBeFOMTB9DH80AmAeK7/EFl6p8HI9/M8NEhuJvpmV4ZzQWNTjHk2xRN3S
dgm2vKnqzDtWz+FfgRz/hgVaOUqj/CAuRa3KqVzude5T66jNGO+b07RWQh45gDfgfl9ubGnuHZzA
kcv8NXs9P+oP61Pm/fxjU6AQU1t8VGHYKGq84OtPzNSsRWsg1MlZi1f9QJl63FMii2sN3bgCIZ9A
u6vAuOjTqmX7hDMor7S2fQa0EFJEeumfcZxzJYAiiUrsizBcl68TSDavLR0UUVZO/2JLFaAX4Irp
x5owLTlEMDR8TYUOX1jYbSoRZH8xuzIESvuG1MstvLYHOlV04HyHsxJyCnCgcUfus35Xhb2vw7ds
yzT66PhlUNdzlDDpO4sr6CWwjuB9zsQAw4nXCd3jqD7ryxrSOM1m8eycTOKu844843Q/uSIeYhdM
QGtMjIJn13JHn01TZnwdR59Iat5CpuOKucITtWmSOHQsMGObzjV6OrVe5YDLgEHyA0zxEY5MjjSg
D19NeyZ+bQefkOjBewNoOgIi+g92BicsaGetkxEwrsrDm+lqdHjWeTEjqLMommRCpT4MMOTj1bOw
S2kttJz/aQ5OOMTFSGugCoVVmNaQgwZA1k+IugTWdY57MR5siTczmxl77oy2KG7GVsh2LgEGL8/V
JU1g2LhkxHOOZAdvykF6qTjuEKfq16eOoQpJpnZD7VEmX415I7C/JwcP0nC3yPBeAa6AIVYrMiIQ
IryaqYE95/0ASRwoBG5mAMRJoMaMHU8AA+7MWpXuY06wlEtXvhLylRmGjPGw3qp2mfwYv3kcVFrI
Ll/pKAA7ixuADEqDc86K3YOf3cAjO2VxLLfnrxZNwLNmkLOo1iweu+i4shl3roR/LI8lNQDm00fC
Uj+LTJ1E4VbggCFrfc3bNe2cTR9eW1po5pY072JOnyRx2NY6iF8QG0AMChL/3ft2NexdCLnU+mFw
hv6JRVc3gVUXgM93ln8+Ds48fdxXniwaH3F/SCp7pnPDT7cF5aVgUnbgZgOZ3hMfDqQMrVLxCoJ2
tf5NAEPn68Dq9zkb9NMW0E4AqU0U7xacJvomHbTF1e/0t6FqI1DnMNyvUn7AD9gqc8TIFtasNHnj
1tgLwhVBu7Qk4HzqCkwTdx/lls0TWy2JR8xJgfUiqNquzO3UigLROp1oTF8UMBWZE+/u1QjPuGh2
MNXV+SkYWuHQDi2XcBXBRIeziljIa7W8YoJO2XeftsKB5jl930pd91ZxWdswtwajzJ85XNss6Nbw
jGyYwKUcn91wS08rRw5vBddVzuKUqG3qMAfqbXSKz3HQW7QXPFr2XJ/9TTEbJ7VLKmENtOGGNM5l
+oaoanj0CAYscFYzfJGqcMP2sqCevb+8hIib9nZYNiKhJU5Ql65hTLpXd5ze1+v22p5i4L07TTyA
jQ9UyS6+NJBe0WLSM77OYrypsPcQTRmArNpaFchkWehU/TnwRQVVtR26sNn9LrMQq5jdAQwM0VTp
dbSwrjFYwxS0/LrTl47jxwl0itw2rhzHVMA7UZrF5/rAIEk2gtwstDbC2lTUJJif7fT2Px9P7ZAB
Jfg5FG/KxSJymWAXpeLKYjJeY7So7OsPS1ZkpKBAdVaDFCb6OpY1S8mt+VrYtzYhTJe5TrmsJU85
/qci7df3yq6k7qGPfJlCU5MUiDYrSwKR0OXD7JmSifOkNb14E4HB3ZIWhh1HV/pAPQRsEJFId1zM
lM0zsIXLysrIzD+oGg0ShErU56W0RzjVotqeQPOdUlTyPyB2gEQUgvFgpYF+smYQBaFKTS3HLLqp
njcWuA2SobXsP1ZjfJ3z+e6dadaO1YgqJ3XlI3jTl0bQUC+yifhB73EHb9ydGW1j7+4QSb3IdoVz
OyLWOYu9cJGgmCzGns4+0xM5PWk8rrmRc8d0e6+03wZLqFQXAojAqK7kitJVSe2vWe3bapL+/3Q5
zhP8+WjVNBv8pFBVkbI9+4EhTTXkoVzwts6gnjgv7xOMVL3YTRuneV6xa7mn4B+/j6Qh2lBfgU00
nCq1obhDD28nTyhS3U5Mrea9fRXb1OcXsE9SLcEQZHgrJr+yshn0aqLkP6QX+4VDTe97Wf4lGLjP
CkbACV6DF0kdcbE00uZrUKuIAysEtMGjlhshJEcwsc60ix6ryikpODmYXjsHnBAYY68GmAeYnB6U
HNNmdl1yIPHKaYw2/6hmOUL6MjwALgCc0hilstXQ/7wBPPw4ogBlFJVtdTOoDDFRTKOngxGYnChc
k/4zIyLwAZxRBwtqMbDpkE/qUpqbB/oGyD93dshBwzSoQaFF3SCYGOTMAzxZvodZ1FOEQRr59Woc
BPgOp0+Ye9ZFUeZXQoaBA/YFpIIIRPLdRsWxb5MFui9N9c5d/F1TIlcQcjfYpJZpnBCs5g6SkpfZ
5SFBwgHLOGyC25C4H0esrH4Udjngts2G9kdEBkbKS3s0W0pnztHxCYxZccTlZxROz4l9w7aRGYZX
B2bFixI4PUbkTzeovutdZNMgRFeqEZvX+K+qS9rQrW17/8Us5HxmhzJn7IFiAeqLC79kT2Sc8D9e
U1GOajjHsRsXUyLujEkwjI3CvfgIOQKCRx0x1vc0xtEEkdzoKX+L0vREtEfZB2ISKxRKAe3Y9myc
1G506qFoMZ/8w9syAYqDklyvYXkd7g0ruY27tqtrZPyOx5sVn6jzXkr4I/eNXCj0er4UOUZqHCV9
X+T558RALLR3I65l5U5akaykZkmlBDaEluH1hCXretTdbUthSzDkuR2OAdIu0zOWAGxcAhi588zh
o57g3rLXKnSmZORhC4jvPF5fNHiE1YWuYINk+Q2EP9cUAt9diEuQu7vW71ILuroCe/qYta0VMEfw
yTO21WKO2phX8cJlbFiRjouJiXAm8+Y50+EsX4diV/HvidmFjC5KvsbM7U/n4D8yTX8udcwODFku
A+eTX9W1qCuNPI8VkTK1hijdnVFopgIaphwApDqEZ1o56fW/vYC8tG3Ytm4Jf9vn8Hx74Fbc0ile
Z6ynexGJT99ii2vjVktJTUqUxoMDOunHE1kAmh++S/jpnCfbSUtqZxiojiut4M8zyHUHE9Y3pbU7
xD4iwQGPSkKdLR8MZzMutuJTv0gNBjOl3/sqFyhAIx7MjKHswSCXfHQ6NOVkIrKgqYgMIwTWpFcv
UAHFsXr/maFGh0Ek1SdF66aJl57ad58FMFr4ZkhVYFzj3/Bw7qf+mOpDUw3iUHa07dKy2nY9Xs6z
scRteUpp0bavek5qxt4QEPqg3DfdSktJeppAIR+Py77q3eSmSRl7YKr6HjScldF8QHKwX0FNHaWv
mbY0dggRIpc768ICupIKNPR7169ml36qO7GIkxFGGWYJgThIpbG5tDUKtYt7DQzWuKhsMwKt1O1k
qA3GIDvFkGnCWcAPwcdPndZT/m3z7haU0AisqZsjewgJQRbgWF70YfjnLedHFP3TJ6h86xiMdYGh
Evf8MHyVP6wCGKZaV7MuHEctP3F4HaFW2vyxiRLXw0i38JdaNg5dd7bMOJkQN64rCAxGRBTYD2t3
a12w0/D99Fap9+lI1ILEVLpwryUS3rZLTF9vjNq2pmBNE8gJpvEX+iwKHQXvTgn5rVmoARPAtA0m
gLT4iGgaWL1bwSk2tD5J+dPvGagsgo/MSob7ggqnX4yE7P3/ZtGL59EhBfoQx5BPJzx3ha50IxQo
WiX8T9CLmvdhxvF1A4Dk5jsWYbv+kJ1RiPrqEIY1K9BX/kUejAvHYfPcCAevKEX0su+1m6AXCgvf
GC1w0y8Q83bdAEyJpKzeSc9r2z9YCJcNPufdOxGkGw8MRF5xua5NeoM+gL1S6wpE5zLm1lGy/9Od
ZXKAfdhCckMPAYEN+nywBaGfj7NV7sj5DFvxTXPOcn8cuYC4BmwdTumbkCxO2s5X7ReQ4LkGFE06
0aE/KYfCGAlRU0WmmfTbGoJy9EzczJuWQxRXEL3MHvQcJVIqKhMBgu//ZHLQnDS0SrI017XnnBgD
fr5ZrzE5EKEk8vbGKJL6X4frO5sn0NUC5dJ5XQRoWVK0zEEuiinImdlnPl139B4WtfFUv5WM+ENl
7nO1lq6hr4Dkndrt5dTqjaAnLmFdZxJBvwCoUBs6iOvb0baHs6Vj8A7jms4wsYZPgmBjB4m32y78
oY6iLg97gLul+HvApJfkkOMz9uWsx59qlaZ9xgefILY1aT/DstR3JVLgZpgBE+bpXrDPlcOPjscN
mye0S0e2a3gisTO+xJwfwpuq1lGKcByvzwSuYXOeJv6h7upf3fdK6Fx10VJ9fpn58MJb/W2h1sEX
FpdeaFtnkQTKl7U3003uJZIueZOMksYButspnS9ZBajGjFiHGcMGtAEgMJk5zsa3ZZ003gmvRYMn
JGJZ36qhM9MgmOmBHhvJillkiYKazfXuA3vDOhlWZ6Jz0eUIA/Od1EKysiWtsK4raSbTBoHPxqLQ
G6jSyNjmu7V1hwrl+ER0R494f9OwxLvSa5YzgsM/JW9fScOGER1q5sKmARUC2YR9ujagVuQqva9K
NblQLZJetLjza0YUuj9oyzbs2SzUJHWUW7z1R/dxB5/JXDuKU0HwH1tw+aeiHYDxePgqgi2d/lKp
I0uWPqLMUkCoCeuXUCjHvNbgG5b25idPMK7SONJqAWz8RVNWWnHfw+z0VhyhVbjZY8ypog6DYzWg
tMd9nCRdfkIKbBla9PXreHCmnPqiWS0EW0K6PJbDv64jINcmfhjOnxFzT6Q0Bdri5lJhOWIVT95n
yKGMy2Vn4h/83dEcYaL2QUqzRIPWC03uum0s59IK+omLuJ9N2ELbLI/lntzsZ3X+36BtaLfczAve
zREntI4mADNM15XVnb9aFRr4Xstaz9A+dpzPLZwbM0ZB5Hm3rftRQ3iqCuMAr/hJbBqvavdpR2cH
UOSQizyh/JJQowwoWaINCOSCBHHMwXksemog7RM1iMW6MJ+mMpVRzYxveBKsn7q2KsV3979aNJpM
DAWR2574uBtX/iZj3IgE5YX7A25mLlXjUMy1s3/Os4aPDh/hwWf0K/AOpL/amftpPp4krGySuqS0
GQTl/IQ2cwC9Ft+B3b/pV63ERZqPB76DwHipOdt8o6tclwxcwNGrvbaglOQTN+bjFW7Yd1eAh1L8
fxT/z7fOzJ+BbVZV/Uw8kit0EGDgFsvigDDRk7r1AzQshGDSppiho9P/sctYGA3cD2dFEx1K2POs
sDZdAIB6fuHGDqtJyyeXFhNikYgqPJxyR64wuMLEg90mz75XeKg5QbHz6KeO8j845pf7VF4Prx8a
npB/xtCXPq1VjdjRj56furTXj/rmRFDsFnYWDoSw3N6ZRrHz6MBiCY9XToBvbPr0EP4jJ7FPZ+j+
ttdr0fMgzFghFnbrZ9qJRloDuL1QduLKNm7ZWG6HztYut5o70kXKsJ1sYOB0Q4JrzUUJbFlIzAUw
dSZkEk36A6dg+g7fjum6DLjH9UFqj8RzjIJ2RjhG/ufqL661jtWYjyU7meLrM2uibSvlXcc71p5F
oR/VcKShkAyM4J5KF6gVALcUQ/vwkgwnTn0xu9tyQLLgEKotqnNSHoxH7tb0oiGgfMA7eRqgalE1
QppdlSdoS+oIHorpGqDZB6QW1IvxwtT5fhaJ6RNU1KRWR6Uh/UuR9Dby/QO2C+JFiUF0eZWvoPeg
3c/+Pymgu/94ySr+JNtvjUvyBIJN3TY+uetGu1OQWLdsO9WyA3PvYljHUNsA05aZHTy78MLQ/Pud
uhf4ibZVi/R4i/GxiuwEm5duKAivBGhf0ZIPTs9QchNceZf72owVEOswbKkkjL3d+CuAckihNv6f
UEmC6vlc7c3HIFxVP0cDSPBVTGl2YvU3csBJoK9PXXy4qPqueVHtnnYiq3GeuN75hrI3HbEZI/+e
OiJ1/KbmauSpQXgpKeuAqH+Ru7PeyhPOXfL9iCIvwVMk5Rrp07KqYMDpuI/kXI21H+9yDAdx32E2
DS1916GLkH8s5O1hdie5u8e8P48DL7sb3xH2SuKWbVACA2jhCZMEyOVWCXwlRMxSG86t0r+f3Uqu
JIZxJwdKyycKEZ3x4b3slD9vHDMd7r7B7ZGoWiSXeGsilEzWfNh4qCXkjeZUMtw1cW0IudpGIK1U
UxQAjwNSKRheopJ5sYYnKQ7mHshdWob4i/z3qDVjU2Z0ShUvUUJuE7KJNkE4d2DaCz1DM8eFr4Yj
EvPfCzm0XLBEtUp66jmGpeM/dPCaGplexGldhQn/aZ9lSL4k0hwceHgYPp0C+0DbluRSGT8Hnl2a
5ADgap7bR55JfJJLN0kMz+K5C/ZeULSUcWW9ZzSH+u2hLq06j5Bb/9gyHRx/5ez0VkOKEJlNVmQp
t+neSi0Ej3R9uxY0t9B8Qbp8dMrrqyDJ9B9kk/6GNmnRulrla1WkSN7es5IIALMK8J2W5nDmCl2Q
RZYL7B8Hu17FmMGUHKMi3tQ9sWYoHXrQD40AfmjBpIsxnYt4UmhLgbIIFYHoVvb64tT87Xiogg1K
boUQToLfZVB29JzwFZnlKNMzVqSdWwdzPSxlOVmK1qQsz8WUjYEV80sB4HRXOeYvu1CbdAbjoooR
8bqcWDn194yz3hPsOh++uCOC5/0Q+wzMzg72AG3L9DjR1wYG2/b8FUUkosLrgBXwdEPOKPoB74GJ
VPs1J8cUxHIp7JgGDwhxEBSa0nuZ1fT9OqDJ1HeM700RyQcigzzv4aKnJmimtAlUT5Zg8lkG29pE
l+wx7OTYWA/9SdKwG/1P/R6gfz9H4N6OYlbNSw9eWsJvt4ARrfeDDjxEkCZ91nIsfLV05yTahh6b
yzkW98hJeOaV4mAHW49niiyQJjEIiCEn6Qpdw2m54wF0PdZ1BHssgrHJnt/3bCn0oq8bMnvxahVg
QObkrfFPSuUkdW8+UT7Wa0sJSVEpfcm1rXy+Jyr56ANipf0gR9+f6A6LKdlY5iZEtrV9tlfcJeEY
CgIFfQLWCODbveycPWkbiZetd7djB2mhKVsSX4f3JloNFON4XJ2Vjt54QQ4ccAUJuPTK6ZLA74TG
JD2sUS79HpUVmb7TzQ9LzjzyoVVSsYlJbD6W70R+8izOZILu803U3JYyLNlmG57Crz1XenwpthPy
HujtcA0oR41t1s1/uetFnFZm3pLu4+P2cYApTJAVHzIggBFfjBxishfFeisG41QcDPWfzqv1xPDp
fp+L7lUymNo9Z4LB1QjFJU2fCabP7vgbZpwgmfOsIvUd61NEcQJ8xSAJzdTkQ0Ym38jXliIbgYRQ
G2sLKnNvZvS4IQ5BPhLeD90ZV9cSfzZC5gaHCeJQEhdnh/nSjpk1ifO3o9UO/OsJyNkUOPbuj+L6
3DRVGGX5274cEjyixX2cZ6Af7qhSu74l83RQNhswKiygTC3lY823IApFtJg/K1SnnPHNzVozK6xD
u8F18Cy1JkkrWkIdic9FXyhqjUeGYoJVuMt5Pmn10fiN3mBmbup3wjRoBqe8MrIXt0XS+y9H9uf6
j/znxRpxb2tWTCvtvb5RuBadc1BTQ6CQh2Z4OGue3FYQztNZjI03UWy9ysHmisMsnmDo9GcIorrE
uKt9AkbiE2dxEgKBLE8hDcfhhNGzgS6Wg4BDvUKT45ZX5/dv6hrCKboxPWmd4d9XiVOOyMHcVTD7
9cs37YD02IcuqzMYiZAZUg6FIcnE/9eb6Ug8PmoMQRqcjP8hARarGNZPA3DkAFwWNsVu/aYdurib
AbcUG3RNjzS9Ck3Y+630GhojstPjHSKYCJjqDAf1QrPrY0ZNfyOn9v0t0ypBNXa+LZETG60dnSPq
c2CRiX6fTK1J3B9Q3WvLUUhzInREeTushfLEZ0eGRgG7r0aDHJBqOTZliu8kM/meZblYAbcogIWa
LfE8U5gwq1Es/OgMDmDQ5CDTJtgSkAJDTor+NBm8WQnjupc4EHQeRLvKAHO2bGsOnOBo58Vb3WXO
OAzyIA4IWrRSFTOhPk1gtSjKTGDMamDMcwKtRkNusDu+2OmHMpnirdd2RRzXlKFEejL0g5LfTPb7
YipmYz7s+uv8fKD+EqGmPgQQ4Ew7lk0q9mNIaFZY7NAXgqJVZqPhr7y9bew28mjBWN18r8E+gXtn
HCtT1WHHFXzIinwMS3totC4hPw1T6WS33j1k5nMbvFRXRRuLl67w/+5mq+co8Jcyjg56NW8q0JRz
LGtOsTGuIq6o3k1ZVBrCVKeN+yA1xt5gPfgN97HtYnCETkpktz9HZZulsc2xpv+ltfWsGN/DJfm1
4NTUAvVxZcb71smg+tuA6+NqwuMHlv55TopBiiyYHbQszKcU4gr8Ok8mRuIMSY9tnuE99NLKDtxi
Lucjz2+Fa40os9uRmiWLSJvO1qlpBYh+qlWnTFEujxlW0n6uzxSe3kAt8ePybUm6R3UDIK5LHZ5W
1xAMBhDsodqwmVV9wG7508g9kX7U0fJLnbr9kgXYuf7PWOKfg7kCUyTYn4dZZagnIcBp1GDetoRp
sQBQelm/Do4l05uJfMZhup+/TRP7eGAKKJOz9OU6S6JJSyPWUUSVAHc/+pb2P3ammaJfDAmDS1AR
uCvWzlFAnBhg8aF4aH3mNxTwpk0QgGKp5T8WfnHfUCiKwnnxhqb0Fulexa+k1ViyUqvvVRFj4i41
9hk/TR0JLe3Z671v5sSZXw34o4mKl91fRU5Zq8w4RVeaW43fpdO/4ieGQq9//yWbDrtI/ZiLGBXH
cTXUC1XWWBh8krkFxRsAJfmuVZcfsEe7jyHi75Vgrl6po4krTXC3SLuiTBUeIH5GF2qdnZyDVZsJ
rfsDzkHtsxhobhw988LwH9gtTAipkMAybdrJPqkYx/VuFd2uXqUX7/PrlDAVuIMSSMaRk9eU4UQz
Y/RUzZRF58cvmUtvFVvAWuPKpxmNNSOuf59a+h/ooKIulPfO09x0miDgJRv9U4Fp0gwxEr6bvD3H
yPIICZKzMd2efF+uSIDeZb5TuONw+RPsyIzoHriM64mo4vc/cOAfnjPPlNieopYgo6AnrZb2T92U
GdNNYyXcYuD80IMB3h0mR63+hACNm9bdOJhto6KI/1lyhttHT844PiW6k00TMj9x+5YhyA0LhEsu
JZUPQOpY81FhZ4pv7ztRRa6QJsDlON8KpkUO5azMI83NWMeV1vaQcbiIYhObyurXjdekfUkc5Wfx
SbmzV3l7KJ8FfyqXwAuzRUg/C1ggMWEMWgSILIWENrxIcMiR3acYmdH5aMtWE2qskfmGk/NUoK21
vyegsKsNRJpHtm5N1AZl8UbGWA9PkHA+XVAaTDcQIbWbQ0jh/nybpZCohLcmAMFxvrR2Pua/AO8S
9mVhvUde/WkxnyR2AC8hNn4UZIL42oYBpdfahqAMQtl1aJ9kpQAXa7/gAhizsOD0TkHJcVBmW6vO
JE13PoOv2F7aNwb67Z850qRrBibUoase9AgAV9ARw/16cGAJXPp5ATUBR8ZyFMbn79gkm755PvVA
9JmnGtEy2Yln9Ii7Q15OPcuhJGzVqQIH5WkoCF73xlc4mVYGXSxFtodHV3Ex+rsYNB98f4DuPHFy
w3Kk/oL9l2w94DkUKr6e9yh+fUC7V63mUhD96fWvPZQO5h6NseDTez9N3f69+2GfA4rOjFU5SkcS
onun4SO005TgVcusyFy2JbW+y7ew2AV52XpLDm3AWR1Eq1qlqoPjvLA15rYnNUWzJrIl3CWxDtwd
RcNNX9ZT8cYI4vvkw9TlxXsODwPvFJhlR+c6cMnoGYLyflBZSrChKcpbzvrTbWD1xtId07ZrwLQ/
ftFYYMC8dF1Tl/XWCmbE7GX92qkQWcGV8gmCQBi/YQJKpK08dD4GfOGw68ZNfZ/nXJRCXeuGB/yg
DknBPICPasmUPdz4nL+yaTBxLfWfSxJ9n1bMOhfkoRLehfzELmFbgTbm8M6g6v3ANwhpCUEZsKOf
RxRR3LoBkWKP+FiEjxBRvq8jDlfi5jUPXl4hO9r856JSr95wzd9UuGdCNtT0zjRlziRttuNd0/pB
Hxk/rw693wN/vChTFPQe7Y0PKeMTiboC8ihgZGwRr/qDlVUaXtsoVrZ6v+QXLHuR/Si+FaFxlDEY
otiK4ZOAxIxHa9kd9ayug2KI5HQVf0M5jQBkhXmGsbni23lavpUBK+uoiWw6BGPBwjdsjvw7lejr
PSP98buRnXMT+KskNtiw2PsHKiZ1UKr6vezxhqkbkXz9rkMkt6gXVVF0j4S4SogsRWbqEE718oy3
IQLYsEtsNxooFygirpq1WHL6neZwvWm9csio5/ylZwE05hJMJJVIDKPsE38c7eEeGKk6DnE8GS52
lzcA7okY6uxIAG2i+miQ9M4Uhlpna5RabH+EZQE++1EkvnmYOBhSVEeNJL6Ew1jQXBgF4GRdxUTb
J3OVQOIXhhmM2jMvcS4q+NjvjFvwENaqhPaMDvz1UZj7PC30mSscJoK+mluuJDVDIBUzp6xDnhsU
58fahhKABjeFZREImRX60gsbBR5x0KafUTReHCquuOO45M5VL8Yy/MwsUu8GAC64+ZJYumqlnKSr
rQojc89F07668DioPBPdWXWULCuXkKWN3KANWCbfKFIUU1uOGbOAM4k5Ohr+5tSAhoJxJSPw/jps
o8Zd/YpvTDoQpuhstqOgQffxaIPcUWDhbHmrJv7SoyqNbDxAnBniW1a+09jhAgBGhYo8MTnSvjoN
8fAjaIGGxBWM3imbSyMmqngDWUHAb2E63hNmbayIi4ibunaHV5W6Nn7vCmoO2/1rC7n1XHFJ5iXS
atSFf/VAWCv0dI939hSWur2wHbfy78W7ldpoW43ZoCB4QkiJJynCewkzILGDww7nPhpzPJOFrEjF
fTv9SpEd6dyimFBX0xPWdEZFSnSs7VKw3LiYkjNodlYXlq1EFWYzD/XlhFXKaaYLGlLTKpekMpha
IebhC+5mXfFyZxz64XjAnmk/oPsSs1G/D5NEYqhTYheSLReSz5eShsvxBsLjo0a5owJ6fxXUiJIy
3XKdAcQYHnTcWP+3++MJAKrrFnYvIqnNjHDslKpibTXcWmdR7QGPxhD8YR7ZdXZd+xUIDh2T6eFT
vdgQb2ipXFUEkEvCg8aROoR7V34/td/fkw+NXfsvxZtXntI1PHlp4Uj4GxMWAIyBY+ciOHDFWAZo
c1MZGs2Vy/s/5jnj+bDbToVhm4Ppu/PWOs/cqrUaesvh8M+nT6AX7KOIjOzTeaIWyRFI7v+LWzoW
4Y7c+zW2XWj5GDNBB/r6NVxf7H3y19hGdtFAc5+j+fz7qraEq+te/xyIIrbnrUHMEFGjGWCJ80JC
YzVA9O+ry15F3ooObiN1+k6xLcGczUD6Wxz9tikgCA6U5H/T/G/cYOsEsRmQRpGanLnG+85+iGwd
lfDSmYdG7hsoPN3Zb1HnVkODbFN+QBPT+wmosHM+sEsHxqsECTPsvbgL4DgFGxoQjo8REckvl88q
+c3caYJoNfQqeC9lNMNMbTEtGjS/bYWI4vRz7ShT7hO4kpsIA34OPCk5cqgwqS+H+XgLkLH+F888
cbJYLygNVEgieTRaPhXfVDQPG90DXjis3t0xHnxCNX+uN0SpNBRnthu6vQt9/HHyamyV9C796ygX
Dl3eovClhn8a0yzarFpB1gPVhtklXkuaU0aZW1UVpfV4PbhwcKQKzWOmmhHEC5REflij9oaZELBL
Yl3BdXAm2lcfqdpP3g5RmFbAPZsTIzN+Uoh6Q9eS2/jx07BviVqa6HXucTU0jqyEXgxnJScb+P7N
g8Pwuei6xL9FGSn66rzJ5sF+6AAMR3/IFPu4fPSaKmBHAq3Dn3tiklz8senqwBnltnVJX8H9+zq+
PzPfDZ3+skObM/f8nmkcvaSD6UHw+0GwPn/Wl77IJ5yF2aV6WTWRiXJ19VlKBtmnG/pBRhvRaW21
h+SSIC6RaeYA8wPtTJUTDD3N9CjVga9FE+CoHyzduI8tmRdaPv977mtOh7q8hnig20bo9YF+kKu7
PsDsJG1M+uVFHJKyJ2m4ykZc70BSsV+kcbgAHHkydpuqKJZ3uHf2xkSw2Dq78D81F9aL0O9ZenTs
elFdrOqrkXZnVQne2d/WHlENcirFJ7V3dQxUilX6RJ5B9FwvDZM9LA5VboC/Pwks/bE97jBSBMEp
S1exFlWVEexkv4XJxkHyn+dXb0Cvih1ctFWiflk50k5/MpKtmI4tnN8cszzEANuvG6oGhuhqYVqB
Jaqyq5dljELxHNKhxllPA1JukEEytae2FaOkewG5HOkfsDHk7CrTVvmLM0n2mpkaTiWSFPwlzSIV
4XzV7oTaqWUScOTucfx1pBBJjtmOQmYAWyjFD3YZ3coVjA9sI6J+1fNAAOXsiSdNM9Ld/W3R42oA
2ObHkPq8KEsjhfYxIq8+U1MPQrG4CfrRHnFEiYb622bKbC7Tc8jRkp42a0w1dmCfiX2KIUWtQ7Hz
m2sOw+L6CT1k34cIWgjeD9w5KQP/ev411PNYhBelKmyL3yHOVVwrRZ2aCbAhTygOYi3YYF0im7I9
IQJqvCXqleZBvC0X/P5IMMYF48TX2/4dask8fuWUSJpQejbgYIJrtL5nI1kDLJsbNWhfNzSXQTVR
ELrC+q64D52MBh0+3Mx3Besj8ah1YWaN7BoqLpQwZCo0LkqAc5tAEuXOrBRKSA8OLgxJUv/SZ0uo
WCz2LMmwLce6Hg6CdDbUuJY/oIUKC9+pEusuD3nfLup0Wvd8aN+lVogV/rED1DXzJEFDIPAnBHoc
8mRNQZDhXahX6qxZJMFypFlvff4h5i5Wl+tfswe8DBVId6YZ3jc25JxCX+Ah0DxGn4Y/hYqdcm9C
hRZYrQmvr662unz9btkJQQrzD7uJ4ORq6/0YSFI3VQdS2L4DRj6KCt20PVx265PHmw35D4XNYuri
/asTusT2oN/LvsbaCqlUfyzJNwLF1/gwDYLpBmrbn5WJXoJfjeRDB0xVANP0yxHmJF6sZ//yHpUP
ej6dQTdgt8MLgCcIArLk36Dx19Fiq0HAUvQWyaGyezMxp3WUhrDaDHfKakzP8Ic7CK/0F5D15s0h
v7Qj5a6pp0QH95dPfs2DtSVjaQkuIonOyL6S7lIqQ5ixEw8kdiCBZ0+gCKJBzZxfNitdVbnBupU3
cnhS9g09OGPX2PAXiUX7QD1CL/uqeN0ksFJYOL+V+1SJQnra/ubkvNhHI4PGxITBiZdIRZNhCQoY
/7F9YNBHT9115pFJdpPlO50jzFtwWspwDVo08YCFUadIjpw6EvhTCK9C2Fxlk/SNCQyISdH4DIQ8
lemTtUKACJCos6rGNNFmW/mAAPxxl51Lseg0D52sFJSfhIH99GDDhXqfS/TnjA17uQ/n/kos3bj6
OurLw1DXS6j2jgtH1N64qTRVA8oXL/zlHfIofxnIJCb/6qGX9u1iNpEvjPQ3Rse3Fkh9V/EkM1xp
wDINMliERZky9MHrJ8o24mQcbN8G5tRYK9j8pIhB0to1jp2GLHA0zhHBHZbLVqR3Z1WQ0EYY6Tcy
Kvnlismu17mxl+v/QML1B/HnL+2E0T1EtSzp/eKimUmM2hmYcd+wx2oKXu8cMj9ry6+cmbpA/U89
4GKW+P8X5Olz86utXk9fF5TksGcV8LR2iaPfitPDTgomWq+d9Mz70LFRSwQSzT4ZD/PAkOzOVKWs
KooUQvo7wYIAyXZ1fcf+pwRxIo60fpq0CWSNOfou8L8hOWxtpCoV7oVu5U0kUxgsNZlPdlgl113e
WDhMcqaFd1bRWE71Wx5U55VmCTaKGW9oQHp5v09lwL1QfpSkiQwHhLCjh2z9bOC9XIvyGPv/hAPZ
yaZugw/j2D/URvTxtsBLzASXRwv/SQ/7fD5KvUZA33lCf2ypxUKIy1sl9oXIaInpp41sEBqwNgqe
co5etKc47Yk5xq3yKdKYfYz6kfDvkr1CsT7r86BAJ85aeKyFDOD/fUiuRKwM/gBh8yhfo1HbvyXr
rbmjRCHxn1ZPTuhw3LrUClStqmJSQaaLhedr69aNY1VXEqS53aM2iVf+/rRF5nIef7fFgH49PE9J
TO3phtX4E7LJzBkr70lYOU8kxMD6bI/Tikvt0bd4mxp0cfEQa1humF4DxSq+ahHF9M8+Vg/1u5Sa
DnJ9NolMP+BZHQxhkeVIWTISLBCAGi8SqWHowkpD8Oico0wm6OfwnaeB2h1EOwAf/iweWi4b+qxd
QrAham3l4+3b96zlgwxx1TM2ft81j6f0PJF37kS6sK5Irl81A+SpuQn/I0KlCNGq2rN6NCgnPmFr
xBt+w4ZxveTi2oGHDr2Ub5lij7gHSNqoYxIANXKgks/2EnrZJV2A/cNfW6Pblm7fZSlrdmuCk94d
B533vnrmaI4LVLrTKVJM1EOiVHrsY1mQ0+LKOUNpuFS9+60sPcAnfOeTf2uT+RMcYHrmO+3CbR86
KzCjK6hkZU6hV4UpBeH2Zsr8jHbxl4LR+iN6BZL0f/GbEhg5xdAUN2cuevblg1VDvC9tFKbE4ZXi
kTg1fQrru9BcMNLF7ct7SHn+hFxKt0yyBszCbQP82g+lhr/DOsiwzG4V/PHJqE+5DGA9zm0uhyxf
qWBsFHQcMF5dYrMMQrhom/2nyIjOACvQckjvp8Om2wiNzeSx4Y3ae12XA7hDqH37cVyCG0QvnNGr
abgtw/QQntIYzyz7CWMyGLfKrLcXspZ7XAUi8JHi135nlExWBCB8Le/wGgB/Ti74NORfI0vgvpwq
ALbS00P28ZDVVyZMmv+WfHZ61FI3ZhGj2o8rim2tQzfFvaqEOaRtKILrFlLwFzfTWUFtmQD7YFFK
/82z/LQ2dkLVByYFX8XDZZ3sSwLqQRVRp7rEkop6MZ/vnnnay07oJ6HVTskTHSNsHwA0q3xGoUMQ
0LQIgPOPcOikU8RlLbCaBo2U/q4NOCApfBDkL8B7gfeWVg627jMWlhoFvNYoVHMhLcGqQldbaYod
EbcDEakc9OR8bhe/6UrDsFM8oyoHDai6fGbyRMU/qqq6/QYToEQPS1r1RgWXBMZayUTSTEqOelwU
Q6U7aYTEG2japbDWTYZEftXz+PDmS0TmliNOGNDuUu3RDHl6fOWyJB0o4pnk3RDVjfVc/v82Q5tC
ecBWI6QnwzJfI/jXVxeqNwA/sROZomARk6FMfgbHBG4TsHhz5pkUuROLNmplO9JPaSPNBT/DdC2K
tdyRzrSJH8ApY5Ze71Tnlr5/DuWWbXNYPjtbkUrZnMw7Oorx1cgJjBYd7ErzhDYrTEUspdAY6xfD
UKfaBOlCw9KIPId89YZC0LAoAXrGa74sXdcR/0ETyhBrLiQWsV7MVLX6WOsQeBSdUgbFUE1ZUZtO
Hcl07b78DpSu1sbxfqhYRG+ieOQ+H4GOSWQhVqfkPcPlMKLRBSW0UzYmKRBhiUjgkeVQUOwOLWo2
hL6BydgJNG+wziPvfqfhX1B+YZgKZQBmuFU3FsqeCzWl7lyjxZMNT9EdO055DoiNTdc9FRu9v//k
8bHDncJSNnDLmgxiIu+dGlBSoqaPvBRVLghnbdjAID0LC0qwL6Bs6D92YoaaGWV6bC84+njnh6kh
ZYT5OSTv6BYPsSC9MH6PxS9zveckYpemR4ydr+JGKWScbQ0WaigqKxKrqaR9AeTBC9yQS5jevpHC
HdnxApXXGQjMfmlFCn9nQGhvbEEP3HjQXS6G9LWU7A8gxoH9bEvqZ//kARDTLpFUDXvpmSnmrH1L
y2IUxRq6ZflMS2AvhqHFFpuT5RKmLOAVgv9vk4Yo7RrsEGpiObUxbs8CJl4mrF8zBVCfnDAzhSX5
MGpXLZbrxD7LQoOEPIm7pSzWdMGWaYUc66pxEAtafFnfC2fmY0nTaogz+EtCqvo2oYLVyZ6G+sem
uGaXXLdZaT+FHDwuIjDVt6lHlEeSrul4w+1eenBIZxzvjmaXgo9pYRavwlvIljtIEWJh4VWHXa8+
657vVQgrKlM45kNumXKpe4e8HtVwtWrMHmLUWvQq34gck+8hdLZwACpB8V3/RWN8Gw4iWtx27Lq+
XpqYHPjZZI1Q1vU9E1J01qLXgPcqXFXWXQItKJ3UlckAE3SMpP7tvt9J9o3KfhmDneHqyDUmk9bn
dEfqQL28mBP6BuhTWWrbH4Gwa6PZPT/rPE1XB/nLHWppr81ibzCGpG73B8Cpnw9RV/kWpvxILuW6
0CrL9R3vbK0WAlnJNTSkp1y+hbmEKp867itiSIa7Gtmn5w8rg2OFTbWcqJ9lk4vnoVDjdvqOyKDW
0JvMQDHHxYuO41tQ0+jrFL4tUVFld8yj6DMSBd1Bg3zKIiyLkZ69h2RI78DMC2L1oJFeSllCEyrC
UqBBwgbYgCtxAgPH2CnQTqMruVstAA0g2F8i880QROWRVHO+eBX/EYigCTM9xOnBceIteEfBWKiF
v3MFuSN34eOBdszr2EqcNJK3CjzYHg0H+TJjjEQrjLTKva79jEa62lGRMrjXSiWu6eneXL9sFB+4
a5nZlE1EGojY6/s8ka087IN5ix8tv15f2kJXgMUHr65nIx2lqzJNLkA+J8U0Uik1LK9ZTIxQypwC
7CcDydV4EYfClmy8tDJUu567d/6N1azB560r9jatp0z7AX2isgyTTnyVhy1PXOPO/yNsL8tBWWra
TPtOx81Uz8h64tSU4yVNbDmFND6V0/nE7+k208+4ZF/JzjzQFXHgrnF8+arlTc0FJFTLm4a1/jWc
28bMxPVx3AvqgoyEPtMafhN6JGPaJqNSemIECyGptZ7K3+Qxunq4eUzoRVert7khhfd4dYVpLVBY
hN4Tao2relUgZD4ibEgEPHXxGYKmC4tgBh3J/g0WEeOCPqzaD6wGQ3XyFfysvjGDrvIpJlebbP+4
Pd+klv01lPaMCNEf0UsBbJqvdUHEkUJlDqvdxqVBXEr7CfjYBFSuHbTYfPNcvxATn5zTo48AZcY8
DkLIs0yYvrszCciWkKlfPV2nTiJ4+tDuykepH4LvfOYJpgQ+N06X8ps1EwtW1mRVAwc5oUqxCQwY
Ev61inyIX3y5dSTVr+RY0NF1Dxx1MOuVTz1IYTAQ7uKEUJQRF1zuDiwmtO3ylCLDZyxqvEB8+PyU
FzrNgy3b+RFfo9dTT1cE1268P+DTBgACzJDwydXTyydaGjkaT2heCH/yvg/tu5FP81sMpnu3gFtx
zdt2X63/jw2CpbACUGqRpjMdkdVO17dwm+EC8/S1uK1Nr79obvl8Iq61pOxWSR2258qm42hpjg3s
XVMsEIOOIq9C0CiImY36DBRuveex1ZtggUqPSzz7t8PT03ryFbcOIHqfNT6wUCIh9Mhhpu6B457B
N/pGO/S2NahpRsSAv9b9frKu7D2sDpY0oro+/wzzRx6ahSKxWO3StilmLYy+m7fwMI8n2mhupdOb
L9SkFJ/s5h30PHrmXb+GasoZToUT5Gdbp5oHP+lA8BS4vYFIQW3w5ZjVJ3uScz5ywUyUSQEt/+MK
2nJQgMSDnsHRktwIF37xpTLUhYcR6HTLAbmtfa16BPq2OUGiApqVzEOBzm3+KmWeoVv5NJA+T2gg
2sdPNpzypv2qbCaFRSaXIVIPvhhFtxGFsKA/sOZ9FOZNzPqrSAjz1/JatWjjZWJrZb0hq1BZqZKo
JjsiLV5uHe3AtbBsgF4llLX5Js6RI60ErAUZ+KB5WJh4YpYSim4bRwbYDUb3aLQ/cr9jSfZrW5sm
hHXWVQAaYVjoy8T0rBqgkhsOPCnQxvOhQvLDNul0SlFKXD5EzG8GWQ0ZVn3+YPap7ebbWP2jB3nE
t4TaHi69Hi8vVwLGrclNuaQ5JVqbOtTepbI8cugmCOvcXbpOEbi2uBAZp3eCVfclmkLZ5sBiGGw+
zgzEEU8my7LwuhsWXMbSwiQDMl7XVKICpdQs1DBkPJR5nQhq8nvOwygoOHBuLHtasRhZwjKkS9o8
oLI5Hje4NchUKsfkd3I4pr5Zq3MDg6g7rsEhehLKE7ycVIlFeb0y8diPnRQ9moRqGChbdY8UO9GO
r/nHMw8paREWV+03llaQsb4ITswsrM2dOXyaXK+vG1fKRgdJxiHSzPTGPWX9CJlDU2CWd7YE7ZLZ
k4umtG0mF7UATsyS3SMsw++Ca/Nmw5gARH0HxTqiP7gcF1W6+rqqmEGsvHdWFzrJ6+9PDmdDnfqx
iRfUouB31q8vZ4ZYMsPdx0iU68joVX2rBPURM87Lqvfn56QECjBTuznDNEd+JrT1R+BNSnjRfTqw
2OJB5gkE1b0Dw2nQsJCI42cbzL8RwJ3flz7a7ShzaWLP/IqNfVJPQ1T4/gBnJj3/iGkNiUV6SCRu
zgfwzsdTe1WR/XhmjKQj2KadmsoHQV9JJj3CkZQfsnJV8FtVF2wtDAVO6/0BTKRwjuOG2/IYnWXJ
S1yAzlJzzjs+83CfhgJM6MdFBubfT8PAAkOkfo7r4MTKbqHXl31O323puugCLG9oU1ObtKjnRnfi
6L9qmRDQptI/AzhZBUeZWqDsY9AKL4xGVhkWTx7pgi6MwjvmwcHyWs5wv5jsWAe2R9O8Rcp38LK5
3g7OK0Zjt0exopOsSNa1bHDRYGUpTC5PLQWXRaLcBPmKDpEvp6MuahVpRvQr6jJOX4khrd49LiYD
YDC0lBU3H5Ffq0BsTot9uLz8VlsAFTO0iXBUZ/gxz8lvk9Itm22Ea852MvIzo9CVE6+qRfYALmNE
+R9KShWGT9rvPme+DtDZFplLS4Ch2V4miPCwswHBOETkSTi3R01KtF16m21T+mBJZ+/9r6DgU6OY
cCZr61wcH4fz40/OpJHGopdyKS3wo93nXZD8Yva9btkKNGFJHcuV8VIj57CrA113ZIX9u5VTz0ad
beNGzF1nqaYDCuKeFZzUrZwS8h4r6x92y4vpWHOBtSMlxNdSv+IlxlZFtDLUHqr8aIQGWVtib0U4
Z6vb6WJLs55nZ3zSwXlEjjd/0wXUJPKStTeVvNrfTcl9UKlz8Qc4u7YmY+kBXsIZ5eOryN1kYvxb
bSXyfh7y2AG9K1S97S+m1Hs+VQ+0W9p+zfMofpGVv2jjku4HsxqBGDhlPcizid8Um+SGnPUFK7uW
gk3IkPLfTlDYfPe+oefJX7eipadRsvWW/IZjkrkyVa2WHFz5/pwX/vrInDv1eh61lQIs3HQ9Gy5Y
0MSAJ5fyP/ftRO+w3AxZG4lS5ePc3iYCBLTZowvP6sqVoyHxoQx8y77hKpLAsqIINOR4Wxz14gd/
aHOrWrzugiRqDvlMfn+vmqBvgcd2URxmnRh4DK3V19HQqMIr1nswCsmQeT54g+6zivemysEprmoQ
YgwCXysI2+uIG91r9PmFEVnpbpF7F0ESDylAPMM3R+dbwjQo7fmKgBeyiSp52vA6Ri8kozA7tx3I
cgxOeWOlzvk7xsfWnIZXrTTGmYvou0PdmHWhOEEFWw8LxQy7sFGyCAjxTX06BLReR93+Yw+wxDWb
IjL5t0BKhmzzfRdWrnCF4oJNTOsTtQwkllsgz/Gct3WUr9HRM1mQCUsCzHx3/f0yqF05J8pOLqhA
bEANa6T0ugo6v4o7FU/GTTvJ+I2Jhan+De/KgX10mz0Ldofad5hInncwvHQ2qYLfUXXBXockKKmC
RrcnrS3Am+Lc7qBEr2DMLHuw05AOhoWzKBiZCyZrpBm9+Yts5viQNe1EGeAphXbMvRYO9trEpz9y
8hzq2P9/Vpd3oth5SzdzMpJVQ7BMcS1OdB5kOH3z8MoVoRlA10CO+XdPNl+nnkcNcpUclA+aolEE
RaqsynnO6orx8ur9VaZ+pM4nQXtBoLyomEpFxW+T6H754pPnwksx98I8n/Ugr8yNenmhpXvDFhyh
D3JRkLFP0UST0EkiiwUFaeOOJxHeq/uQ2waJY0mgVqlRJ4kNv7LMbcUjKrcRR/rC5aw8OBAbZ3WL
RYj+y6FbJBujJ7Rm9Y0UQb8BBbsjE6zPe4uNRNUrjmLSx9xs+Y1lp0KtPbsbQkZ7c3jyvpO0BMyu
MlkjfvVN1qwn3jY+LinPUUyOHCFi7RYagqJVEGV92GcAnSThOiMdLQ5Ov3puM7qGd5Lpvqi2Ldla
0Ecx9goJHcFfOc9g/8uFSNoYL0n6JnpPLycbHL6IUaZLmN0K6SfDvOuu+5IuHXYQxGaNQR5sH8/k
ojbGBGceYfTYVFkIYcYoUvzyioTYRtlLUzXv9xzQqAA/mMLfrV3vqHsLBooUWTxEi6dGMF/7Rso6
EQ1jvnzZ7zqVuaZjPzi1ix5vgL8At+e43p+a+/mH5gChszKY9oRp7rVYQrcICFxPyZOGn0PUDxzx
p+FaTxH+Usj9J/LwNIgdoBAfbyKwIp0NWQ8EwNbV6OGUsmuxbTRGWSdaf+iqaR5RO7tLK1jvyGPG
8bgKqp3LdLPA4DwWiBuULGzrKO4FqDorovxg8efzTNor1lbYjvvbijcU5Ob/yzJShUVLIdVBgDTj
5Og6qnziFo6XOCFtSCsQdcG7p928ZpG0DuOYa4wsR1njZCBBoyK+UqTNcqxqhKMBJIQ5CpvNamZl
LahDbYGPrdtXkjEXDunE3iyQmv7/AUZcvVEZTwBMP3U8JNviOlAXWcz4gdPwEggKwI9tRrfPZ0hG
5CzdRnbuIRCmpDEsNIaaDuTLRlASMvlA4rQ5z6KKN6Qp9hDvQLoMP8nBjSbzu64tdhsXtNaJCAip
mAWqp0nS6gUlT1yj57m9/BCaTg8vuaOPxeti4TjyqwtJd2VKaQlTIpq3jiDIdi7sXCsg+OQ2rTFJ
mBvpbU0exRzRPHgxk+FlILYuDQeCXN/ZGeEilxpBkioe0PS0cUox1RZCvazclLgMpnTDZiUm/PDL
eOAKgAhCG9sysEoUPH2ztRr/Ra3FkySqSQ1/+nGTt0Dd6VrEfZ0GNBs/un/xWKI9NXO4xqctx8Hq
r7qr6wFcpMV3Ik4uq/Ns68NwrZQb2O4FcYycNUH4WZWHtT0oW7FZ+4TXlhROCKKSLBAVOyw71xrw
QQP0izq6VezSofEm9YSnZPyRuvVklE8+Wd9pFVbr/jdpVcXE298/TLto+vzRCroLbZ2l35Za/s/T
Zv1num+U7n7CfLv+//v1aUj1AUHIiHsU6B/59QnzwaikzG3S391rhh+wdjn9Ajhx4MJXIeFvzl/H
heDLeSJres+aISEOXSoMp9hvfqdbg84E6y5ZnELBTLnPBs8ARyf5XB9mn+Rd3YCF8mhy2hLianha
WLVYSMgThLQiPOHYtobraaKhoDtcWjiBnMNfSnTlSFX1ndhvAngjOb+O8ms26PFapcIzC8Zkfu5i
miNOUz+TJ/N7nskBouE7gU2kwuIHBKOZZup6X1zf6jdr8ztea3aPW+A1a7AfbfGck7j7sfnT10pr
DuZdsdk71AygcoGiEuwn1Q/FrzaGKKp88FoUPSq5kJggBUYa5y4QM3HN5AmedmB6EB9tfhiEDYA1
BwHtCapLSTiNUS2Cfhl0pxvpB2I06++JpNEBgBUymVS1E2q9XPjkthqFgSGHuX7yV2Ru47uPaS0W
Oncgw2OHvlgEDlKcCIR05EePQebTaxyuwg6olsflnNE4pdotEU4LuycGg4XpB6wUcO59Z2B+KWOS
9py76zOLyTpGGLMHMMo/BO3UXVA0mkFHUrE44g1sDbTKhdNxQx7of0dzChmNQ+BYpZI62EMBVS3+
KOs2TntAqpFgE4EjOWlyDqHvAj2RrheKNls7A7fzi4B5aBkbN6raMsps+fwmAS56rUkDUiLyRz12
KpE2Qq3HSzSZkYiTEQlzshvv5Hovq2jTW2kIYewSZ8UEEiZOaujNmS5dY27TCRFDRsdVq0kTmQv2
mro5LwMUGwZP3h6KieCL2ZYBgu11DYvsGrnfnf5f0hp6BBwdUoP6J97PfqImaxyFbrO+5eVbzX/M
4RM8m2jY/uaStsMDzY7zKYcJC14hZTibNqh0F4FWC4jNJeeHF4NgZAkTb3ONi37sGoWjEq6X/aPo
v46IAhUqMrlPwMDDAzMSvY9uxBaQyXkxmDMgd+5B7cdObPJzMktHRdBSHX8MpZsuiQboqls/RmJg
DDGl0RttyQg+Fy9g+HEVewia7d0GKSPVPAl7FIrHIcUJ4vILE5GOJAxNKxt/Pa69bcdpEGhqmnTf
1Vz1AfCpvJjMpOOcwv7SGnFe+g9WMG1W9dKB5V+vtDxrh7dhmmSVIppwwwJ8bLbZzUwx/lUCMPNB
J/iEnO7eoJjFM2JYeV21Idk0fuAwsLBGGFQXthpMtAvxPXnYdu9IiK7Gr/b4YkmhmGC/0bN3gFRm
HCL8TWYsVH0nR5PFOPSQTlwlG5a9sgEF9riVM4UNpTQHcN/txCQXM7gKDIF0UHBM866biJj0/dw/
1WagT0aoaKuOKUk14VSEet1l+s1F0qjP5Pd8bZFRcMc4g/tKDG/1sBgTBLKUHWOXrQH5kS7XeWIG
5tdnpwu+NE+ugNkq+fGsKdE5wCol5IwQo93t4Qpzq6t5eFoTgHFSpH0X2KykgAaBZ4Q49UV/WIOi
PdSgaW7Pqi22TEHT7DP91Qt8hNwIdG6PN7FBrlxtLfKcqN48eh6tyXVClxDfAFG0vFDLDtvhnYiK
09smhTnA4XuQpSs5513Va8tuKrPNrXrp/WSjfbFsS8MJHqDLqZeMbmegTEFaLJDvkhibFG9BgoAE
MXp3vWcC0Q/WNZKy3wsF6ef4Mv5pwifn6RSIb5xjmKweTmPGPnuJoT967wjd9ZkSYov4GSr3qfoL
zFLJVDjbdeO5TwDNtctIMzZ00m4QSjc3vaEtj1cjuUWJ+GmcnbwdFspI3DugAVPxgonim4I6ShdQ
pCJuZ45jt0tNy63kIiy/ONxu/ppY65vqjxv+7NHb31urf3t4nVs4Ph/MIb3esMTsNW2pw8jk4b0p
+kvqs63G3/1KPaUwdBS2PuY3UqLMd/84s6TLaPLF0Aw5t84lOmf94usyn0m22agwSDdLCkHI2Xgi
ZciZ6t8nYCaaKIPA1RVNPozj+rCvVk7s2nL5J2UBM6isfwP1Lc1S9RuxFCoulUcYaQXvGIUhIBLt
Cx9BIZ0gAP5YYVVZl3bzLpyQ7W0k2PX/Tiba2IqTPuxNo5nH9ptdVeDEYcYjuURz16HrL0jN/7in
iJAbF+0MBOnv/A2AnzCg6F+wl7uSn8wHBKlMqBKCey7acP3gxolb/+nhexllT+7faGAIZiHqJOgH
L00WVWnQ9T71q2gXuZ0761qtHGIAgNXyrW2d+c5HsFecmti/cTa0+cLWEzrrwK5iZwsQcWaZTnX5
+3te4azeyN71Oei3Tpk6M/UKinD1+PFWQTF8OfkeT3Z3oAREs/LroQmwzHHb59M+aCHpmS7ZgUj5
lWq6eLFNrKJoYyhPaBg4iRbAt4drdREaaR9xwkCdRTrCXtdhKUIDlVRWZhXNhqjGDw3deaqSO0l+
EgrbTYGWKARP+Hlc2QOS6qeAkyLH5W+Gn7NtNUJ8lFuO9Yd9gLaOYLZIvLujQIo0bSyRGnPJoeDR
pwOO2HqeecClJe/JiScV+nMD5G5JD5vwyRGn0a0KV9/WKTuCoiXZzeqtr95Bgl931RMgJ4aiM7YD
7QhXWj3e0x1kVP4C9dxKotua6VIZ3YD47TV4iwxecri0BS87BIdrDArf4Ijt0NenM4if34PzrS3p
hCekRR2MfBxcyBPlAuaRmCJ3DgrnL3y+/xYUKTC2HBi2BzqfDeaEVlGFeOYxeITjIreTKi4+WI8X
TntH/Ft7Nfadri38NgVj0GWq3IDwiYT/piWIr05AtBxkV6MYjnwWGWmSNdD7AUJIeKBxy66NSOcW
McOqZVMBWZZBVKQoU7OOIKY4dnx622k+AO+wrR5j1VOGEJXMBqeSELHAaAREGrn2q1BOFsg7okNU
MJdn3uX8WZUT02c4ZVFg+n+oeaYXUbgBx96fPV9I08bBhnxX7PigJi7HnZXriWFDhiNnnad7ESee
x9fE369EfVJK1QZ65M8dBS3D43agSuM7XxoRDg2HdxGs+wvq+L7LuQWwbXk9DX+0fd6JiANN6aNJ
L2FVTe7VJI+lfU52j+qGA5axYffhmUHns/xzAJ3oDxy6AhsUcuiZtc29DZV/KupUeDBkFQDAhTWW
HIgtrr10l8/3DtQQK3hHTKc8errn+7MEXZ17sXAm31knLWgrXf7J629ulyl9XEsdPrY/tjpHVB67
j7kBpe5q4jQMPpjLPzUCS4Tzyz+PWmlcy6QaGYQBJzHCxJJcsAE33OtOFiioJdR0HkwqlIZXzr5N
CYwIDzB4AMlsJnqxHL5iwqj5uSDsvjBN6T9X+Xu4qPTi4jtSxdbbnkjjE0U7HECVanK7BRj7kUC2
cs+hUrBScGco4CpO7gl+rJgB8lshz3K7ZjrTvqW9YdhGIglHRwo+hKZBOPbHpHwPUPzlBmLQN2QK
/PwKAGZsGpjoExA6Awi3yF8Oa5sLYCwOOBEzRh3bIji5kkcF4oS5redcRK6Jgg6XjoUjKXo7+bsl
f5PFnosBQ/uxzUAuLDL1kKH/Mury1ZIZ+2QpEb8XgrzyfcSlsMwttPYLfCnNHGF/fMHBqtOiqKXl
LfE45q3k/o5W8WR/lK17z2y25h9H0oS6NR1R1ExgzFxElvn82QyhdL2Y2Ip+UhJYfxIzJ/dR0o7B
oHKsrGI/b9EAt7fWRSHqtrRpBlfAYc6Xxs/iGoXgbCTNwNIwLafWlE4uOFLlOIHZJwxTKUe7LPA0
FZ8M1ow11bwX4OFNN9/xBK1iAA4Fypdlx2NNxB5obZKHebZTjfh/P0RERASvrlVucIuueJZczqf0
iWbz1WmZ1DJLmns7PIqiAbeJv9Lajh5OQzw4u8IdDBDOHtC1Hn6NgJTLUUQxLY3kIpzgnGgAWp03
RiDbPLnPKSZDDxE82bCGtQ8ld71nMUgkx1H9GVF0qqgmYNRdG1uSVJVzQfXeui5G7eOXBr8HaP1J
QhGlRJNOT6U2ruDO0lr8YEvSx6hLfYItCa/5nMBOXfiPpDHmLTNCDMaBRyroZIsPmI9FBmipL6nh
ncA1urS64ucuFg1YOZaDxKWVCe0DWbELi5PK5hJ5ZwdcxUXlO2VAEE9z+kdt9S1DcapAgEr287Kx
oR8VtEd7WIziMVseElDhxRsVbH+GxtG+uHHcNWShhQ6qHF2x/r3Xoj9lXJJQqxK0po+M+mqSOBzu
z1I2WXtQ/Kjn1oNyi9HxtuRc/REV77lTbEuYiZQGW9+Q9Pafim4dw5KF9jILds1sQQufzh7yWOL2
ONkT8vdkM6QXm7b8QUyEOxVPNcnbrmk1X/FYsfh9vhEkCFD3W/UXonAVytLZjfrpdjH/TUvx0j8n
oeACj1JQuo+5BZRFCSDZFRAlUYbXUBE1HNstoeEt5+1qf6bxZeBiF5vMcleORV6ArhEqRUbuhG8F
svEZ4IRQsaboqg2wOVRjMyigwUhbWjw4rH2hj2UCPjsmtBMTUpnWsyArnUWxEdofI8y4UrgB+v4v
yEKyDpgx7MFs2c8TH8NFSvNKGRavECJrT+TRH2icQzA6jsedzH78zmdN/yRfd124Ywu+G4FNI1yO
XuW6fzo1osQjg9IbUfKCEA/l6hwKXaZgu0ZBM9BPCfTEyt4J2r/zV4NEqFxB9+SC0nVJDOKBkkSn
oru/FWeywgdUjGMGvoak8MGDCP5HPC0zSQ5+cHiMB/rkwVrc92EzTqvxBEB91C5Z3OlMkKSry7L4
o89CLw2hsCn8dxVqU21cNOypD/cFeBjBicT4C7ysTYXq6ioUOi94Jy6aEi8kWWCr3WM+NIFMaIVv
MBUBfd15ZK7ohDTsLLQrA0QyUES9sngkqrzMfop5JWzJLKtmRHxa2SVmjhLKdoCbn+qlTLSN7WHM
8GDNgtyItNpMyseKLsyfWCdZM+SnWqsbChUVsxs9VnJxzlVeszzruy37hcPnihdGj2PpJAohLTRR
/2UgPlbey387Sba/DsUA6AjntAGRBlOO6yokqs66d2K0SGO7YGe4qO5m5sDcshJ/eWHebvrLZ+Ld
4wni3W/aKZiNrLZPuso/6WdCtKWAoirV2in8FUd98SlwlEaMKoFTYCYE3a5uQuRaqsi15JQER/Bj
qH3/obfwAL91Ge7J9b8lZQVaYNgV/j51sDuAQGULmElODuoOladXtjTfN2sN/XgV+LN/x4U+Ji4A
ugMDTYSYazqMFrRarD2fqnlA4VbxBELLxC57VIHNl88WWDQkIC0u5QDF/K93o3nCPO7xCY3obSCq
YARf1V/m0XWSQIIaaEbXMVnpWRSgT6wdhpNQrGqwB3cA7u2EJ4gHZEMa0Ka+cvFNMPPVXaZukAjr
ZAuuiQCpGzZUlpSQL1XMCkNNlpDIlqjkwwck7Ugkt69XrYiKd4BJL1sqsI9e+0gBeow8VBb5kjE3
E/1n+JQcexG3mD5mfc/cRx/0RjwgImZkW3qNuIQo2sOhyc9bM26ESGYc1f1sovxult2mfO03Mcn1
gp5O/vJYGVmLqrvyI3M+If1FRN3j9oarlq3LF3Y6HY/R2PxgcxNMTDvIINd46amXjp/TkIw2+B5q
oj6E4VnTU35/+X13yZ2AbT4Rs5V+E+nrf/U3ZjjRXWLHT3goeDRf4ldsCP5zNN2sGhCDoA7XFtm0
T1AZFoH6KrOKMsyJNnYXv8sC4m92jnJT7wNC4KwLJg99t+WhiiGsDL5PGHyh1UK1iI0+a/y9xk6+
qXriXdnJaaHdQIoKCr5mC0qi4+lLjvJ+tfDqSnGasUwAIitis3QmkBCmf6dzYzzPSCxUQKFEw0lW
5obQiSBYJ8oVb1ixXJWFwsljl5eEAtTPJKVNYDNcTZDgj7rAmhG9l5fsztz/LRdDCZf4gSAsHUki
iLFUx5h5+VAkqje5gWtpf6uSVtzYECl2YMIgml4dlAXYcsLsHanuO9Q66MCiu3eaQgH5x4pXlZ6Q
90vSkXV8gKs8n2ZW5BWfTalU85iQywftKmhyq753W7ToVATzS5fsPHKvD6vtAgSNsFXmnVDLvml4
UCE/CUISxf3bUCo7k/FHW1bu4LbkETJUnoVakteTj/aJAEvqJp7eDtMUcF1tUxVOibCMXrR2QAbS
f/BJyvH29UBFOY4tXQwQZ1LYyoMTl/8/lEQCTKXqNEJAGIMfiFfTmDNICAgSl4TSElg6+TJ4cCx/
vs0hMv83qacGqPtrLg4/ZWlsVphrjkaSnD2FwXzDYdm6OqZucSxMx3v01CgDO6rPEOAGcA8MkAm9
67lgIdUh3aPc+Hn12wMfMIekoJvbLlaspg4WuOEhr4bWzuqQnoeIMTUP93/g2puPtFJ8a9NLEs1g
C1QpJhfqvx0HswwGJnv6wJOk90VHXaTKky+U61sSHq8CE8hLD6pdXBOO7t5EDKunu1I0gvO7syrE
H9BgbQmW7+XZ+3oOXd71J8Qlw5pAL62NyIpwz32c3aas61yb3FiZCdZ/FOvpUDPk/mHsYjMDrxRT
OdHt4cxcaKzogs9/qxmSeBdsxBvCY3iGEBdpUG7qmMoXob0HBSmkV/7JxAlRwyqwTZd5c5xQHvGH
AN4pccWtGmOcfiWGF8nhgYhfCLSY87n//m9UsJtxg9kiYtePW6gg63Fp1CvncAh3lcIfSmHm4rN3
SEFGI/4z2eeLDbVLUz15tJpkQwmZht0re4dzspdOmiUFVfToDpPvesH0oJ+nsHeRw0ZUQ1T6028a
hs7EylBuRBc/CvjOktzB1upLx4JvV6NX8ccURO+U7lf4JZSx6QrcTksBreLDVv8f6pMhz1mah2LJ
SleOE3BHpvBSyjNrNZKFG7eSZIcueks3/N2a5LjlNFPOiN6TaNg7iL7osLC8SILqaupZTnY0sxp2
cuHOZ2fALP16p3q1XznAwd0vx5USiSEXxNBrt7g33vMn89PGoHgUmz25yxn7kpY55DwByaggc3fm
CrVm/jNswV283Fd7g2N6ztvJi0ryGTvir+PyIUPq561PaH3RzZr1eXFnhdUsxu+PyVyB0vXHRFzl
oA/J8mxBSUoFMKR1xkd+aJF6JFLqEDqCLMMPfyT1e8EiMJYo6GoXlotMZX4AVaQ0pymKmDkeWFcN
LVavyBqdujR0jNFxPeRwXARibgSFXiL4eQzOZY7sTON8nklP7ZdvDqUyC7Gj2jDIpI/stA4eAAnd
miUm3BLKz7axc0NMXeOU/Yh6yK4kxZAZtdjKHJXig2pmEIg6lCdB26g6fPOnRIUz4ni1FhWcU7iR
CroJHTEGFkuQ9S7r32kMPOAhHofbF7LBWiuAvrEXfDZ0nPiN6ehkwviHFZUFqrF23rnupZDi+6IK
Enfbxty+0itV8LowPFMLydho4FEn1AfUF9LROhXwZW/2dRXwUVkOdyiKVZjKbggNOKk4tvycWmh8
RyqBJEzjfrqLYwREVMaEhGUbMsEUkqtaBAfUMzzEWDWqC/eN3xFd3yjTHSl41xouEDZH18KXV453
+zqUDpImQSTBXR9bMYIImkucd3dsbomUGVxer3kWOnNGo+Hj9AYgN59I1UEz9+icaNCeravvQ4YY
u9MR9DUUY8TzkgvwsZg7hw9QWJAcgcRcbEbLf1fcucZJQJFQiesW5Rj8Ou1LhrL/v6BxUmqj1FQP
2LdVGk7AOTHF2u5TiCPoFsE7cntJRxK2P2eDcDrmWTs1NWhvjl/JqjgFA3Wh6xswPds6tH7NmpLK
15U+r8JiWz8tlItldrj3ml6B/XfYaJB8bDTfAUFQlse45yQLjbJ4NlW+bDTUnwK/JOm1be7wJuX6
0HAWb4lvVfp7uIRcqucQOlMskWAKXqVJvYTdoky13ABruDmBqG4HuGAw0HNPmy1HS7CDP6AryjUe
vSZvBL2Bhcbl/SXGG0AkrH9qUrXYXiuGOtc9AEDF0yqQ3JNIrZUNo/CVJB3a/Y2LnTEqrFduu/cr
bIn+M1oN5BsC1brDW2mqHEF6034Uwahzy5ksN9JUADEaRsa/UwTT7Eb2C+FyGGwLFUXBX/2mmFUf
tyQWIfWzjZ6HPZIBYrMbaNfnhtgMW7FtAQtxceopi3sdo9J0dzRw7Yke7ZLVeuw0ekhiO8DdX6S0
n7jmDuWdawInw6NJfyp7YJ1CAij1zKKyGDLnOV9UMdw5LobncAzNDm+nVY9VS0l6SNnbfS17z2+6
ZNWSAYBeZTxvd0folfOe5WKg/KP3hw7CYRIGMENKtHnQzMVFl4dMXP5N7nwnSuEioBMqwzcBx+dc
551kgNV7h+qePv4LHfHkuV1hUhiANEzJmV+Jj0iCTACIOe55i29RJhEpCptYb3hD/ZwMFlwt7ygx
vz+LynMT/jYrWvqO4MOKdsD6WybxocZkhegSNYreWI0Un0uIfDJLsZFn/yN8pbeqj1u9LCQfou0i
ZmGy97TXKVdeWOKGPBr5sFw8tQXEed2hjZ/zY3/3Bqo2zQOwA8sbO7lEgOHK8ZAS+qULbdSM6urp
p7O1ZuBCLytzkByBgqz70I4N/KgO8VB0juYaK9tafLzdN69df5ClsD7BELpxFzTqmFqBteF3Lu3S
k8FxQuaTzhM4maneafIjLL7p32Kvw+shR1FPrEAzZm6DMGMnkZ7CLDEpdRUQQEq+8MkMQn6bHz0s
rTt1ogBh3pgJWKuVDOf9crMypG3ck6Qd37SvJeY3xuMMdj6oeJD3KFxnFVJlSvuxe0bceiQIZkjq
9oa2JegRjckSp+7AfDyK+6jRLoxJ1nTG/mykUZW0pvtLThSoThLw2azAnOTOv3sDenzkx5TIfvgZ
0EUoUZaPJtYSHf0SCeErj2w7Jux/sePzqsC4w/4wdvrfb+YNft58KrCZFoOyIqgbKxQ2XBKMU+le
iz4FP2vlWvl2KuMQiHmxligiVfhcuhcOIP2yUAR6c96EjKkqglg+O7TiA9npVLa8DhahCPI5T9Np
5yh4+LVg55aOVj5N7IJV7qDTH4v0xV+7FpuImWdNVYNnWthrRfooKy2uAlaAXmda/Hdq4G4OMvWP
2EozW5D2laLpirOs3YAhX98XK5xmk++M/Tb0/XErmszzWEKeV5cYdg1L2Bw6yjjdipCGMu7rf7lP
+lBB4fGL2KbnMxivFnNlmH1o9K/yzbGI6ov1zTD+ZsVzAqGvDgRlJyDXYUuAgZN4oCB4rSckC3nO
k2ymTS5TV8hOexSs8oo4miqNaytd1/t3AvTNH39yfoCOUV5edOdymwbzleX+ZuEcRefeXymjW7IO
YNFzMIbccoMXeVL0jrlXwC3BDEFSfUvGihbS19NGV1feV2LLEPAWZPLIrQuEI4pxWGlcgjWBuL1g
DCwxLaHRAB62e26NxLQ0cvtQn1YiwbbZhrwqO80NCfH3OMdygKqcsgAw9q+Y47sME58AKCrzPS0V
dj0vCABLbxcoHLlyRxiF3mU133BDNSayGiRL+Go/kKxSNatkIAtH0g6uHzxzlsrAecwAhag6Wny8
oJ8oszqlIBkowf89BVz6PiJO20rrY0TfiWRE9udqDkqLjUF+IlMP6+PSrpsG7oi0sUc+h22pi+Z3
DhWPJKWuUhuZKuJvALSFVepC/KHPVUe/3HUYaVqi+UmpBr30vt4xDWTAliy5UNgfulZQqzX84L2d
0i0XWanCybF5getvbyGRUfIfU6WwnXC+mzUprT0LdEeADN7j3/Wh9oM6I4WMEvXDty+D32qdddhC
aZZJagBb8BYPA5VQj1nWxCJmyg9uRk2lPlQvcT643Z9eqMfhw+7nKE6bc5TzQkN6JNgeTy1Qyx1e
gjlgOhVf2Xtx3mO/Yyw3AF+tZrg0I0D5kSNJAZmVFBTk6o/66h4+UkR2z2q8A9LE+IMF4c4QzwGh
CY6yZh0Ubs/eLTbT2Xpvf+G543ZkgwQb7q1BpZ5YHUce3ik9QMkH1PSTLzMvBhXGzsrlkCmzjWY/
Pn8uZK0i+ofN6tsTO5Mud5LyUxruJ6EyOuqaNNvMQEsmSfTmHiR/QBmiJJXWl7dGQUYEUsp4CnxC
IA+X1mc9K9geTTBsvTNUCvoqYKfLtMCcZyUr+5r1GlZJWvvzCTnFSH/YbWxcxudWmxbUXJ+SE6Ep
PykNGnqHe3mcbgHL46YIxllnzTfh/82+MUj/DGCNUVA2Bgp8beWzSbKapGGhWcr8/fDQZRMAgtHX
ZUdcTwh4ST8KT1zWUKUFHsjnjOdCJsqfW1xehDrbvKXbwhRqGkHGz791S1up/O+nYjLvoANPoohj
TqK7XL1EasRIoW4eP25kSRUh0sSadoVn/ux3Wq5JFA/iDvQzIi83ts2rI7mmVSLYRI/+AE5Fx7AB
+OQQadp9ILAj1jqQ7DcKL6Bw9I1nAgrGdlgBJ12Azv62dY4WGSvgLgnnH0CEYdI5wmJLmgiOr5mM
YdupLDCp2pX2yfo2+58niWC2oUy13h2cSGkUiwfqebk9q6Q4YvzV/VaClI72j8IZlMPCDHQDdUV+
jKfThkmguPP0uIASz3xTc70viHQSl20MG2QQ7y+CpzClclKWMQwJky/lxqaNMt3S96XDi9GED1PR
QwgLLUJqolDi8BWtGey+4WGj2ppoLLYh6ma0DuZh392isVUZYVhvP1Huefj3RjrgQl//7NPV1O9S
8pxC0tQPBAAIvVqQeWyqjpa7kQdsV+odAZO/Xx7xQlWOod4uHRmTW7FaEFJZY/32Eck9Vbc9torv
06ZG5+umeHM/7cpfhWarnNiPOlStPB7kPQDBBKBn8ZCfLrGGK/YXqRNtxzAPMbBipT2qBMnU+VTF
VnCiIUbzTmnJ+acPTiYvPBIWke7SmV/g7BdGQhNmvc1RbgclM3EWVTv4phaKWw7H0bp34QJ2X9Ly
vHBmBHLUWVtErFjjJzJAbhrsT8aFNPCqw4+KJzWqq4PMSry87Qc6FCEBjs5Uo2LCjcaiVWUvxl/K
8yj9bfMcAiPjBnUUjIlNkwwDRu6+gy6UDqa9WgI+O2/nJSGwb2JZ9ra59z/2BLS2yjld1HxpLXEl
A2E+CpzCR5i87vmgr3bNZekwK3m2YM71cWTWOOJKW8YOtEZWzFqx1ZTXep3MfK7HTbx0Sj0lUos4
2ppS25qGo67w83oxK5fYGNzp9166VJEesz+UO1iKgsG2LD64eJQ9nO63ExQCCwgXQSQNY2v3zNOw
WsaQto9pnNmxMGRQ6QjX4M1brC94+0cvgF8Rza8IplymSGZb3pAJU+J/sMjlU5oKYAW+2PIOPVal
ZBh+BScmUW646cL1SpaxfBeEYKv6WLwh3KhOJ422hBLlJLgniJr/PdTqHUDt931dbCVZCQLtbhlD
O/3rEpF8NtB8Fc8LU2xHuKlCJNc7FZH5lTHf4BtnlbRKlgoChv0Rn6JyjbPXzB6INghta2gVyG80
F3uhcZRU+cAZqLj1o1ikkIydcfpse/eCMD12BmnEXTbFgOxCOG+dHGB6owfCxjceJLBXONCotH3v
DLnCVpBkDVqAGopSELHBaFaKOoXk5/UWrH15XhKrCATODuZpiD7eMCQJdg31ywCbgr0xcHjCvzeo
2D6X1FW39/1gAJf8/Mia/AkfvgI0MdDmD+7iRQM6C783YgeRkwh+HGFS/X9qVEZTP2HwuSqBSs6r
y056A64lne4vrQzTvvhVBCMW6Nsmc26vPEd3hN9UT+RoDWNkMvXQkiE/K4WgzaHWxdrBywnLrVPn
XcU5jeXtQVXldaxEYTfJtzAipzJ1eWWqH1iiPi4b2UCJL0SDLnf7YZdceWMhpSDeuf7snKvn3ZxE
/69Qj4kA09+aG+V1RCSELILWrLfUv4vMkEe9NhVlxKtldrIduOIg34PtsG7uArlvxFKCnQGlUVRg
CoYWAS2A6QnhWjIV4AMjogpeOUTB/+fZFCrY2nGHimRi5lxNl8cId6x72YUo1iuFiyy4iZDK2iag
Qls2VCq2bUHWgUAbllgAE/5wKo+fAqT94fYvaTF0oUZG0a4t1kQkK0NLXYHwKU5CHQIaET3gsu8s
pYzG/MZuMvw3+OAlJlku7UnciQb1czHXC72r7nfR9yVzo4sCw/pLSbhK8GfCV+Y0kkJbQAHYFDrv
DAAusjelxFTEbEpngb5mu3kxjH4+Osy/fd/KzE36Pl+IMBlgPK8AkkW8VlZlWMPblvBnMyrAfSJu
vCXm+f0tF8foIDAAM8LiJ/UIsMq+7gpFurEK2DENsBy1gfJpjgCjNDx5t4/lqqctooDu9526B3Xc
tjBmPBFu4dHG1F+TbvUevPYOBh4XRePQ3+ebSGmdQlKgmJcFJ64ugqCLmRb+02xVLq5NLTJK2Q/a
UZPymASoLXbLlljYgd+VR5PtQlpcZhorPKyFohNuFVSaXyp+yBKp9IsFp7WRowUFMkcdtj+vHeYa
6L0vt70or0B7x2q+KvWXbQhX7Ubd4GL5QsS3x/6CciMrsRjG+bqhY8LIwbj9vG/SegdZ/p8iBvMd
66DHHBs/aXj3yIzqGTwK6e4I6RJYEK43nXH6yCkub7ujqfHS35dDdbIy9QIDhbFIdaFgf01dnRtE
n3LzYClBbeNhbgWnMm16BmYhfe4fjILPubUPzoiYiW0NOyd5d4eaoGxeArQw3IhhxfdaReVX22wC
3fms9t91HWctzzsLEdpXS22NB2UEsVGRn4Ii/AQXcZsUbT94GQyrdbYq/yVVIMU10L2UPrT1ay4v
wmjzG++MrIryTVK2j50bWbG6McSeXXHljs5l5zbTODq4quW3zrpRLMtOnt8VKFYjIxhOkDlspJkO
a8++UZg02HektRXfkFPPOFIYGZj89aUZyfscwWm3R/OqAwe//s3Ywg+VB3/nDOsDSvEkjDYjNSdf
vyaLzBZ3S8pBmqg9PPQifCDj6v9jSwRjYdIVM9QXxKof2ZY60PhUj635j4+GYb0mey8g9g4Bkd+4
F+CKpPfDow9OI4yK5ec61XQ0WOsQZx6FSmlmfbqyVPtlwIlqzvRhtPZDHBCAdItXswfWbIamSRes
H+FnVEVkhnO1Jcq0SMeBNwcFG9Q3GthTRqm4cdNEzmaa0eXlo3fNwr/b7s7g9anq9/gqNKap9elQ
mdI1wN+QJmbQ/PEgZGE6fHmoiKApXRiAhqOOIiNOaB2i3wAMc4le8AaEZVDlQ3D1DFeE96vDhvWV
p/fCVYvNjBUaAOX+N3LhusrM7Y+r73/VYgBypL2qLhgrB9vpJB3DnS5L+NN5H3aHJucHqCrb8uPF
m6S2jImtTkM2LoM62YvOVxmewvsr9EXxfQxZKlB5bKg+hLyXEQW1Qaq9YB9YcSXWlwtipOpWuI/l
A7wNKvk0qZoZNSstSInmgUDco8MmaEtRupOWlqkrkm48Wni15RqZABnbhpR6lGrSeij9nlWzWtym
zQxSzEXSQjuB0BOtevx+pI4tIqEz5UbhqRIhOwWWEqYeQZNtOBmCITPVYv2OZVGJ0Yw20UfUf/3y
th114JA+V2OXeyrVq86HzFCVhO/aG5E7V7ooMQSsHOPmuhRC3hzqU3TZQ5Bi9dvKK3yJG8Ok5Fyp
dO6G5YrKQ26E6f99mEkl0xdtYCBa2ebpCqAgPFQKGvDz/xu9vj22NHfSWIsEr+bBIGhpNyyYSK7z
bEideZZxosb9aH8nCSxTk5QJ4msqLW9VHOTfdLDf0H+RvvI8n4lDXv+7e/2hYlOagusOvrQ+HcIt
Xq7yefDl7iz7DSYJQlbl9N/KZaRA6XftbMrKitgNCqd0LzRVwAkiFExUtsVexDGmyji4hf+IC9hl
WrhDD0qAn9rdgMAt0LuIBtJH5bkkYW72uN16EpSdio2ClkJ+U8Tr8rimVBM987F7XDUgHvKgkL+g
4Brl/FzMTEvRtm7aoYGJZlUWX6pnLTJGjrA3ra7k6IzZEeXdAsgGfcCpNQ+yfeeTq72hKYznbliV
Tt0cgczhXSQ5j3MM+A2uMea3Yq9QpBTBBVXJIXQ6y8q8194bFMZBVCR2sIKusAZwb34UkeTsPZsJ
X0frnxdLtc+aKUP/e1dXQmHPRB9B7dsfr5wDCYSYCxRMen2CxwRLSeD0agyegnRp7idZJniUWozM
supFwy4qSs63S5ZjsLQjZs0h17ut+Jn55p4weMich71kLG/jonZF3ta/T21iv6EiuDa1OLyDvWbf
5sN4g92LhwlT8MZrEewt+08CuOkKfAKVqbJ2ip/Qo//0OqYOKVocTlsQ8dW664PmT2PHkrtrzyqX
okcu9W7BFPI75woqs0Ptifnd2yNvk0bam2FOdcTeGMMXuXZ4Qs+ztXwxQpNr4G6XLzxd6DzRHasM
TCk08y55w/9NDew45jJZwIMvMmgx3gEnaqrQsnu00pA+Hr9/lkLcZdb06WU4/IIrlDgRFliJsc+O
liEoczBosLmgqDpdFDc/QnByxl/mG23CL+vK+9k7fmlGRDu+Zm7dGclwuXr4Oa7lVb9ugC6RGPSv
vaMutce49mVVRbWSuoff3pakr0wGwvZqGSEDB0QpE8DXusuLrBMndXSUVwa/Bh+Sy2iEm/P7FoQt
4s/MFPdwS1wcPWbg4rJLNRe52DRdwtPyBFfZ8EpCX85nrylhLCaJRKaKfXD+nAY8o4kToOgUEiTz
3jHpqwvp+4CbEns4Lq1glp/Bg/S2cw65Ou3DOa0T66DVnPeeuG+8CN7u11J9TDepCvTKZklwX5ni
Pe4rh/Y9msPjTfGETnTbsyAk43aUNimwF97s0pNX07uKZ5uMtbiUVvHt2GYhFdLwu/NiiuoRKchK
NyefG1rN4qrc1oN20gHB5TUeyrWfG1cGrb94prKv8IUT/BtZU+5HCDwXArt0FzKtscMjb17fLSR6
1CFNJSNolBcExfdjsOdUlGLyn+RkKaAUowJBu/8Sa5kvHGI9CZ3fmazCuU1gEv3vXJ0FJBZTZP5o
9BHxr+bKTzcCt1v3BiYU6Q1S3oxVtuqhOjaUb2xLGxS8SF7Oc/pl+WwW1NBqPDvPKqI5JDPUoh1F
Muf5OwJ9L5ov0bD3pVk/WF6YFhU7fHeVNwsWshHR+HFW58yqKu8nRM6R84x7pTxuK8RHhxzhHKv7
6DABp30RnyTAzniXu29JjpkN4k/qFDoAQ9/6vMNDkFnoAj1GIcqUl+rNocJaoMbSJJcGZ9i/E5B1
lZq2+uYcF839J9GgI5FZcMHBGw2i+I2VbSffFDiwyU5pRPFe6HA/fYyRDk/YnABH/UGRN7u8j5zG
rwGQMDKrqMIRGgukBjxMnCJ014e4gu1eWmKxq1UWThQ5K1OY18rJkEmRB4Y1F6mAKJLvLAW+ib+f
qPRFQYFG8/Si2KJLFd4s7695/66yNofWiXPi8JHEpZnC41j+vp8j+4TUWsYxbqtwtlmTTzxYltFC
/OQxt1AHzGNp8WC7T9axTY2K9TLSWfHH8wZ3O6BdgKQ0i/sBrrXQqeCNdCw0zL8uHS80KLYOOLls
f8mOnNl1bNmLiprF8eqZ7CoOpI+3AtJt7GSLqBhdjMZ/35C/lFAOKjI+SNu2QCVWOBY/NrO8g8+3
p1zxJdh1LJUQ4zqrbGYOBUsFezmc8DBw/sZHi96JZrjgs9U8bUNKdVZb4rvAxNdr7MuSKOX6gDcV
edB2gFTtaIIdkZ1Lv1t+CVKbsjgVkxKXJIMzC6qVDD+IKc7MqeMWnYzuOYU1qgJNhkYxzPjAm/8+
LRCDRFIbnlFCiqgYO0yOXPrdihgc0OtO7z75MkvWWE96T9ptJ2E6XSsZ6pJcbhPTVgY/kojI9suP
E3vblELMqzqvBDSgdzGwHtwWHUqteCE42F65Lu1zOPjLZNzYTJbI3MKqxUH9Bv50r3qqqPf6kEyO
ikg4mARC6wEhYrDw+4GkuvlaXOhBmhBceReQiJMuyZTx93TWB1BuLHKCCIA/mGAQfWgQgT9DRJbv
CGU3YfTuQTymvemBM3O02YT1uJIAXGgsSnCwmeRqOEkoYUh399lXuqx0fj+CkUUkToaT2CbmEJAQ
oSrkkDveMkTDUXBAFobBTUY8UXM66JwKU81NdKum1P3HM7ZG0zE42hQFiTfUXMRedq3kioNi4wmz
usDFNZnyWL7W3O+3Xuy+fa7hBicTqYY+wSypl7YFtybfLZalwD4F510lOkr5gal79MgPIbfseLaA
LsG02BM+TuusnvcgkZjIBJY+lwt+tJow6h0hGvpC8rAhCXGV4ti9+KD7Tdk/KoO9po8ahSedD6QK
QKvKE9uHcTYR4PNURrrZVo8dVp0KR8wCuKBOcazEClf22/vqbLbEUOfkb/WLK+qbMw3Skn/YSBnH
vYwjQu8qW/pzHF6VzWrQG3uESumDknEYWFxZbesmuqka+yyJV3g5MFgSSZCFivqtmtZ7ZBUQIA/o
EXCy6hg+i3RVKWtV97SdYiuHwk0PKcDbpr80HoT5wo/PjUYbNsaDwle4NxFhHt5OhWWUYs9JaP4A
HHIzfEFGkPJgX7xOBqS3Tzi/l/TNtPxSgYgKKiMBe/S7o/aB4FDYQywFF3zxje3Z+j1kfMxuGeNI
ctT8xslMl4MqLqjsjSR6WTM4Ie170rysHxFTqOXNL8aSTS5JUUhL/9vKK2sLJDv7sW/6HdbiYFFN
ttxOSbZ7eCDiRrE2A2PBrfa741KVwiY9vBw5wvkrrl+9Pb0ecOIPgRFDO5zHN5rnLro82xu+XYkZ
TlQsJSVzNRIeRBP9B0s88t+pprAzPZN4+HpNawfbYTnXkRqA0BBuCyO3lzirg78LjjYzTXbNb3ix
Bb+BXqMsd3fyQveTJzVgILpAEUZQVdH/E3gdpY9kjA3honKv5ttd1ybckcPZqAOSejUBQh7MEsqo
EaadGIcAxKtTJbCd5F3RdPpAeM04QCODfwMTgaGimIJ9YdoW06mrSqhZ2cxjXfVnjmYRaV8ioBd1
5w2gNRK1E85bmmG4X9q/M7gcyyghB5UDSVaRtLZoCdx9/P+bDoGsKpNP2O9qsjry6eJrwpOcIj63
gGHmA/4/vVg59dZSwxxX2Zt/je3PC4icEXWS+Vbx96Qz146h47GlSAI2v3LBMLRmkyYGEhMaL+yY
xglsmpLJTNsxcfLQxmvB5Mq7eIviKtnBahtGREp2lNJnet2SypMsCfyGgSIsHxl7xg5OX1TD+rNv
PddiA+u+GsP4nbLO1yb8ltk2g+02HozCd/J+aSHz0kEzNac0u5Tm08HdduryynMT+igFQO3cFXVq
dDE+Qj56XXOm5e2bnBAhCYrJruVozVzNv1mwHFO2gYAlNXCJRkPQPQOlo8hBLnt9ZhmAKWm7Ch12
FYGFIjSZ65A7TCORey8r8Zbktgp2D+nT23DtvthKw2g34n76BBUUa9mVJdkxJabpXjGQaWFbnA8z
1Zrpyw3id6hmCQ3wsyJLRXiQV3Qd6xuQ6IUS4MFxsKdrvhN4LVjtlcrc//KaC8RYDSNaBsTojEwB
kP083IrOXnNThzNKbgPvOlXUzU+26/1VNDM8CmdH7XTjhO0yshyx4m9hB99rZU4kFeB8FctKFB7u
Iuaks08Q+8M/4MnPdvISo5BBQxGgDcqmC8sIGoPfpo/mq6AeWUel5p13lauyvBv22B8Q6LlXsMkB
hwQrNJm8qZE2EIHVpBUTFJQzZ2Bmsjhdi7Tc0Q1mOM/IpmrXmHaHtsUSHQIhERGKvLrx4TQ5v08N
bZuJvO2D8o0LcobYqZaXcHAaud/6kGKk8D3O5QJaivzz2+nTbJx3P95Aakddwl9R93fB3kHKNbtt
Z6KrINhHMNRySETOHUyDfcx5giUwCLLV1QgAvIkFtiKdOJ/uGh2UEccR8gJpg+vO4QVcYKn8Rm0j
/PhOMXhbzBn0+/75eErMgfdz8mB/qWpxtBgrgHYwGx8PspoZaLYPjRcZdCEddq+9O2npWqJbikir
G4GATYXJmFpuTIc+oNXqXVz0h0aJJXi9nku3/iTVNwOhfXa94hKySedx87ClqQ64R4GiSVWdqvdZ
PGDxcoClsR6UpbVgc5PhLbQSjnQpTlWsEf4GzPDug1vVkrj8qqYYSwicO9m6YKDoHtO5yA7t1Tel
iVe2Cey/ZD+GvwgNdeuYf2PwLdeSqNSy4GIMedsRVsV5OmC9ssPFv8WrYCdCHmX7H9Dgc8drnuKv
bDRPUYD7ejahWjFYwLZhuymfVM5pxOlTVvE9POAsViYpkg+nlwPtFzrDYsdjgqdHbi9YFD0kKcpn
Bg01W6lMBH/+n//Hd25TkYfNMdE0ZhkE/OtkYtTXLjbHy7MXrsAN4iF9CBqmlwbodZCeU7M6j76R
dcZ0B5saHulxPvZSlTaejW+3X+ibBzotTjN+UMGlZYImQU8gPzTnaO4NP9F93xteTiQNOxD5hSei
p2lz8ArDgh7w1blGk7WnwS9nCNJTybhTgbaQERO0APpDL9NR2OCKK4xUdGbQQcVbFdu3TCinxPek
gszBgcF7H+DHNAK+jARy9gZCnorgt9zt877naKnTLGLH5qInqjWzeHxrwmy34yIOxEVBDTcFrYhh
IyGHFXVltMomcfy0bi7LzQ9u1zJJ+pdVcOCTrLLOf11m2va4jFSvVuTWcM346p7uXBjz3ZE2bUt6
mj370Dq5LQXMkFyZ6vc7+vu6bphdbhnGZjQ45Dvzhci5wswYw723/OtVfvY0oauBkdZXFWeIhkX6
iALSuZLVXhISCt7WuwutqbethNyuR8Jje8lp4zQiSegaCCA/Bzga0aae+aHnDNZcYbtCFhsEwMgY
OKa5JNHRoVAp8ogVY3dd20OH62nPdOxpmLCX3jU3nOjoXhfubgdGbgJv9XDYmxIlPFM41WUjaYfX
lu9QHqMi5zjhVoO/11ZXC8Umq4Pz6LplgjoezEXz7iIdJxpl41CKChzu3mtNUy8e8/5X2dDxC6uL
cibXn8IGUGmXklWNliO36yxZAXHNx6BvNpwWFDawD6Tc3xYen0iSZVrrGuVavT+GlMUfLqIlCRpk
WdMyM5GoR/KzZXTBrTFKc5GcyJ5VCcCKUnx41C/vlQmvToHDiR5uMI6SmDTVrvoPdYnKk2Z7ObmS
XU8Ifp8Dg2/swBu8b7qh+ruA5bhcquII7qahJ9hfOMcbT6PXKcgf9SXxDI0E/wYi3imMmyxmHagx
Y8l9Cw259UcR/zJqbyORMwmax4gf43pELWt4L0usrk5rRzm72cIReBydYmCrJqDwCHXhnuCIbDEA
oFgb6lvt82688RP3DJtXhdtSMRpEYIg//FxxXyy3A9Tb+bOYEiP9mTihTeQUsu3rBIzcWd/+SXQf
pAyl4WNy9C4gyUHOmP3zcSFYznQr6tlVbBMZSS7eLzx048QcqDaWAoY6nM+/x7bd4xGRjvneyuLp
U8WV5zNDypySiTk4OSBaTd6z8yE314quvlWOOtpsJQfRhwGz/93imNy55Lvemj5cyW/+a86Bnp9j
e8zutS1Tv+leEO0tlCWKoGptRXqjNlWIailZX0ndoEojYs33najPA5NZkcls2eUQzB0su6xf+i8o
MDFMNCw+dXNhsPQgES17Rziqq6FZMO+8FnpC4pjWo2dCcI9W8mo7XYd87oOk2U+j4pK8gdGXMJBK
W6+lSP7oZRuKqxWIu/gkCa6wrTcl8Nj5z21EkC20zPbrLM0vuaYvcv9eCWVyWFTi+6rd1QaQCJrm
Au0bL68mzfSZqiOdFxpCZlxfCxajTjoduTLS+28Mw9s4dHp8MvNw0xw7idmt2RbbNPzGftmj/qaq
fZVgSEmsYzaQBjvd7C6JGAYte1HVXJWw2Q95Ti2poosjPEa6zl7HpQcAXzqQpifi8osAUAKpxFZP
sjb8VxYcgg7fyx6dTTKsJZjR5gY3Evdj8a4Z64BhaX4QXN1TmIXwd1UblmFNQmSmV7yVIE/icj45
Oqrauo9Yt/k5sTvJhixx6TsyIzVDfFO+Tw4GcANytNC1ImxyBrdWNroAMmomHNaNdTQ+SKMrdsP4
Jvdcu3ztt6y5RoywL5xdlBvqx7iqJezkrAMxm7nTv+OrYXplprF8pYEYO80BQ+XSSfT4/8k0HDrL
KnhBvSDOg9eRlPH5sTUOhsqg+6MAGFeSpxCRlDAwF8Hv5Nk+ni3VY9ROjq5S70mszFdELtAkk8pb
aRTRQ+H8Oh4F/rGYb7EAV00GrQ5sryDicPXN7XAUvxVm3VY/EYTZwBvuFkfTdmShRF/ryEbwUu9G
FWjZRhbig5HoIh6GlH97tXmA3lhqgTPjuIqp+i4seTkl5DleSfIPb4bRYtd1pMwVOldmiF8BS8qv
5nEu7dY8ZjGF1i0nLlFuFyUKYsH+5QWw9q59bqlLipDqXa/S3L81HDLg4679mWEXnd0PJwzbQqiQ
Offp+voMTlv0tO6GnWpXgoaHamei1aczfQYOdnQOnvRfBU17lVJTOc7LWf2LM18NfaTyWczXZSLj
0duPvN92Y4XsQQS7O+ge/ggQpF8uvR4BGeGdDrKURaNOR0mkoTbLED89EZZyAp8pwaPq01V+cVu7
YCDcacfobP3Y4qdcycBHWo8bJBNW2jWSpvWfGKqgVoKr7fYi/DdLhiDh3NOuK3+0DyAJbNlVBrPR
uh9FRtz6FFcrCCeq4xcR9vpBHW5i+vyq39s+plCcvCaC4Ccc7y1OCz8CCGVdTRzwlmIxDkLyTITQ
MI0vvclgb3Ci55bL7NFJaBjVsfm2DGue2Onw7std7OYIffh7mswNNvoTDxVYUHFu/dfaGNDG3nyb
/u7dgrUDzmINsdW86mm1PR30WofjzfiqTsOF3nQcftU4RBgcUX9dcp2RG8GvErfv+L9ISEmN3Obi
MLcEvDj28emyWd6WlsxB67FZdZwNJPuecTnEU4mNayaY9FUWGCApf4CjVaPiKHoj8+RP2j1VP7i/
dhDctyiFZHj9f/9+FtGAlVYp+2QeeNvfSYvLkIWT+gZhzWylO3gGPLBt6wLhQKrz3yELn5eiC4+o
SryzC5qcYoxDGBo8nBbfK8ZjJQRmnlNerZKIiINIKvsqMhi0U5uYHpa8eUz2T4TrBA5tWul26dN3
CzwQgqL+7p9vfGGWokbeKdgyRKkGLkQYPcoESn2WZ+gwGo7+CDD8KbomQB/9EUYDKRDQxOcakRHG
4otNSNYTURR8MQjQV7BWWJo0y8cHHiC8q93EvEhpFjsdYLasyWvtgdukWqJgpgAzpe3K9B8hWA84
NGB7xKqXsChxgP+aBiZ+LQ7kSQmYR4ejIrcP4xTw6gFhRhhw0zRkwBF3CfaihpBs3SV/WYFtZ7lK
me2rJTKKvAGrA7/FwZerr8xL4SvLoLERvau4z80KwfVmjf/iFlnpEEHIO8MOqPijUeAM6y2eCbZl
UVoHcPVuNeK4gFgJqHGHf5Gd34I/2jBAZqtpHogS+Ib474RU4wAGU4e0kVFI9Ce/g3QGTN5nLK88
QWAHwvOeJ2Z3AMwtzd6AN8jq1D7bcm2NgVU0eiumwCtR0Btn18IHD0LwR0AWU48M6pYXGeH9CVHq
9LrUGFlCaLoSYEo9P4cHwRENcRHRtLphi8HMUZCRzFqVTjxBsnh2Z6j6b8u2MbUith8fkdNvj0K0
20r/MzazPiIjszeJaKpleG8P4a6SeIVv+tAMgP8yXx7M+ZYeD/moubpc8OzZmV5P7MEOkWnpkyF6
OVxe0vHAOJNXhvayspXNTMHxh4Ih6s++gZhSBNPDaUaGDLIYD4QMY07HhDb5s7A4Xbh+Yhud0L5V
lm76EOgddxzXYLpJ06lomPoNX7GnKwf80Dz36/ycmQniV1w2M7vQKs0ehw+QFEDt+QcKLH/gzrec
AZ4/Z+RYwaRZIXvQbuXernVY4Mlcut4Nk9tvqaP06v3vrG9/KSv4T8/MJDwxdMsxY6mplKn2bfj0
AvUrgz62Y5HUqpN/8jzN28N5Omflkc4Vi2ttjKqtHmvJi+0Rla+nhPlDvarH1m9x2kHa+yNJnEK3
RYNXr1HyrPRRyN2hdEEyBmaTCfOqkUa1YDsdysLs47lSltaGhoX0AHV0ISNj99DpPfktv8lDm8rJ
AN6kcM9FzijG5jrrGiO0HFTb++C47YKW8eNLFiK1fY/wj3iasVPUr1aEDtfM8ClwlrKWUjv7Kx+K
VNo+fjflZBvl+ap+2mt20uhL0h9/OSmXWZPvVibtj3PAn/WJDVLA7PyE8sBNcH4QL1NORRlJJGR8
XiJZHFkIBNjZKFDWNZbYErWD5jzApTrCKFbtNXF4DdDN9lkr1SGafcqtQicVRSc/ZafYbvMJ7oJV
l1tvdMyEfwMRzbOZmp5TO8tx4CdKNDU8kFgNijTvZTrBAHf1rm9ZZuljkakno0XJTkAMHQyNt3p9
JJLmmJsWJwy5oi4uuUfV3omD2FISxR/uErDTfsFLbwZNld9A1cyVUlVlzoC+p7UNYGQm6GXycHyz
/Vyl/qdMUcOTQPZeJ7QcqaWMZfrIHaLjGnjphkFYC5FRCZ77wLxI6JbXY2zzsI67e6TuIXk0rcqs
pBHbeVq5fFqKVRwz5SzraqYs6DZfKpQWtMKE8Bk0PitXjxnnbRfmP3Ru0kPs5CjOsAfyEFb3mymh
xwf66ay6KRoeZPO5YCm63xGz/quN+GKDf1XTTiEtpJ0AWNs3OzDK4GvHfMK5YPqiGNAaV9AY7BHF
pdJZD9CVYal37aBy/1bVvA5hszEj0IngUi/nUQ+6JeE5FbVeKm0B0mlkW3+jvHZgMI/cGZ8gf+SF
i8vcXfWyU7+e+i+2wOHuIKa5N/qtqriDO7u4xBw/uJccY9NcIRlTXLdkXE8pvgfTDbIKRx+Iz8RG
wHvgCOnn4RaTjn7QtI0//SMCxmLIKonXvc0xUTBJqZugoU7jDLDnVFq0Ryc7u5zZtaJqAkD5Mbba
VsX/huV+7Z1N0HRJ5AsNnMWgYqpKYiqDd6L7nY1vhKxvwgxYkYucYIkXTpbJHmgzX+b5VHWp2fxI
+go+0oUbTsp05NwQ+Jj+HGG8TtrD9phIQB2dw9XzVPfQNQTkZ1mL3SKnM2wMTWeVqY3Dcmcx70+t
zKChbDxhCsg2Bmwol7nKGjfueql/IaeliSeeoipDj0C2qRFJh98NLp1yit7uFpLDltZ6lTSbWsP5
SmDFCm0vvhir37/4Sn/HhcWc/w8t7JTUbJK6r2LxYkfk3dtBoeBDo++9PiUndRhS83QSDozR8dv+
6QtU857PgEHSVUjsTwEYa5IBIAlW2Y2D4rk3wyXf1stYtCKGbLgNFwHpG4mM4H5KE+3W3hnG430K
LvBudfn9JV0k+xg6UgWGdzKssQEvYAdZzS2FBmaNJaorRmuL0fMoOguZQ16zPOuUDzKh8ZYdWNx5
JyBy+iaiE4i2PFPtenapRi/haGCufAxYpAdsKpRLiFV9697ViAf+9GiQIb1XyV8G5JLx/RhCbt9o
Xmak6/PWKZPSyzfDB2KthkqdRsXW/z+sX5Rr5Ud+MGTQY6dzvTJiGDltBmpd2aD/szikdExH2KmL
5J7CzsoX80hJnQ6N6tbjUF+AQk7RfOIpD+4ndpcIJ+jrGHjwJD0TYRXnOZUCuIZn0OgN1F3tlSEA
9VGEVQQMaYUE+ltJAyAqQ68zH9YIBpncwcdXjhPPcx2RXB/9NZiFZugbCiHZwUzua0Hi0sCyCba/
0ib6Co807PZGeLwZNbduAkVGP99Jwsls+4Fut5xGAGdAkuXCnNK1R9jnl1fYaAPhWwaJQnOx2vtO
357uZFv3RQFKEaydT8AL/0wb6LBi0vARYyOqRHvtWLeRoRMAd4lYvv/rK59TQXQ11xzDP0xdTZH2
2esnpt+Ov/pJ9d0sbtYPUWMjOKbcZ3V4idDacM8zDOGZ8Gn57ngP8rH0euYk5LFd0i7ruZiLS2pV
cwzFt73E9NkKrJaafUMys6m7pGeUSpSlDA0o+0LDqrjFPs/cH5nxTfku8P2bMmQWeluw1NT0Cqtd
dBlbQggtAL8Fr7l0WCQMakpcdavh1ZE1I1+F/LbI6fCnA30qdU0J/1JzmH6HyUld5CtlHTc2bt27
mVzVmKAzhLNwnIzfXUvzgEOSQdNIArLTHRCp0Lj7z7myyGKrjqKotagKTyIuYsZvHIdf+N25I3hO
wgdsUriEK83V5U7jDj9WnYalgrtKv+5xb0MbeR0NuE6mLoCLMS+GC/KqSrAgS9Y3wxp/s40pJ82e
YImbf3cwShJI+IkJUHbMLa7YryPv9JdI8WvKdtsMIInjVzrAt2aj/GnZJDOSAZbAprhsumJGdt2J
nUPoS8xcq4bcGVZ/b1rowcrAxIfSgqccBOTovBIhpb2KtPodCoN7HE2N1Hj+0wo7rVeWM7frI2lV
K/vUPjeXMRetENY43xOTdiXk3vctmbF/D0cnhex+k2WBiwq9zER2oHYckvDqv1Fe9a8i630qZWsj
fBpCFuVYPGbYSz0vSCn98x/YNnuJncR8dFm+R3ZhAJq0ruB6YuuTHk/wcaJTLwrzGWVnzLGBMgVU
Sv/wuYcE1G7YSEIijv/1icTW7wrU9v7H4hMclgEZtMztZ954lzt7uC86pgmfjbcdtOQ84znyJbOy
GHMW43UXHMkn/0KxH/hAllNbCwH8QZQvMvXuuoYWZcW9DTZrngXk0QRL24K+ZW391VAcJ4Bvyb23
L81U6XluMCDGIMad+punoELgZpce/G820G73vXSmQf/HBtkeU8ZEb10LwH28aCEbTTH/QD9Je/OD
k0RcL2Z4A2Vp+K/aVHPJVGR4Ahtqpy0ZtLZlaALTS4C41tlQJctLFdwxdV3EMBN7jEix0SddEilJ
aRHt+Jid0LutW7Ms9Kad+JWdhYIXwy+8v29i9dBzQv14twOfljQI3xbEOz0PUatUu+wUBPJzQrVi
WsLI7QGSHTQiIk0jM/VCYPyGJgNgewJzBnSAejwsb8h5mEnku0/qFkxsGt96lwMUgnuqLZGmJl7l
N54X2JTPQmUB5JBSdNXMd+Kg4rG8dE3EnAVsR9GdBzPwGMkPXUIwqOvU/eQGWpumY0mP7Fe/Zc5b
rMbRBEspwNIife4h3K0uEhZkahVPMMIrqTmBAiJsp0LoprZSuWkcYYgWcsJaBUf558FE8jK/tGb3
VxutsAJrLmIfNWD9XrMqbyvWAFrv1NGjG0BW9Ztt0iILhYI4UuIeTv5TLuOi8i9GlOB3SNrXUg3G
OVUfcrLokWYVAkUETAo6Rj/uipYfmBZ3fGxkgugb1bZl9H3VZLRj0lpjvB3FUFOOjcGvJzx4IyYR
0fbo01PecqhfuV/4GzrAUNgUl67jJJRgFpOrD7h0XpUQuHl+HBoBfNhiaGUNf8qMjPGKLNFmY22D
0dJ+veT0Sw28qAnaOgpVHMAIbPpc+7k6lsVqIBDdY2Pm4ovaNprxl5tkQZwRzvWmXNDtsR8h4Erj
X9jGysxQs/HktiqcOXIbxydU7Sw+mORGiyS3uPoqPTTjik1KZukUFrXLAZhEiuMgJvtb3N44y/bD
NbpqFKAv1+RvDVi0Lueiu/PC2PuvmC1GGvaA+a9YoWN+DaGTutsQMnljlBwFqZWIN9FlnuOYRZZY
eNcn8AbrpIwCbZL0qi7IphiWjeiTfiHsTEMj1AGnpjaVRJhapi/HU3NpjId1t6jIX8d/CZy2i2SL
QpdhFZP+X/1QCjMx4Pa66TmT4sESoOX+8/L2vAJgwBH5AxGC6IPBqOihuXn037H9l6X0JXtVj6BR
WapcmAQGevjBUlHY/++HLWllOAZgNIb9n0QsArj/1KegTqEEMfZVCpa68EuikvzzrznAw9u3s+Ub
JNKq1vvh9nEN2jy4+7EuCnzUdrewJN1SwCSC3TaUoM52Z+VU1hHbRy/udWkduZMaa6kMrFsfU+ZW
Pk5FaA+R3zHan9Ie1hNP/uBWmS4kyyz1RcI1dkHA6viKbVFxZZsFTpiP87x/vY/EQ7Jdxm1uLPIm
mJOO9e32TM9wG1VwFhmUDsHIz03Z5EYfL2lYkX8Gyc+RtrEDAQnqgsheFWhYl03pIDCGSnewvmK5
WCxN1INAE5X24K9OnCQ46QuocstEcoiJkghbwkOXDGiOisZMtW4Gq+IGxiOzfdoCDzRpNVA7FX5i
xkQYaXRJIIVunXA0E1cPFqnhmXwE3jk7gP+sb42jwyLK0osJm5SsNqx4jkKeC69iYz596ymkOs02
A6/huB/7MKN+LUB4ZirzGXfnfeuinaTD+bVjg+7FqRPYbkvMD4J2mw9LgIpy8EGqd97rfcRqPDfG
setgaG7RK4ooCTwTzMSBxG8EcDVGqXkH1H3tR1VMUeq/XVMZPA9dngmB18q37PoPNYiz9Y1umTgb
diN891vaXRXgmP2JQ3Q77FxCsQ2GW46RjQIiOYa3sXQPlLR4Pemm6pnR4f7v0rZ99qkrigSzh2Vt
snRVc8qshaybZ0exTH2FxIkICmVsPrsQKR98gmCKU1I5450KsZkoXkq5zkxemD48XchWZ1Bxa9cH
xxDc03EoFZoJPbfljETF1AQCCtAl3lObcgz65VQlr67nHVjWzQlFgh6lFWi3Q77bOEiVa9kximmM
SKitte8Tk598dPcTWXSCLDCRsyVCNdJJGCdCDnBQ6xZmGnZKSWoBhsWrYGwa3Sscw4j2QY32r1+k
Hy6p/lbd7DDTyqfjluXpj6jT1KKUmRAQMbBZ+nu7I1FvNYVy6jVrSUUAR8+ONMW4CqFbkaH3joqn
eHiwF5ts9hXvZhB+x+ayDzPDN/NaPZYhiB4+QdPojB3ykugxN5Mnuic+mPk5KZzDchG28+EcHff7
UU+faPGmmr3+4lTvkClAfeDbV4DgFlIMVXhhagkBtK3tV3G+iZ0/1qDGk1+vziYeMz58CKHBIIj7
GtFT1GAQUZHxrlgG2rG/gU/ZegOu5UK8NVXrNLaphk8PzIO244aojMuLpZKpV7GE8bylypRdIlIs
DZzyDRmk24TLOzoExFZPTuD9ywXHa6ebIs7dgmBHz66+LeF3RxQnkzhWjMeqOZfsMiaSaU2K5CWE
sZ7MFiybfWNB/Lkk4r2SMRO9ppQ5+zJaycRsu5GRSF3MgdPDZAjlDdcBWiNKDlFcuammSKUs28XP
Dzp23CMLvGQ8shHft3dhq99ywxsbgOO03CJgLZmVY/5lyHV6MDqkExLyKmBwP23o5Hie2QSNFng5
sFzMLvIFivj8mw/pYlr3kc6Rj3wBqaP4jF2d7SQj6DgaufGscNon3O9ExuhFLg3F1KKTitLPPcO3
L+E3DkPYGkyQodN1KUg+tp4yvEG/8TVy4aSnUfQ99SNGKPhPzUvmVL++m4CWL+34XxlMyy8KYsug
C7SIFu21hCdbYtiCUi6ua0di5dHlXYDWwD2CqVfekIYXI2VH+kroZAvb0t2P0ziGtMi9T86LPo58
8k0YhmvOl8eQsCnKu0L5M22dMukgzX5sFRIRSyvGJ0EolvGqWUVYN6DghY/ATXZr/w7EifVFzbLC
KlpzdaPccrk3NF5RY+e1GxNucnNdwldIZr7bTcxa4OfJii93Pn9uW+rr5j24oG7b7CfolXsGbMzQ
N4LgmEhAdqM3qP7wZKJJOsT+WqWd10FxKy2nrw6DJdvUNVp75hGsX1qPRgar89XF0etsMeMEssCr
yzB2f8ZU0mjoGQWV7OKm4tspz3Gm78ivdTeelzNTgeVm470R95kspxVsyRQCo5RXuufCKl2+kTHu
AAxTOPt9A4I+37dZEeN/gNWbX4oBQ7UbGTXgNlDtiHHt94vAnGHWPOiNodCURDLVJc0wBTqUbcMM
aOKUBY0C1e87cxolnaG0B5EgdjbzgpzkJy2uB9cRfJzShcKQhTa7PI7n8M+cvgy1TcoZUP8Nihal
EqCsPQWE9faruci5jtpWeJh7DdcbGUFy5KdWBUs1jjAjZOZlmTfxT1kk5cw3B7uVmHXct+fh/KWg
n/3NRQMn6VIbPIRtjLkPAoK7QAvZlXsAuWGGx+CuvR63ChoJLXGosV8QKTggTscRWAiKAFbxjVZb
bafcq6dyYClHqq7JPsxe7XhTz/VrAlK/SvnuIGLJN+faxuXG4DBn4Nyjx0SkIqNMp4AQph8szQEZ
Diefh8jYQ+yYHmXBRn9V7W1Za5likMZzZy3qt9vaO2zyGi9wTy+cBhPRVKvtKXSobbymq7J0e9U+
9X+RenwIc18Np6K702/flY0YXWDUr76jwi8qdpVTT7Rc0q53yEoSvTNvpfest+idpuxJtsA3piOh
QcHnbVj84vVvhDuNlLt1xveP2NPZ6+LFa9s0W69Y1algD+3P9rnp0KA/Ha0i/qt7zOnwUGhBI7/p
gk6b2udPrKhT06bP+8pi6V+ovPX6JDCZffNnWMLPhcTzv3ByIZ57SS7lyT3U+FK+F+vw+XXVAp3k
I4PMOfDaX+yQusOrywTqV+A5Z0GThjbxMP5ui5I8QyPikgy07l4hYiVUREyRg9fzyooMk++IlUZ5
hUfxc5p1ilSmMmjGvK5lcsgYTGr1RwBnskkBaXY3lGtaPPMr8wk7JR37gM+wmzt+1GALoLgEhIDX
6eyQ3hDvE+5fJRnUns5O/0v5cuBFwlsVjO/yYs5H/rJT3Fi129LIrzz/TPbajEZjrEXwAyJBZRb0
uH4sZZiKrlKyiPW6L+I/fAglS0EXWu5UWRyFyDcNUC/71qnLOVAaaAEfbvZD5IoRAehE0Sc4j3Da
AlX37sD1YEWooTwyfHYcbLNVqndCni6NtSvekvRmbyN2Edt1CWYKzvc4S8UsGElvBTlDVOVjLDIj
2CHJODe41Pcqk1Y0iNkBQcKPVDFGVpQ/mI4pKZO69b2TgRUKeqNs8EaPZSKGVzxO4DDq12UDy5ub
m35IT8wPz6fKE9XnkkuCWH2FWFkBkUZVkCRADkhQLu5fjtdPRIKBnANlcV0OQcxabZWi9EPNefW6
9D1HNg6OPi61ujCvVj3zPU4/orGOgg2kjz5HcMJLXo8Br4F1cY84TRZiSB1YMMAMUco/gKPTJ8EA
Jik0Bq0aGmW2P3BIK3n9RPp7dsl63mX7nRxdhNtJT4T1Q8vPqVT+qR0MgitpNlRv83ATC3wd/fye
9iI8+BHADUSEtXZB9Dfo2ggfFPnFDt5y+vLVpyWzoq8jKZjY/v7BzjXeDlxhcIjMsyg5SAdEyKj/
8hWup+f3e1G7mZLRrQSlqhiwstz3mo98Zc/HrbMHTeHplWrtwJLWsQrLetcHsmrLBnPoglvVaXpE
AIPXDiM5DcmO9FFJG99llvGYhjk25vXYcBeWH60FpJjR4vZ6QzQm2FHsp35G46FmJgMgNyCrphxC
mtOaJP+R2lEJABPx0M689YETSXPem8hneZJH74OFUBM4PnNoY7AdiN7Pni1q0cr7Y80h603p7oxU
w8nukZQBSIWYkUF7Rvwk9j9yE8lYnBvRLWKikgrLh8yHDcPtU/NbQPQ06ZG+o8Wypf4w7yw6PVHl
G7RcEkZ/XQi1bH1aprLDYmhexhMG5Mr8j62nG4BrMvRthFk6mdvRUeFJkKvzYV7gta8//h1hMhSh
k8tcayew9ZEdP2Yui56V3uJ2C0/rgH4c0KMqZkdlfeRnSVzsqsH76RD936LLY/dBEKJwtTQDWRgF
8tk4QGKD9GW/o8TJIw7zrZdA92mIOOen/aWRNYGEIY1OvRKjX9Q3BeYFQQb8/ZvSkH8u/2Ro5aAk
/JVBkFJckEpIZKxdwKKXAvsadnfXl52/yTffR/fZN3HHjE1uPEYMOsIwncxU5zV2jErmNWchC/xF
Ow39Ep1isrUxmI5rfYDnwfdjjaYVXar5VRn5LQxxX0IwdFi3N9r8yp6aIT8mqLTK9iaQOwIh3zak
1dEG4/i/h8bE4yR4n/ES2YQPNIWIwfYg6Q3r2pLKGSIM+bFS3Rb5ffw4aX85KxIuHWa5psPu53NF
tUkuEklbtaaq/Ri4iqoZd7YzTeMglIZHMfUgRXC7Mox2pVTiATRnIp5wZegr8CM/o+tyrJZVOXaD
PHQ+5Ysc/MWfZW0y8lC+rbwN4qy6yXjQE899IdXMixRf6/H7RiihRjYyqYt/+2pWpvlVf3e7cUN/
+Qo32tTeV7DtgXF4nKaWUaTT14ItGCx4f+cxflowsf3SPJi4jBeprs6holOGQzeB0zz8owb6R6Ck
9wsx/rDH2jVa5KR7x86VG9gG2dWcvXjyOUS+UbXJbp4BiQTHUkk80hhjilygfSw8xQcMYKQCVh0P
ZLzTlFRGnZaojvY0KEtU/pirfTrTaDaCgDiOQC8W4mPzfBJ+IdOLsRZU6Y51DWX+ocCCCEfaS9+L
7ZbpLQ6EfG7OEPXsRRMO0UdB/Kz0t0HV+r42ICFVsJSrMPVgy8/iRcrgL+44w/Harh9/D6MgH+fH
2FXC3REhhfqSLa3eEcnod16QWjSTPfwugrHilAyugrPON8QLRwbWAFSukl/32zvrvWIHa6agzXPm
rgM0oI5+uCZWEe++5v8FwC5zAck+qsmjUxWIKeVxjadHPI3zwdpy365wag2BGd8Dava26SrTdTOP
jAmEwZRPiCaayqhGGSEiu/STeIbxqqtP8qjVvOCehn1uTGWFwOC89z5duJ3w5fSBqWMcYxcSmkwQ
5TfIX+L5ukEDWEIj5h+4p2/M7oanUXcq8e47RvCJZ9Fc8dg1sfSTqo7E/hOasf+ixT97y+McAibu
ymKk6V7gJcHs41nkcXhWKoNxK8AO3PQqu0OZk6LZPDLcyCwJoUV2DKEPXawfAJpcNw60q+8az77N
1lw3YGidpp1Y6yzHvb+5L+IdrLwm9+XFzsb1N23uQDh0OyPKSYiortT8fO7Psba8dCeYanUJLood
cHzEWzFfYaQymf2SW/Uon6xBkZyZaVrdPhUV5/7uq8+kAigzpv4Tdl5dQ2ugGX+76dj5VgZgcsNi
A4rWkr4/+t/7ykNcH4T7zZ6UWalyz9hvULA937JuQbNJVV2mn6I/Y6upI9WYpFNrhEN69oHR45q9
8qQrfTwIVVTEw0AUhPi7OnzPtnmY+zkT9Z3nchC91yVBAZ/pOfWWDC9iIg81b5HBICudz0rPqAKB
ExcBWPMs71HM8JRdh3YFMzcDwKtEh3sCmdjQbjAzLnsDTEijIM1aZVNyudXaT9DUe0EJkLxVcjTM
CZw9ibVUIZpUWgRoSQwET3iUtMb1GIqoHYGGm/iO3blQodgbKNdh45DthZoUrERI3XsJ7UN85LXk
28iIRoxB9sgnGtPPJPoF1eIb9QnPuQBkrezeM57i4esmy5G56QX4mlo7XbcHpzCuh5x1kVEiP7o1
VO3pw/qXAsul/AjMe5nysYWB8GFc1s09+ZXGvu02u8r0P6N5e0RKgqJ9T7yC1Hlu+TENUihi+VHr
6w2F84kdxf5JxQ9YxGsQflCeUwPDfm26zGbQSWlj0jXYeGihhSjR23vASHpblMutefTJ9h9R8IQP
OglVXkU5uxe8fwUyU/BBGHWndT+6f0wUr3J0Kg76ml9vQQ34GOe1ESwa6A72005AviCJJoPMZxsQ
cntIo6RmanmggBlg38CE+X0SifG5Bou0ygqB2N0zMBh4YF4eNKT+QvLlx7JrtDY9sXTRPXV6fbKM
GmvN1Zy70x/zj0E5LYOa6enTl+ZOMBcV7wYjkLjRmirdW3OU9j5K0VIokhTioNhPmaZbt4SOYLk7
OIjakdsJvhvwK4zD8dpqVOc3hxIgnF0hVND/eG04ZxCHQkIsLRrOZUbksTySRckdC/FhG0WQuJAU
0+TRcGklfd1lpzlQYQZVWn4OLh2DpG4QtYQXsAkNSxWAdsJyUC0IVB0jbHCAEwqdzmXHflnWcN3n
kiP6aEGjy6AlWtXDj7aE5kgxDnu9t5RdHcvo+/2ZxcbmgWiLwAvu5m7dFVX3soffHj+Ak95R95f5
5DpLYlXWH69j4w1TfvEYRq8H4f3M0fD0bCGJwSAviJ21s7gRV8Ynj7k5zO2xqc2ILnFEcu21FdLU
PJc43440cTlx1x32mg3RNX6ApsLRGRKZ2mU+LJ/ZzLkzfhmtAgT5tBOQ98JV4fZg1CyAauw5hdJQ
9kJyZu+871iCAyCodYO1oJ8epI7GgQaxO9qEQjoSy35WU9F+ahJoLWI8kiSHoJ7D6sgwQqk1aOjt
C08pbxDzyOMJpQ2uhz+2obrzproAqhaMe7K2n3hK89P3tg9R0/Y47k9qpqKDoHEooNBR2/Qfpzhl
uBYAHjwsK6AUnnElVsPkIQ5PEAmckh7U9poLyMruy5YHzWqLAx+k4qeeuPf46IT6/1OnGds1zXWz
rG/gA9uRVIl9kAYbGuHf8B3GbptLkSNEN5jG8BdvXZUtdzduYzqdbMtGyCMM67YqetWk41iStkYy
oAE5mVoNYtGNWrxjJEWXCbvYqa9yj6ZsKw5rmtE/a8Y++eQyB8W2/5FKMhXjMYaeIANqaLks900B
46F78pBOO8ZjLD03emeD2HTGTgCYBMmsRsBzOql+X4UaxGPdUWPNAH2zlIL7g+ifAF6lQCW53Cfw
gf6blS64g1nylQNQrffOsbjDM9uqbJHqlmrkyKiKtJ1qc0/78cwPaQeoDQzoaFnX2slK7vi/onYM
w33FiUnC8jLwDgp/Tck5VQFATA/jdjI60Jt5ENG0VognfGlhLAXY4RI0AB9CvtTSjgOR3fQc3DqQ
M227aKKQSmYDBsOe/Yv9BNYRiGb6iYZwh2QviGQB8vCPi+o1WSGwvaMwSY2CDXguQXjckXCXDwPG
XDK4ynVP/gGu0Kyff9Nr4nDW8rwZNMQxrZQx/bN8yPk9JQY1XKMqCz8sNkbf9aJrtOuj4y61NxxZ
GSuikO+/e5JH8xK2R+nAYz76Ji2/8Dh+cqwOaJYVb5wLIr+UD4f6Sh4yMxnsT6R8OBT53SeSRqkW
TZmC3EVwxwyan33Hl0V90jwVLcmlyHP71oKfn1D82Mtnga7ukyNuQdvk/ayXX8ACbDqTyfI6G6AK
/gGtnqrTR4EHfXZA8O9upljFku9mAoRBD4Fg+ukDpq83s58vUfaE4PERsWNMLAbJhSesqVAXmC8f
D3EaDWRGW7Rb8Y/iHE6YQ2wPVBEDlTObroZzRjddLBut3JGXO6TfqRzfEy/b1xmqGKFssKvu81bM
f9nrLyjahifCDLdXp302gYlMFp57y4UpYi24bSZC/5s3r6seqh7+JRvO4UgBcaF+A6T92uttHfkD
80XlvYvqsXDfeJrLfkADzlyN+RM8icrmCjkDU32i46bDnIr3xF11Nr3P8cnGDFj3FrbNt+MEcsJT
Fxbwj0q4y1C3wIPIsst06v4NW4+KlMqZRr8vSALPJ6gQI8xSmUCPX0Iqi/QqGIaHwOIPYorOm+Wq
WW2odI+MdLIhmFiaLv1e9xtXy/uI4IyL5PPZUQVLh9GmfVGURkxgn0m/mMRFE71dI+JttAUpfnZq
kJTwoVafZNLlY88Jb7aJ3u9jjmjg2rMsUy/y8+BuTRL3F8vplqa5IS68970f+MaooH46sGklMQB9
eGkjqt+Fbo4odBMbh6CTvITV/0KHDIcwzmWz7XQ/3wQsr073pMOIh9sk9BCkphxSem2ts3EDjJ9x
iXR00jUNqmaDq5vO+V5QccPZo9pAb1gBropPinN6zn2zZVTeIjDXbQxnyibIUQiRmsiASoMeVBXx
9F3TnBBuTkCyA1bTLntkEhIQQkWU1ZQ9fkGreZrtU8KVEqvNzDmyC4J4fnXTYYO9uJcQXUfcqcLI
GIRrne+THmiv1gCWdTLuhM/t5WkSoqodGUo3HCXVCKFsO878e+PXtYDP/ijIE9URDlXTghUQl3B9
Naeq3UJf7/Xu3qfGwtkNEaod4c1rtTkmgPksu+uSHLy8t4093TRC4BcJ/zEFWoSh4YQQ9oJYRbtC
O5tl4VjJ6gf+EcmSUlHrXzAitTWHdFgTTWUgov1YDuLHibDpnYVcfSrs52V4IGUGJQnsqtbi1Ww1
larGnLGdtQnPrfgtBhOk7HMvpBpJskcB4HEaoyHr96H2vbOGilslaUfZ5mNDOj47CuEkNeeBfYNK
kfZuSRX6fObXMH0jbmHZHvjdkYvGuL4jUu0TpbTYp2kRgmHCTDUFD6XctmVMlPDLQkvcWWftuYHP
m2OLB0d79sqfj8s9zFJ79e3qmM7agQgqi+9OhFeuzO9QcvEarPqDdkMdAI3QmvtwgM+X+qXXbA/e
oq3ozXCx66GUpM/soIWxpVpMZ3zMmqNu8Ffxp6sYZP2vAxsSom+kwrv9RYhkLFQpm7du+Me3aJNH
MCoynubV20LQ26BoZMMeDUuSsMvrBk/c7g9OqMrR7GVBVOmMkv9dzHXN9ZBp1Wh8hgiM3cWkIavi
hOwRd0fqdUhDo884XN4a/0n5UO0wj7GBhK3b0piQ21Enk6jd+CN6lB+7rIfXIv4eOOi76WkM5iCu
0THrZ4bpNqVIoDFVPdHuwE0qEZlmPBf6VHOfh3qfPVAUekkiwwnQkNZWuAZZxE2ZylxCjcE1U79T
6vuSW8f19qlgfloRd9a2MEVWNiAn7q48wdObqBh8ZLlPPjbDsXXRFBzWlQI0LK6sJcY//HDiBqcm
oYM1Bdwo5kVVvNiBirYQdy/YXfJdpnjZWvr2VW9AbJet9dr3KuEbVwgf+NsgbUHP8VxF+4BIARqL
mVFXJdAoa9nOYhoTmINnNCpMs0dzF1I9U4Jgm3jzfRPY4Xi0l3FhtziucJELqjQOciDI9kgAeu+o
s01TUlk5RRq3BU1zqDz4RCepkmpacmfeQzK+WioJc4GFCY7W7HQFOOrH76GR/tMuXPSthOcvzL56
CzmS7Nji9f5elJe82r+1lJmp8QC0ZNhDiNZRwqKoqyaQ+0lBG9+Lm3kuBeTN1cnQMtg4tOfqULCS
yvV2JFYlsYF2yGeBV9VB50ODMOKWQ0P3Y//MVqzWfIixVn97ev4p7A3x2N7bAaJ/4DZVCxzflpfj
aj9oNgNa6+8SwJ6MLe94UH9S0Qdw6QqAo0FW68og9DC+4o3iax10uLG+Yi1slLtdYOUX92f2gDlX
ByM5EsgFhEjrWEiiYPCBQJPoVBeCpKycuiSLogtlcaNRJHaLVjOJXGTzuo7M/1q3jEANlhhOwy04
e8uJUayvhxf1yFnVJQpOtE/b5JVT1jK3/J7bGFx9CSdyq4svwx2bTdJKuWeciqEC1PS4qcP4Th3R
d0nCuXNRACeJYYIbNbjUxfoZ4EREFYrM783fTFrB8nvue+SB3hXpoDetlUxkcm+9uuwZd0t3cLgj
NGDZJQQhkPIbQvV2+OFIUfi1wngK4RKok8uRSOePqrj35/rXYVNCscqu8tRBYIlkQpn8RDngDKz5
lKlwmRQElaVv7PhB9hAJT8K+1gZIfS0TNqlglFEZVXoIi4msxN2L+GreW0wBgsvWB6EMORYm2puf
srazzGTE+5zycWJ/0oDev1l/W/OUbfDDKByT8VOcLAT8m5pTLjcCYJ7hxZ8hpVhs6MpE5JR6ctfH
cVg7h4r2vje8ukUYlZ60yH0Eq9buzKGW9z+BwPoY0tc6lwR0FO9yW1WHuHSWb4Qeindxd/Br16wb
UUD23tr1NDx3eSmbeyhGTJI8tR/x/qMra147UdN3fNO6l7dpVVcPeQIVM91KUdlNh+mJvNY4Oy7l
b3sL6/DQCy0qD+/BmGveMsiQh4LFYQXjPeGlJ5fPxsrIj2QtaYskc6PEiz8LEbJ6iYxAgvDlvb1r
bZkYSkhqBuXjb//GzBk3toYYQCQ9n1GYYyijyhYqK8sTcCJPMSbUW9Xh2YbiymOD7DdPG/Gn4kn8
jrbJggMc6bysNVySlto3S34wWQuCl75bly2nqudTWpFl9kS68lhJ+0GvdFWjtSlFdd07A0SDNFdU
aTG6S3UbqUyLXsP5Mr6aUvY3Ne6M+xI4vQ1u+eoxUqmWAMCByrhPqVtIyy5EkRwLlkVQOpiMduLi
NixlGYhtMf8Vhk6hXQrReNqoG/eEhI4wRgHZOju+fExG/CTlaSLUTCCcJyqz/rXpUHyba914MhI+
34ObhivtVRRC/std6QnXWzc2xw66iK5CBuIE1ERyQ/V6NGjz6TpK1D4Y+1yE2HG7/5J04MAeOJv+
BqFlmA0NZC5jYZh39K+/IN6xcrQjcoGx0tNAzd1GRSjkf7ePCFj9BGHU+g7VczUbRu+QWSDTn1f9
x0ouP0OB9A+MZ0DpS5eBDIgzWB2hrxpsxzQOldepsNMIyNJLn5TJdD1bdybuHtSvKZF6j4VCkuht
VltBib+Hr3sxSDlN5mWLzC15iOrmASCBdOdqlZNUv0o8/3N0pfpjk7j8RIwuh8CFss29e+OSNtQN
gYa/H6SjFGrfX1btEjuY2TILJAKPqcZlcbzKR+fTa/pW0ecexAGEZX9l9sBQj2FKSKD4TANEfYK8
EEyo8VZ/gySnjdERTCVY9B7E84TXEqaos2sDOmCY2eBVHlSzacnqqSVi5hCvHGHI12+F1xm2wC6N
DkhsF/+O7XlWi+IdxNmJPIHntM/DghugEglMkC2zjHlQptePJQqlo3uPrxolPGODiHuryuXcA96j
WNroE1P9rCyRWwmOHG/J/f2Bd2MYqTYda4v5jT8ga3PGIeD4Pb2gYvB1xWfAjkkmNESJBoq1yWMY
QB0Xvp75LzUJbCutkgGFVXWyi08uwm9ENQNNGghh6qSYkzrcxFftddTAnMEwLe7uIkmSFDcHhhyW
n90YIA+d3DgxbK4fhL1SIZQLkLC4WVumJz6pj9tJ8X2NTX82ujLJSCOQ2PVUekGO19cUR+PyNKz9
DmNvhWj+qKx0liPjQOP8ys25cmy57+hruBhnkDGusFJp1uLHnap2MAonNQhF9ZuSsKnaxD52RDVz
sww9EPdS8VuqgWSbxk4GSmeqS19AKXcH1ZNA3eCEJDqStG5WgjTZgb7JWgcge03zRCJiMW1l2Zau
mxtwMo7R3Q4o18exNKH9R7oDM5Djo4jK4C3OLjn5jp5v32qqfYfAVMcislkI+zWFZ/My8xaELDQe
+bUud/xCktFw0Ug7lVzWii0PKqlEJaL/6HNdiLFhdendgHY9vzVRdtxLMv+0gevcU/q72M/6WMBA
OX/TKRZRS+1fXwS4Ak45uTUY+0sZO0JBGoeSz1qqH4R28ZrnpdtOAaGcq28DxW9xsiD1R8HqoMMW
PUjSAAFPMPmh/yFdk10StMvfyUVxLsRsd4i/WmlUwkd3KvJ7RjoSD87hgAGDLDAD39ZNduj3iVdZ
yOXgkTtNskSm0FOg8+H88eiIZyb186AA1wivb/2B1BFDMCB2gEnMZ/K8bC+W7wUAoeB3AiBNvK13
YM1jq46d+mEY6ms0hPzJamtvFUQpxehtJ9RZsJ0vWHtg9s34qP5k803ylZ/NEl+Sqr8RxMZsSWoS
jokw0t44bT/uLKIx5ENiDh4lwNMpQ6IIK5c3OW06XhQODi8FztsJihT2SAfWfPe19VRX0bpGfCrF
OupbNDfVS+Kf202tR39WPVJhFCGuqwFlYHYozN4fPh2/OsEREMWNV211oaJM+w4qXKSA79QCahOp
OniTX7ytGcZCqppHj+eLm3A0XfK9/TYFqdh+Kea5QdFM01RHm6SnulT6pdElDa1ZRJAkNEi2/ObP
xDWdwCzggYMuRq1RfgEiw+m+3yI5Icd17JjX+4G0qT6+jYQvME7j21nIwC5/HO1vRzIu+Xce0nyv
NeUhPHABpCP1DhHK1ymlaetq0FsPnzNWp0B2vDyFbKX9zFLkecszvpejleE2PHLMP60i3oV/jW7q
bOSYppo5Iy7iY0yOzMGBsjydtvzIyAaYNrIJU59LANt1xjjD11E4GB2MD72Sl/ORViuz1qoRwkqM
mU3TYwPCiLeS1hxpgnGLpbeLn2fw2zu/1eHOjU7OCzhCN9+nIQVFoIK0wTZA8C/CFV6yO0SUUN+Z
+8PlNtTb2pTr2N4uXlk+7f5XaoT1BVpgMv/pKATZyJwW2s7wd2AhMDThYkVXNQOeHwz0M8zt+NpP
pC69TQLTJjctlDnJbIRFSjj53k74Y10duE8xCwa7OcsL9avZVaFJAD5sT7bwOlgVAjql3Fi2U496
cXPuvz2vNYCa4KFDDtn12MHNdRNH07uNMR9O5h6W3809nVMpYlV0kiYBawy805Q4LmhVpQLfV9cI
+2vivZz3mNlJR590vNGNDF4v05lM+L4g+rege76L714jKREk3wWdb3BWT8pDuLGmXyNKptQZDdQx
SNDe0yCoZvtqYIs6J70cABWKv7tuZPJucyb1QC1VFs7H+iONRFz+94iVr1AFM7EdtKc1iGyT3x+F
h361MG1DEOtKEK1WfqlaGQJ/01ibcx2qdntedEAIngGhdaHGo6X8OaHChPvy+CQGEbgc/tTI5KI1
6eIMq6+B0nudhY8tVP2jMKDv8Tf3IoHmtgxtQQYsYtg8ebh1bfo4O0rBO24F62zfeMH/v4nG4Mm1
ZiLJ7A2dW4mcrKkTpNVzHFGmjIoyc0b8+LsTKvSRKItgoae5cRIgSGd5jsbjlu7NB65ECNfuehom
KxLoGsHdO12oKUS8yiOrVhkTBIEaJqlhtx6arDnZ7CcycsEh7X0qaXEIhDxbneq7Jwti5g5sMGmq
oLEz5yYovL9IjnLuy521G79tm8r+neWhFJAmaq/rYYtvwg2TvMzRQn47IrGghZDZuf0EjbEjHPGk
rVOcjuPI8Yl4H8I08uDNLLyIsZiGIR77OaZBAWHk87oteMkpjJrHHbQxmYsDbcTHPNUkS+jN7u4J
NzRyqhZvePrHJZ5/q29rdhknBBw9O7xIkOXhJiO9nvzOYbjdb1qPdPiC5E6bm4TJIhj/mKq7F86H
/iOJReG39ob+dEtG9OOhFuDXc3XoDfT0/eVwJEatNxeZ4s1D/weNp25WYbOIlEr0+H1UdQwqMkF/
1pB9MfirqK/ClqW6OG39cye1DlRjtgCc0Bbz036y2q8Y2OWGEGmxx3V7j5x119Ns3vmtL+UE3nwk
hJthcK0/M2TqyvHgL9zPBhiuEYAulB9nxQoNlUXuKYNG0QRvpBOjqv7xZY9+XukfzydiyV2ofMwC
Gnxv5Zui3sWaMdNa/QE6GkABIswpSouSN4wVW8i1De93Gy7KmwUpVa0eaK3UDF7yJA97IJqNkzuu
y5CjL4or9v+LUcBTlVEGGhQBke1RVw0z3MJBwBnfVchttsgeJ0NHUGViQrvqFahAq6vm5AKTHK+l
AykHI6J1Vlly9QTB2KqKxMzACTIu/Vqf3MVwF/FD/z0MHqh9uUwcMrPCSX2MaNg7RaPv62vravMR
vwR8JFLAvgZvrhsGmG5LZDByJqg1fjiZzIJV1B2r1Tl12uELx+aJlh2LmC8YwkjaZpnFJ1cb/abg
Os19MmDITfqGupE4g3G7dCqK9iIorOighNjut0lBHKzcWTi4NDektuoKyzmVDtM/ZA32synIg6su
BQTLkDUvsibV79yCcYLAumTHbBjGkoD6p64/lwNcIlXo9OoiVVpif1n0D2ffowpjp66hE91M3wJN
ZDDOEuOlETTjqRbNy9UMpKfZ/bLk4P5pVajcTfL+lFXZKa1fYA1CDWM4U1Yk2I9tdrBGMWCAVIFz
/XrZEeTZdjOONmBmBl+VRC6jq5j04ScRFcQRyKjTU+BFfrouwvevvJOaEDE4dwXHU5uHZJFWudku
DYz1OCrpZB6AEVdp31n4KL6T9za0GP/+ugBxqB45wtXsoTLqwfpP3AaI0JSK0saNUX9RQWkrfmmY
PpjtZEOIhPXhbV5/ulk/ibM1NlHTu9TtayhEyBbNRo2/Pkp0hhLG0CnPdxHyhHwCO2PI8oPfdD4o
fpOBR5z2MerB6hh6qIR0B8q5jdnbGYZVnJdyhtpTMFitvF6rGg3RgOWe9Z9go0xA752lW4N2vJjZ
tOJQqpk8z9RC4BnPBYNa5BgUnBuD1yeffc2Z71tlgTXtLdnWuRB3VZLjtd6WYF7AKtVDDJ1lOyHT
g8Os828NrADosl+r06101ZEDL8MNa0cHx18OUjLk5Q8eXaI+4w2E3zCeqyjfnBf0Zfeir8u1xu8C
/ykFqr151GG5adYFiSDIyiAlfF3ZfXE9zJbn4fbVcgtFZRoPtAQS+HHVBlGa0FWRW3qUq0MFTLZ6
PzjT98ntt2AKlEMofJmlu9tmyJ/wbnaf++2HwBoBT8SfWUDWV5QL4fhcvl0s/N/3PLPv9OXVRFt+
tZOmLhgErAvu4DNSckTiUkU5tjQq1l4rwIcBGUatab20xEvej8aSLuWf6/xmo0Mk0tZpbUN+uWdk
UBLcRk3UXDJMHyn0n4PtueyveOkbfnEVUHRL+uOUvWBy0p7JW79XQrsLSrT3EyjOwy2ZIvF+R1m6
8TnLRInUtAc4A1LZXf7CVWiq3kdTOwulr6wHf9pqCDQVLw/tBqWNSZkshKURYUSVCaQodbW9yoX9
tYpiG8HwtdBEX8wzEfVMRnRRadGwsP+8a3K4goqlKr4ZlpCXk0UOgwAjmTAbfFJksTqLXKOEask4
ia1db++HixE2H8uNM7ImVW5dH6r7PVAloy4SYHUKq5K6Ub5pprqmBBQGLLgX6iE3jHaG1eswJahs
Lt0HrO6xBWO4NtqRzZl0nb9U52XUEq+TqDwv1hsYcOj+hQEgQWboSjRsRvrLHLDSzeaqNvuerStN
bDiXZDu5XZ5YdzLqJla9I/i2OzNbN5r5FSGH44cO1AvV2j2ixPGwrW2Oe/hwb9NKeL9w3LmEUa2p
TW+qce0j/YH0XUDR+hIIob1FYh+0kbI+rsuX+kGuUNdnzReg4XiV/j2pTW+5rbszzbSBPpu7VEXF
gdBMR8fXz1jMJagfgCzVdGhnF0ckgFCqD4V1gfv85iyPPb2LQDhgWHQ8dEVpvpg4sRTJ/q1LVNFP
CDCIQf13kTFZJDvKyTXIYGPj+aM8EIeNEGyQmc42x8hhIFXgQFGFiw72pidn8yimbwX/PLqrxjqn
Gqii1BiadoIonaYRa9axrbkc8aprI6yWNKY48JL6mvaBTbgN1+lqkt/QNx5NSRVCM1nYzAqaTBN+
EACwVF+/pGA5br3bimYZN7vq9zEWiMk64rkNGFy7LZYZG97x+wpjw4I3gyLWUSy63RAYu9oKBDpF
7xwuV7w3QdZnLqOYNcP0Cq+/OxqgPgz2AjulcHbZ5kVUZXuL6UG7jdIOc2999kIY8Gf60VAZaj/O
psL342vHq4OtSbQmjqtmKjdJWAogkt3Jhkb0vNAshMpLLXuHwL+Se7gsbO//c+tCqXa9kXwqlo50
avFcyxXIskdhoHWXVe1DbBjO08W8Rueh75vtqYY62OU+T8yVEktsDBIWxovBSLzQ8IkaaA4QcGXH
x8tSounCBP6WE9wj6rbLes5mdEEBJDnhF3nFHiR2Errp5LTJaTYhgTVY9AA4wRXbCghSeJktBgpG
WPBRsWh32vJc5vSsH9bL5rHOkl5gMEBRQDlHxctpdsUeiTkRwglynYvUQMRp9/RYlLMCs37gjuci
EU6hh04Nj6Wl0RRuYhrF5cGHus4FK95T4ArXvVjGkJ1+R2tG5a/0l5Cc1nzcbbhQBTwNP+DIMSfU
VlYrTzESYCFC8hJde12q0an2MaJYl+UMQ6jNMVvU3uvYtXiSBTJ+gb2PD6vgdn2b5q0TVoyh/Z9w
J2rc2o+/Dl4/91t3i9twq8rQ5/TSnovXOZPjPnGwOFQ+3Q6AOO1PHaOfTsymkdCsdR8Kwbxs9L/i
TxCQwQEZBccrwVMF7YRZ4G0cB4x2TJvU+CJxwC+KqdU1VMwBdnAZ3PmN+9c5Z599fbhHckZPLKnJ
oOi2lFsYbSX0OiCJ4h2WbdTgLTWW148VX1sh3SCI3OwlvWVbLOg6hrq6ZkCPslf+ZwXMVkUhzg/P
sf8zl9yyRGDS06ejRT35SA+cdUiUaTftNhOi5hyVYQnNGtVIcbu4f1epjsnk47q/E838H9TOYYMi
W7e1KBzhDRovi46aM6A32nJK2eEOi1RCUvhRUV5A+hrpDe1rnCQ+QNSPGqJRueEKJbnCo/XH5OX8
RixGPNIDY880WpvcMJZo2Coav4r20SOjfhSoAItS9X24r1kV1LZ/aPYVvQMKoN0SjnjKekiNi1VZ
nqU0WOF5E6tXmVoUi4JpITm/o95OJuH/1u7iGpNhyLe82MVZkMlAqTHRGlp520aoX1yYSkqz0DB6
1D5wI+YCj1m0bHaxcHgawEDl5xE3qejDLrx9GAAsJJheYSPoYpyg2tF9PgRJc+WbtXb1oJPIXO8/
/KvOhEodca1p9d8bB/xgtwQgztAgfvpM+GPX33TRrs7lo7bgQKJVGtGo0VFdZ0XOc/7urhpTSQpi
Udk8NqpjPuYrgK1LiAVj89/tG3dShT2o4b/34xs4tLhXQCbJA6LTDAwaS2EZ8t4rl0a1FMop1aF2
CkCJsbtlbHDEP3D/2CWxSCEwCfQ3gL6zMkuc3UEe8N3ctsns1EhV8GV/v0qbljtgs8gleGBn6/94
NCvuX0yVJMur/qxwSd2l63+UxKW7DYvb+kHH7xe3gezsIysYSp7wz9Ic7QXzqCAFKStia0T+waPm
+sJ7Gd/jpWvPE/3Yk9iCgnsxrK1pNqEMCA4CQ19kOpSgpMEjY5pzuGTnOTkVZADcSf/4uJVBs7fl
hMBGwuZOxxNlK9RkIoY3KX6xVIqgQjwSZ+Le9QZQGLzDwK0lozfNpo6KsEhKORmKOiY+vU3rjxNY
hz1RAnLEvAs0kqg8md0bOGs7vCclntXlWziF84r3FHW0VpzKFrLHD7p78f8SAOVu/bCXMavdtWi0
KF9lTMK0gk64FKSJZsCdESowI0ff2WNDdcx7+PQTheUgERuxFmkvm7iEY8Jgor/kPVuDl3wtnATq
6VXL7rtXpwWy4gPh3Jlrfuvp0RlDXAZiecUORYgUGo4Kqs4wurvb0j5u6stJl/BLc0gzbqi0RwsY
2eg8ZVk3n8IjoC6KH2OjIZLAzInnH9IrkAfUIBp1SkwG7RlDiUHoUAa9cThza+KmBngc6PQ3ULsq
c9qMRXMaNb+q7ZEW4onrNAPVfFeY2Di/V6v8O+wxAka5NBRhQQQpy6JcOVNbJCAbdalDroE2Tm3z
yLOrohB4+BpLtRXSmOLnHpYSyLitLHcWEEDny8D9RI9d14ArKLWym9ln6te1QsTZTXCdcjmYOOCD
/EoAOmTwa3n8D3Toljd8uPO4NgRfrKqrVlwYvsagL8cOtQm4P7Yar7HXlwiqmZSdBrGGb2ba+wYA
1oM+Aas6oWm85fHeRIZJGJAorYdbqU+Fl+m0DcwV12hTrFVaH2nOlg1WhJGzVJwvsJlCQ6Q8SHeR
FYetb7Eu510iGBCBBvhvYPl1dtlpw9zQ2Tp3kaljhMsNRO3gRd+5qnXWr1ivn3dJ4bt5iC/nOjrI
z15PaHo0AIEBUmgKgsn4rtRCd1CPvzg2fwj9FqIsE5tfGEQ7gqqKufmY7PKHOxeQ1KdNMxGr/njq
zszT6Mb+Lbo82tznA0uXlN8suqTONckmYKcQWU1V2N0AO2NgEoerH/JIhlEEGPrgeJIHH1kSP/nO
/KNLjVmIpOreo0WKaRa+7pNVPUHHI3kt4iq1t7vOMoEqYRMfdF9RGFvYVfOoTbVRbOdFoeA8RG2h
sAcw0b9qieYk1B0jr0lqy2ko1zrPIJvZy3gUvylw1A23jdRN2YeXGSpigEt2YPzlIxO0aeSQiugq
/GV760pcHsOPdNyOHQFvujXtH84dcWackzX/ucXgoqIJxUbFFLGMBd3+Ai9hA+tG8kAwdYqDcSah
uRALXLN/xU09J111Rjef7FggpKttgVZ9wu5pzs6qAS01ihMuYPkuTrhrIyohjX68P4jux7eLaOhv
ou6MRWI9jjp4vKF5OX73tMZI6BYuwV9Q3VAhY3IMefF4dwaChbnJTko+DLQ6VNkXD+w7ATzytwjB
OXo8YqXJcp3EGUHubobIkahnvvc9lp2zrb5UtbpJ427SC7o2GAE8tiPrQvfmwf1pd7Bz1d+imghh
WUqX3wYfhF8v7Dx7f+nkyHN8ZGEg40vuBscBAHxErnPFqUEkxGultgQ6T2511NzDleOzY455kz8L
zTJf6/Z0DC4G188xpu/L9KIjMhKKfq9fJoa7pRANjUvrqx0tkpxai7CHDClERJZ6IL5eX6PwB6s4
36O0ASLFgptL1W9pgKkqGmdMV1DC22BEdyL2vZV4pOW/Dz1qQyVJu9OTKtUOer9P+76/CwLT1nXt
FwmAXPPRWGjMQv/e4PllNpsbMjdZU+zjr/0zWJeS1CWxKUQRRDUVbqVtx72waz1FXhN6gOJj3Boj
BmqTgEmafE7Tr7xL1WOO5cuZ+7FCgug388RZdaTxO6SljlPjba9x6Lw4BMV4xOcM/LUobHvfV3w7
ZCWAkweTp+zrdvgTmKlyJXgszDmNEcHGedSlN97Kq1UM/dcGXiXMJzJwlB7sHrc4ubO4PMOUoWWv
qhKxATQliTSK6YnJ7YNSTLtrKd40Cj8/1YdBNH30xx4aVnJnY1rr3ZOTQCPOKkkVZV9FCsOqOaQA
xoJE/8UI67W2gM3EiyJJ+a2eznUfwHOhjIg4wHqZwtBOnBL/GTogxD8mi5QC8pcgxMurxG1bKxTn
k9CwooW+j7R8syz75Si3Osl2JTA+cZ0DJczRCExdEjg+OBi/tRF7Rfrh72bPgluvKfllYrW5V5s7
MjBysjJyQ1y3FnKZQv4n3bonWDL+mJGObLi3iQ93z1x0BByhFoiuw6mbwEStfcLmrX4FLSoedPGd
XmtUTnttH5u/4LOVbjk09veHsEXd4LSiDxM5+PgWEZGUoxM2dRFxlKOJRFSk/3/CRVyBV6coJ9u0
uCt6Mftt/67j9iIGogHdPk9UQKUpE3XdZaoShGD9gAI+J4y8NE9dv+1hH5XMELWhmO4Mo5uZg8n/
VKmNxZrwtsg//HEaq5snhWwHKwwQcHYYwvUp1geW2bs8CW0Nr1+3nqiymEJkKU2r6zjRGkl3CccZ
JEkyo+UVJjPhaVBGsCbxvUPvlvm3ld3XbxR1iFy86mPGZI++lEQ+OwOrWcGE1aYoozAi8vlQkq0e
uRFAgE0JYoOdUBx5nzplWiurXKmTTNuir6Zim8WLR6ccTDppkTkkmM6PKrFT46LWQIGwys0AGGxz
fW0Jc/jg8JnBF3JSwGktyzpbvu7jy11bFHQlFD/wHHoyPhlWn2+v7eybtNODIqo4HvNpz2eLyIbh
9oMxLajAvxbYsRqA7kuxzoD8U/Y0sSrorJFlA/+3tqPRZRguXILTS8vdmYtUKL1vrfd2/yZiwbme
japJsdCUHVz62y0E5ZXCGp1Ii2gpOa3E3+Wv2zsrjIvEdGXFgGtr4EpWP/mTNOr5yCRtb363CnkQ
dR04m1FoZfvimfKYajgiCio1giP+dh0wtlBxG8CHVyg1SeE4ssDDbmK11aaIydg4KOzkYc0FZK4i
DSV77Jq/qglF7lhdh4ElNmjxrMHfoeUotNvBbkD/2js+fLy+dUp46c5PRVCoA5+LIQu71ET6PTO8
hw4U2SNW68xh7HdspDmgC5gqenljC24Gb0jnaxaIiBtAR9QLKNsIbVPOuIZRIrx0F6l1h+n7L7ia
4vUjfhstSn+lKoARY78vaRBHzIZirx1woN/g8Lz7sN88u6GaBB3XC7MxkfWk4AUkVN5+XjDVuX6h
bgEPSR9kiWO5QNq1pa/eY42ggchZStlizP/5UKxB50UGWZy5Q+7vsUGPeyFO4DabYwAzXRJ8pN22
xgWh9zxTgZX+avMf4MmC+EZGyI+ateypB3EqGDlcu6RygFVNXcBGKUytbULimFHlG3AlhiyrRNnG
s9QVedTU0WcR4y4SxKJfSLgEY+7W29WxRjvrs1+KIb5TsY0j7Jd3A5n6nvPItSNbuhXvNYkSlQ0f
xXZlE+4wupo4qy6wbTSc/RXLidGCc7AGFV14EO+O+57O4MXQGWxxB45FPaSEGg0v8KlwKsRJcW/q
gOYJgFIgnRX21VHZcZBUrAVInpuN2QSKjPBTcOWEJe45eP/M06dOjPoFeb0Uf1umTIX3QkgQEv7i
gBv8dU0ImGiHwKnHWMiqYeEWmFD0PlCRtB/cxdDBDAZbUj2SH5/WuX2IBLs74MnRcuUgQm3XafRD
HMYa7F3OLH4g7YOpNW5zRtue4RCAQVwhwq5FocC+9iIxo4WDyT6HprfE0JeylzGGAxxhiEiGNL2Q
9TVkOgE1P7NBF65R1+VncCXLnXTt67JnzTv2HzjT3FPf0p5NuP9kebm7V/H6zbGiXWNitkdzcZkO
I3qzaE8aRytZF7H2bsyYTKCLDA7/we0hN7XhUu7At7zFI/3bhUv30j8Atylp0PgzXaPmsUt09Q26
Ddn4kVruCO6nMTJRlh9VokqZWPMKbdym/GUwDIeh0dmr6CIB2rJHcevYnjhBnHoA/Y5geCUltDGq
4h9g4xpR/34sJZHoo0NH/ZD+5KlawFIDirXuCtW9RoyIIXt7lEbLEg32e1yXfXpYFZWANGY8ZQdx
+RWbaok6lhmcgcCjgkXnwo1IaMe1cK8tu9Khs0MubVz3lQLRGZagnnXHNb6FwMYoyX/ltwgczRZk
Osd4sPWDGt/4BSTYFybzB0jPL/bhvRoFw9XQAcwZI/pSBYHHP4VYE/QnRYNTLBW2BnlAGb7w0ALR
vF/406X+fTDeR3/ZJHs4hZ7mnxuEyCK3Bc/GN4wX6iRLz6Xahz7M5f3YGNEJUqjOBdLXlun5S0Rd
0M3NMieQ30uWou4yraRGYQ6XZLcFmVG08eIl1ZmHSUWl9rgefaZm418so2N1eKj1TOZdqbKgmC98
gamEpjGDa0dQlHPc7dDPju9dihZldNS/cetGMJskQUV4iJRytaQFuxraNxtxA+yLk8u8say1QR1W
kAC3hhKg1vuIz2gd6DRBjrqA+U8DBjIiOa3KFtSW9rMpN6L1K3jvP/ZEcyk0p6rOms7wUdpQna1f
2+K7v2fN70UKzj/aezqqH3IzvnG4fGShZUpw40X5Q6aUMe4ijQGiD7xEyGuxPubyFZmDci44I12c
w4b+ekWEZ7GYQ5qib5DscyXPg4ohZl2aamEWsnYBYg4PIZBmy6QX4yBkkyuPNp4bKted5JzVpau9
wzkm7Xo/Curk/6j7GF1M6+9r2nlbyTiMcoxOSRsxgl9uUb8fb4TmDqOiCrGHARWuB3HPtkLyPo2H
C1UfDK8oE4LHvi1tyKJFy+Y8Z1N71CFPq+f3/i74c7K3MhEgMhwutuhKx+psZg4d871wCs351nOj
VRSksXhcr4ilaN3QaCV0mMwipHRmNNGUPFFaQ4n6jbQIrVGZn9ccf3FEVwnzZ3dYvakFCXIutCgH
TqPKBDn8mRy5baMQJFou8NJGlbIgsQK4Sny+Lr5KGfYg5aG7+0kLnurXOdtXzclMk8ZqqOqrbIxz
i5lkGsjR1yHM49CdkGXTFvWX3tOV2fAhudYBbE2mfapYZfFV4cIEcribnx1MUtpULIx0yRK1o1Lk
NZdKXaK/gW6AKBXVSAUYZwgcRrZrcMjCK103lYROZP85NYh56wwS9edl+utypN25gzXF1fDK0mAM
/guMURFKmz4te4xji5fdfYKJiWrclhetOm5vzyG+UzGPbNNiYUAJX09mabnJDbKp51he6/ayBkkt
QPFSHvo2tqCLR/zSVKzNXuAVkkkkn0Ki/ARKrTlYxkAhS9Mp/+fo0Ca2neXFFfmaksZ/Du1QqsDa
yBWJM0RZWi7ninfaw4RwyiNJmCuHkZME/0sztRImDsb/RA1PBI1OMecRibLmAy5ePUFPNHXmAJPF
jp9EZYgSfbm+Y4Yw7rfbsQywYrmRp3XvG56donyemXF9gbGeuV2TTltn8IUblBtMiGLGlu1SeaIk
5s2aNVYMhrsqGdRIKV6WrlvSE1ifswlpF4Ermgy8WAdaFR9FJettt8T2wPn5xzx1+BAScEfAYEWV
LiiufB1jfow94WX1UHzIDX3YNtbDdSpO6+LX1b6aBAvAihUujAHUa9eXsa4zIREpg4lKZSI3yOvG
c8flQAPYf+P8KY8VLE4X+XJX/xNvLf5pfLHoSSRVVfj2AK2yWXO4Tmf19g5XBl25JMvCvg/BpAnH
lQ5/wvu7XG2COy+mx5KbUtxZLmTZg/frPDIutsXI9lhrLuwtyT+mUQoiDP+OPYt+lAAHOyMZTvaG
9DS7FPnhp7/9/HgQBjqdD3RTS22SQKu4fsgy1+OUxrpe4ofKuZEM5xHRf8DYsU/lfWRJgzu5SjQ2
ju+trl1YOIMXy7PK85FCc49MKtNyCF2dQkq4mm9zFwlpooJaqmaRb9OrcA8RBmWdzNrES8qEX5TJ
2XHtMJLvrrxH6QEOrYfB5LWsCa9Fpkm+B1uqgXqDmXYWaaS8zQPrlASO944TgWMSpnjwt+kBrnwP
A75pSWYi10AAfhYf6przsDR8X5NRv7A6sXL6me98sgRlt+PDASbtupiF7ONsUJjkG4iX3H62+A/H
ZkVezRtXSSfoWlvJZDF/KImOTu9pR7T7Uupo7hqB4cQXMgRg1BYLkhcu+YU5APECQGsH0iKgmfJl
HJ3UhSu9jsmAHS6e9lMTp6r+SA65Qx6JL3Ota6zSqup7ym6mcbHzAroOS9ifZ6ZFPyPsd818/d5E
Jot0ctjIZ31j3fnTjL7VPFJmEeeGU6AyO0dTxi+/j+zA5RfawkPBn4ZVpdTXHUQ2e6u24MWH44MR
rKJgzKs6MCBTzoQuWJJxgMtkuxidRBsNRSziyJdtjXMl4bQ/fdXjP3k5UL5rFFuRhnA8BLnKwbjS
UeIG+oZzfHpsIaRmVRs84B1XxsR9tRFdu7q/ZXPSZzQEeRm5MpZc5H6XUTzhunPQetnlM0GoDeIe
1J1spWBU4cNNJngz3xc5E47uNGErAtftSILiUmPceR9I8ZP7hVR700oeJCV1rn5GtVjgokc9ml9x
gLJARKTxGcedIx28lhCiX0XKSTResLJgX7/S1fzlbQGpRvqEp3bC+5qBjbl0UpBiVP7wNbq9FNp3
ZWaWgQ2QJ4vorMGJ8j18+giozVVzrFAO8FvcsyZ+gsa5m0g5WwvOtvC3FRL7RDz/daYdOqwgTwx7
aialBj8ateqvhmjua4AcfVVhN4oRVGjEuIujfTDRY3r9Q8tlK/mQGh7XijfbdIk0Y0wFmAHP/cfR
0bWRyAwcTuDcb/y41jgo/vGcRtOKUSTqn3f80q6X3232DG8ouhwxK7v19EBVLlvK6FS15TfcC3pm
2ABI7nFb3J8NWcXowIGfDHUkGTwcKIP9mkwQGwDEZ3vvQ1fqCeScX/gpJ+yjob/PVuVWlbOTzhgu
CrHWKV2t0r55LveDc9dAa9Ok5XKYsX8OPDCA8nJobhYiUAoqrvnzd2qk91JAWDslIu6fVU+4ARU+
krq0aPZPXs8945p7NQ7qeu4Mx8yykX5OuaZdCLZJabW9ot10mPP1X7vHGK2g2JIqtK3CUf7V4mKy
iSKdRk6PM9HgaXDFa4quMpE3fz2sNxaubPrCmN/Gv+9Njcepat5THzzFDPCZRgL1CuEDv73TbK6E
D7bsn3Q84zrmM26xh8s+ZV4x+jC1TGZXbvE1rJvOl2FTm8PsYt/wqqYk+ulol0BgEIjb4j6iprZ6
CAZSdfyuyaYRhVYN2tpe8JBf4+Mq9ZanCYb+l6dfOWyreykngaa8KUg1wgUoM8uKg3XhMebObgWh
aayjIST9Sk1bOqXkXm/zaLPu1LPTA2sd4bbQtdno8Y3acKjmFADrlOjjJPqQgYxhRCJL15GAS/71
eiPi3cMc9Iq/bnalnlapI1G03YJZWiZeUMor0hvAEr6rW2bFg8gwsMbLrj02tEKvvY9DjwI3yuFK
n4xYfJwlwI7ItKU5pGdoA7jv+dAeJkFZWt3umSabdvZCya4aVDgLHH+80IpEJMh96lBMB12GNRGM
pcHXDqRNNylXfQGNO2i/oaQCu9W8iZnnWaad3wX/JJizVGClPfkvLJ5yyfuM1+38P+AeSCZgZW8D
6hfQKqbHELSJ7oBXGCwFLE0W/Bmh4sk8I85sw2jtRzn64T7SIvxsGfSVszhSrUO3R8D7DjNxInK/
/p3dFKp6ev/Qd9IYCLj7mosZXxBnECDHxKLsLrzQ8BFeKF/TLT0wUz3UQxNuRKPv/2wOSl5tzZCK
BZsyqgPziBR0DEDhskKSCAn1p+3bTT0LfhvSmLabf/GPJPYpAcOC/nlJHb/dtHOmC3NMu61XLr+O
ielIZscc0WOvNbstlV8HvN5XvVGbpD46bnFCc1vGNLHW+hLUufw6LikfQfhSVerABdagF8YEhirb
hF9PN0KLRLvUduO73AsUd3vCzzskS+YufZTgonNBbtAugtwyJWWXJsOVpu+xQTOFOdx2QMQKiHCR
b/hmqkepGtOR+5LmZ9JeWO09rRec8ygBUElRUlbIaDjbuGftbMvWEwUy8nLPmKAixhukojN951Hd
/5jDswoJkAt48zxrDK881gwZ6O3tls9DbCcwRm503jNFQWeQiPJsaoiuJ7VLqLJ+G9gB3dxp2Yih
mNDnLnz1kwaWf3Tr7IXUDnwVeSK21HIXKjFoxutqDzXw3EmQOSK5gM3eRR2ypjnkX+n5N4ZLTrSL
PAmcx59eCkjrIEQ2vaj+zTSH7550wwG+S120M1uKU49vGbG3HBQIr6Y8WsU62FfbhaVhLSlVBAFl
DLiOghq669e+8HTMeCliW0W2BvfI5y51bYuWeoOW683KHFGuZb3zUVZ18lYklrX+9e9annGTuO5i
dK1BOvRTbfGigu3sZyjEvKmhGpPctVUJ9yLx0Ih8HW6oWKqC35eaaKBSodPQ02D8G+EtPCl1fj7R
eUC6oTYmkFOpKIgpQKTe3mIpj4b+T8+KoK0tR06DWc2p/O5vbyPmZxeWbXcUdtsROQ2RRm2+WF0i
BPI9wEI6K7K35VnigV0xsjnqYz3KN/iK1GdO8ilU+25/D1lRt23G05PXZmRdthNTot38TcVFqF/L
rW5Jb1esJsr4+tnJ4lQ9RwqsAQvXksBH6uzICiHpnIuarkbEiH0BUaE1L+mt7RsXrvjYrLNwQKnC
EPa0nIO9TzayS/UISu/rmW5tPz3d851fP/qGs5Kf77FB77KsoA3Nc7HFdUfiR3mXECWivoMrhHiX
/48D+w3RGFtv7ZpYz0GsAq51JXxOIF/Jihvic+8dFpp01Q4TyIUx2tDI1iHo0/X/hskv25i4RaDN
Wcb1fOvaVZVY5v76EDmTh1mCK2xx6ZsaMzI8buAxrEA3IBBT95Pni9qtwi5MFWZN9kgBFpKfGeWY
2jSq38WO4rFY4ghmILK+NJU+YpiM+lS7YwJ0iQY+Tk7bZSXZVfOBTFaeUcfFrYCEkhCZxqlGbOax
8j9uwhFE3czwfIwiRSe2eRkaLvw+ApnN65Cz2VVzZCGHLi7zdz5kpPEAYdLV/J2NK9cqqELdT3AG
BjpHxFnv4AUDTUg3ACsxe2rMih1VJEk6qRQt2YK5v6AannxwhQLnUEDjttAouGJ9Lz6l6A8Vl1WW
J9F5MWe7fxgagN2MGgteZSktC6kM4d6dRiY3h8gEjDN1lD+LgotKVFhpB1SZQWSOdbenxMqlb17m
XdI7VEpP60MY87I2jih/m1t1dg5TLQ1S5RWP/TEs70+Hj3miXkt9nDVSiHDH8/2VMy02U/S+CFEv
6KE+lgwz2QM8hfLhmFh831iSrS9tybnzsuMw8gupSCV/OnPNx0BLtR4iGEfCZqjE1vVSCesG/d/m
seXtenDXgASrhs7dsKlrD9JXi1sO5FxTdMoJs83Mrz7JGY13zzqIWqd+wTFJvWoaAuj6Fmw56Rs8
3yYuKNUyBflZzncZx7BcLNmx/TZMl/jfdYRWmQBOpRzqVSgV8LkCk2mRQDcf9XAWTyn+m5CgzKYJ
n9nuZfY2nq9rNSrCyEC1+VxyCmoOYWIpG8eOWHlWMI40L5QRw0NioTam1FQUYRQiHpBO1W+lDUTF
uz2ILBbS6dh2wX2C0wygXs6Dy9Xa0bG4es+S4Un0m4/r3VuqUqflLjMPBsOwvFNqPLVRR0rbrM5g
okobbzEV2kUE25WT6rIjyvE1z5zYcYEIetW7s9w5jLeD/BqzDV5oNbuirndg7TPwcADflyJnXaIQ
5AaD0tOkzfwspJkSU5REJMAqMw6BQd3B7/CsI621Qc+PDLnIzXc0wJzOLid71ymw5l+BjKUG2zM6
f7hNWGsVBNvRYs16jy7e4sqU80m95D6rVtFJErd2GzOggdKMb73RYiWPIZwS1Pvx2mtAEzzjnzTz
66AuQWhFxVq41i7pyf1dB2uO/CG+Nnf2NnQ2Z3U608C/tmYwBOP3D6E9kkMsvvgtm4B8UXDh35AH
akSnOfSS1Sgo795nnrNkX83GZbkQUUuTmjXtsTQ1gSKNkRjp+1OvShhlGOe1gtXfW6e9+JbI7uax
KfmjeLxiCodf6Rb79bDoI92l8N4CaW32zADbD5hhyQjHCM3Bhh9IIE1OE+50EE0JWj3jLB8qqe2F
r6UO+6Smj2TvJKxFylnUu3pgJHRU6KlwYVq7QNMDOYq1lehYVVWdgKtD2ZT0y3CAwLvA3OQnSe79
RmSeyCjIXrKfJJ2QHcHHh5JfqjLCsT83D43PrMNIe2w2Da5qTop+7JiwnhQI0Nb7GAlwKydWlaZb
996NArRCSGqod4oSXbfaKGrsJ5AChAks3BpweD+ZVsY4S32VNmxYcQtmm4K00mgVFGc2PG669+qi
W+GLhmdnSFFDVfonGGIoCGmAtte24TvUyUOCiIn/O0eqNSm//wiMArVICrx+C+nJOJNSwLgHJSxq
AYz2nhsVPGZtxOP1wXw/JUZTvMj6jb1Xxs2LeQQKOQmc+zj1u6DwRFvRgumx8NbgYzn1OOlIQSot
KcISnLczV1cieU1eoi2UEXi/q+w0NNQgEtO/NVj49GPjBW+0Ap31lC/3mdbC3OqwlUt04o0zheXz
yDpiTxUjMSj0/SZI56URaeZ6r9S2oKxOlDeGHmo/H0KFtVR8J/imrlSbjxHwhtYg+bjM36bOZPcj
bg7zbPhU8wmRf2zqX0U2D7NqWq1GjO9UyOeAwaZ5W9Lds08OV4iZOMwMcjDUGmjYrFqWLAg5xCUG
SZeFgyNvAOoRKVjSjd4iAB+7KVMlM2rTpRG8l5DwRqEPAXs1v7tgSRomxsDB5Ym0mKeWNqB8bFDS
GClvsh8+yoN5PjfQ//6yFhgaBGNIypdm4njI61aLZ00/xx8O4JvjoPyEQTTHJlcy3rp3DPmyXGNz
6h6DKb8CXGbGNhQB6xW9yPoVLXY2AibB2d6rtUgFcip15fQGvU/nNHhu5nvHuSJetIVrWHxzPgNO
r/mqGOkPzNkk1Gd4Z5uphbPYzClIVBjeSD5y9WEiLNaFmPhsgCFKuR10NgI3bGIry6y6Dd4qaegt
xHYOcV0zh7DJLcMZKlxz/h51UxZXpzDkm41tMh+mw5ADnVErb2oitmBP5Z2mae9yXWnTdCmLeDlX
BwmvadzfoHhsOIJSEGExppR2UkUFwsqctvEsXI0KTsHP2fXwUBbtwTe4uxdnDiE6bUdI92d0pXi9
W0iPLUz1p5R6x4S89kK0usAq/e62ewxCxKsG3So8NIyf7wEwxl7Ds3kB35y8cDEUzw/4Jx1ZaPg0
IT2g3SI9ySl4h/K9VnGraat/ltBQHwMysD7xOhd51+wqWMHaW4jLrw2mbfTLcxmH5pb9sukxkYuQ
JcBD2JeJ9z72E4QRQG6OR69JdJfe8Dkjz2v2wXMoBVAvlnrO/D4vARktGoqXc8ZY+/Pz/BtoWUgv
TNU1eXEpy83x5YkMbu/wx9XAqiZVpbH4VAJy/a6I2vwfymPhGtn4FOcrXxfMClqtG69PqCpkUQ3b
W+LVl9tI0dJWY9ylDorGPQmdphhyktjbOfSyOLKd+Y9DwTiUZdEnl3R5SQVZnfexjEOBjrRWUu64
7wXhrQmfgNZHN1IXK2LXIivp93zkYjmSGdSZ/yBRMF9a58YVPCG0c9D3C3t6HZNx5ju7Ink/XkTh
C1UzCUj05CgBhBJpPBq/UarTkZsIr2qdJFmVj7BZEiK/dkvYQjdfzfBZFgggIqCT96Gu6qxdD6Uq
KerovYlZzcw/h+MeYWqAkvv6aBREWMYMHjvEUA1+kQt2bWzZCol0Z19y4AC9eDZv6fLGCLT9x1zq
Fin4b4j+/EzqdDr8095kzBvBcwdpW7mH8XN796wSsAjeeF9Ex0HqZUPCFHtyaOx9+yevmQg9sw9K
EOhIvqqacbWx6XeLk+/ueB8gMmVT/k4iMD2eEwpePjTkBubVRMhh0hZ/WDTzTT2l52afJ1Gge4kz
eg5np2OblZMEeWkuccTHVvkLrLjOTGcRAefxp3cqdkhCC1HI33g5vxe5SpqcObef+BSEfKh21G9j
d8G1riDVVFH25C9zs8DzTxla9TN+TUN4tUgwdtH6escbatO0AjuXWY0O9gYUzwuuosSFaQfKPatn
/JEWMAojvKynAzX+L66N8t8mnwI4OrXzzoDBOV274reKXsqnihCOExcPVsMoBiIh2h5dLOLAizws
X3+Z7eNXjJ2cBh7et3nZiePjsv9JkPfcwl21lXmPcoHJ28e+6/kiL7Srn36Z/fxdy/oCT4aksEwL
VGhU4ll/i+jRDwD0AMOhF4mRMi0LqIVpJMS30N5TVf24xVbuEJROk0l4z2ZKhDaOmehCYPFNOPV4
yc0uGg6mfz/uwHk6qirjeDzrCpU4gb6caPmbtUgzt9RUqs12i+skAAccya5MoZmQU0KJT4Jcs0Nd
etG8v134Y2QsKGX/TOfv/HS77V634rPvfpDYVXWtDO3l/HDBzDy4q4AcSw2A2gIest3zpwtwWah2
Zdx2APVwspPsn7WgihDJDMk4Ni5asqVQMRw6fH5NFedk2nluYB/Vay3cypDJsNrljuXAhOy1qucT
NbQAByS21dI7OKDSSFFu8acdNq3Ou12M8oR0dbkAybLvEP20V+tSbC6EVzVjk+xAEnRkbTGmWYrm
haTkRlKoJM/jA6wjWRoyUbCzrT5NZZg0nYpirQKbWH1M8oa9pmcx5ZYdhaOuLpPuce8gOX1RQifD
zrDCBVchlfVc4Dr9EzvfEYjisJhXr4bpzOE6HTrYcmVUqdjo1pm6DI2+OUkK2smguwubQAFhW6uo
JWRaotTKlaNhbWTPvjIf4eHns1YRftHmQVfqYNZVmhxZaOTbI87S2beejQOUsZMYVQN5RNFWkT/s
LNO3QsQCH4ofcSrVQRhrFJ3Ydvolvf7M/WL6RgY6r/oqQQfGFRZMw8X64Bou7efkf4qSk8wBJ0vu
7IHNgUY3AsYQxlokHjA0EWIkhQZgCCj9lGKT71BobebdhxA/MqQIeZku4nVqL8DdPtvubhs8lNVI
pjmdcgk3F97dUnhNYnC7YdyojVKNjy+a+8FwlbWRZfSZ8wiR1ER+g/gdtGum/JDVyhYZ7eMGtTQ0
RkQKUfDCIBXPYGqn0/NEFb8xjuNaJJussNlUeu48INDoZVCH8X0B3PXtTV5I+EdF0JU3nvEK1nka
RNMCrnDqL7FnX/bSw2vbUeg/oiJIupNUz3QGBbvDSifuKB1FAguUn3h2szh0CFvDGt8pOlff7pxn
vxLgYqthX6zAh1Q2UYEb8wiEsSDTbsVfAvfzNwqmYcafJm8GEWIdw7aP2mDpKUnoTqdV425btVC/
hZ8S31KA7J3LUyLWDizDXZhvYqFQIFZGNLPkPxtb4XpDtmXk8MZq8BqowJOQ7get9JlpVTbmyrIa
NwxeQOyr7lrt6wQ9zJg1aUFjZbtMH/H9Y40xPO0Em7OHXDRZz7+tcOrGGKK8l16PMlRqLFPaWPiN
2+8AKM40UMiRK40HQbWECYxgcygDLjE/omSMszJXZIJg8Dt8CARpeR6M5RDTX73aLyn6qaBaf5i1
XCdVplKxJmUioqqCCCoJtkuSyuN5lYvzJO170FzzdbFL2nHrd+JC2J4gPLUd9tJYMp63ZA79HqzW
LJaityUkSd4YRMGDxJwZ0o4tqol318CjxxpVAVnCpUg7dWCsp67NHbPwohU/NUd+RWOrgbfje5EW
/B95YTqSZJuFHcpT9Iwz8ctxoGq9xER3tm6jaR0hdFTZTkB3F1S/NoeO0bxNGquz+cAd6Q/86v/M
s9uL/vavx1HoqQKAhxwqr2lH9TEF3/Ja/uYSG/dSFCb5SgKG4TMDcQ+URrTtVxdWVhn3Lgr7w/nd
+zvQ7uAZB4P7YKzyWdC6JNUyUAzi62MExP3RVO1xbs8TGD9xB3wnHOmkespzZtAMpwyMTrt1pFRm
L7dekQe6okJHcGxk1a3qcn730hfZAQkVsS1VhF2BbzgeID7OmILPJldONCcSGvy38Vi/7HZbrzWh
NGiNon+Q4bMG76pMw8ywiLXwj+kHk8kpeSuGIZezDIuSeoKhvn+gAvbQ3D2lrT4lWjsIR1rnt7Zw
dCsjw8iW6eTWm5jlzNWymSo2vft6LGdcuk077mCe30Ntl/ZsF5x9P4rtXiR0kNTjfXNfgr5LmfvP
T90Dzw/La+nLOrjCf3nSPohieqqKt0PKepMLYO2WpEWaF9sCbaro6UVuiZYK/CvIdycVxF8YhiU0
VfXhlRiJ9qY+59wzcpZCFNIyKOaW9Wy1hjhUxJYoiUKd/HNR+DeTUpXnx1ucC0SH+pRcZBBbRBIN
HkJcZYAw8wMCnR6bVra6MsN0KScpSBsQDkWVKqcP2WUD6g+JeJUY56BKzZg5aWkRYP0bG1bS4ScC
/5SYxTsgbborN3O2/R/z+bgFTTvA53k7XZkXsT4jArfPigxMDz9oV1Dowl73DxH7N/X/jbMm6aSU
WFkAlvoiwa8Om1oHAHlWa/5troYeBtRoMkOhSRdRN7ab1F2JuhU4ptmWyNnGlkGLW2MicQ/5uQbS
CmuPjMF1Bc/E2dep8Os3hCqXvKMFlCQqboT81awhkmFWPjNdKkbR24VoQtw37J+TNPlJIWK8w0O8
33BK7qP7MxWpRd9c9wUTsBlGAkXY5ThpSFk7kmafXhWUUMrr55n+Fq3yTOUWx03qUKrFxqYxzWG/
7i19RRR8atECKS4s1ZGDOpPIdkNKLB/Hgu/NvvGc+b802NlYITZXyxW5g7cDPTvJIZwQzZuOYLBe
W1omXfQtpU3EHx7GPpv7Qykyx8fmBDYIt2Ht0ihkL2S4Wd6LrQIhiaK/IDcMUKMmcxS4jQY7XCHT
lJGcEc7rVKK8l7ZbgpOtmY66rEnAJYITAdqaioT44gR36Sqa9P6aZv4XufutiFRmhcE0ykRLvwQl
EFWlAqjDejaerV2Mznh6+JGh5viQfNWIxXrdQIdCmi5/J60y/o1B9c/P1mk1UadlsD4FYWJdqhQw
1prd2kZaIegW7foLZNOSoVoVfXL4FJUrM07mikDXqLJFI1jGEzqfWhwYcg8gHymsoDChosnxkNyV
xFbuiAtTAuer2YEvJ49Wpyre4Ute5mvhYr4DJPc2zgGT8Dcsbu3YiKd4dAyKxEG3e+U/s29yB5f1
i7XjLhJ/cvToG0opVUhLisXWqXneUpeJO21/X9j0WPiB8NCRJnPOT5rOwCaoC3L+XUTY4eC2KVmk
CoJ0Prw+b9XaWXuBkmHJNdPCu3YGLpEWLruQoELTSEV4A8apMmwcDXOFljp5PBRlkLSZU0wJy9OL
EOFmOUi+bzbW8MsMY2jjHNsGo/7gb4jYabAWXVEo+zPAQyyt/IVjh6WgeERiGerjqeTMQavGU135
xWTEttCJv3fC052y3jCoDKBIOjmOb2F1vk6I41fkb0xVvPYaIlTg2tvifOUEwgh3+cop0psPfJF8
S0JhibRsPx/oIRcvB7nAQ51vUuhdXsKPpkmkWBkI5P5VNPoECk4J18mJwZKe6zcrDd+0aAWCWB58
tnLZ5ZIU5ZXAUWbToX0eke4n67jyRdaHfpcC1h9+A72HeTYWKVDe4jjt1+9eR0yfpN36hLy1dp/k
+bULxTIg85vbwNYt7ht2ZmYtdWRO02nNt2y9qs9wbmSBo191sjaZMx0yqWVopjCe8cs/UcJ08vla
U9bFrUDEQ8cCycWLO8+trh9ZjXCNV0BSO+0HtOnoulUZBvjUyx6Usz4D6AjbRe1IY2AoBWOwt4lt
tN/kqhUIdE1EOZXipBTnAF6hX53RSjYKYx2ndbK/u/ornOErLjZCmOTTYLAoa/pmIWydixbDAOAM
n7mQd+Hm6Xhe2rfaMI5oIZe2r8WLBTBHN5zJ03Z3rN4eMC9Gbg+XSjwo+CsPaQauiDTmRBHC5gLF
PhhgY4hqBrc9cMzxOMgcZyGFSltogJAzbWr9ues+CZdKdKr1SG6Kau0Z/4Pl0So0i4WJa9zkCmOW
/wZFOPVIg2JXoO8DwWEDuz2ztK2CJtqNojXABekGLCRAawEpprfwZRpXDmd6DH2SM0XhOjexlNOe
dPoOKmcMg6XMCxwnF047IBhNEZimdLv+VF5H2ao3pKAD1kulaUa7C9Z79KPsMMx6I1gbRZnkp/wN
Di/s2eMPJJaxxco9YmJAPYyqHUUQqa7pnxRwaJhRypU5AuMhPxu5jZ8I2UKL6Zb9KxdfRERChdPf
Lc2lGb3gRpn2qC3P9evmZHwLPeqdAtAX6aeATRI/sWx+KvPYTSz/WrgKhCiOPPbypW3tFkMSMvAf
n0hyBL+ZJErlPbCg0orukv7ChOZoNAs5E+hmltoEe4bB2xVNtY8A/LpevjMy1NvFXxwW3C5XEQzE
jnbuiZv+NZQhqDMv7G1w1bwyyjgMrpOkKku/tUVOyV2k5uLx/2ve5hMVj2/KKYXsp+l+zoRP6oN2
4R0hBFYvOuIsnWJR0PuM18XFfPEakxuXXxVYDRSisjvO0A2DRPmvsHAiDcCWtazrKDhppGyOyjBK
q2ks9WDaJ8ukJE1Yjr2T8PstrPLvyOxjjE6DvGHSqwjdIvorTU2EXhzqGwHvWbr7QFR0QPWo/kWd
pOlHpZ4F3kVbp2iRe1YZxSeGRUerdmCngn/xZx4g2dCQTD06nlP78y+yhf/2thFaM8Jx5dFHor4K
bM77RaEpKooADVvkB5a5ZwTlMhLnsPWcFNgkH1xsoPVbe9tHQ7o5OCctKzSX1c7za14WRpNRG5Fk
3rFKZ5IsuilLaS+oTWC/IDfYEi9xohge1qu2aJ3SF4pkw/WSzIPLUmubJCFymcDFMNw6P0yVvKk0
mow1FhG8fsiURlUJdr1kIBHdHQ432VuCTO7MCQjWX2Q+gYVB23IfDdeVgOkbA2qCMe/v8O9ADJ3R
klrTRYNP6/rHuBQ5jgCZt/bIjjjtZMdiSTcfEq8hLHC+Gcgl31xXMTj+m6PvYt4BqOaEEvTYHhJx
zDs3V3wFpaVnitU3eogMi9o3yBqERXCydBk4eaJy0qlAoND1qtGa1PisvA9yyTZmgQ2aaQgNn4Ht
0QnOGRYf9JMJsb5hc49go0yPxsTbGVthY1JJvmVS3tzDo9kKy02sPEEI5r8YdlfU1W7LxDy1+Go0
qjokrGDMe4Id3ELU21idZYx5LkwDEPoI3MBaEnGIspchVkpxZThGY3MIbNlI0sI4u2Vm/1MaV9Jx
/AyHTImlPdbR+6K44BsaehWpLS8BF5wSoFlAZZQmoZx0EWr5+QW024eMTC/uI6H+AOv1wl6/3bI0
UIyZGDtImR53TpfYE1PXOVzNhPZ/59c3m0oHpOf0S3IbKN+dJ95Lz2bZS7Nh2DDXQGAmBx08FU4J
dkzGn4BRQTHeBWLSVE+B/om8qouK+B+C21Kmc77Uql6lljHLO2vJRqSGwxSTFld6V2Q79oMmxJnr
sQlwheOJPL7fddSkqfyTVKJFJL8UbvGqsyKeQcCIfvYNJ8Zmwhho6xpyl/aeVxItskSsfQNNH14f
pn5LWgpg0mH1VQRVx6KYV4Mn+FEHjR4fXSPWb8NHGxXUggWkmo8VcS22aBr4WW4+Q6wymKgRAREW
Z5IAtJubiWPFYB2oKs0JrVdw3O+PXXpYQ4qXpVEqyDBtTNHElPVtEQ4VPWl6qSpndyt6JVsuNO9l
pPcAtURJBU2Sw0pQKdpFPAXDMXblN2JW+4W+JSDdt31oyAh7jzKhLtI9g72Q3S2VnvZNWNsdbCjx
EVzplGTm0cwXZOiVC58ZFQqFK8fWaWYgg9e10zqW+s6MuGMjngQGFw2D5dXqeCRMrGxzydnxDGc7
puZuuBUrSr69WPAAlWiQ6RLG2Uw4JT2dq1Wi5jB0BVTvjEd7nQyXQ/H2r6TMz/PK+fmfIZcBdkv1
XaLNR/dAsg1epjOdVxmXscWn8E5c48+DErmvop/pOI100442y2CF2EK4ImQ2zYCH2YXLxMPYy3mO
FZu9ih8qhndmIj5wZjnRnvhH27QvcEgE9wexEEEtodCJVgqpPQW8CmkiOvtTmXpbZrS0ZSjSdh0w
Pa2K/4LGnskUmfiejOoaIDopWz8fXmQYUgIWtF7YgVbDjPPkGI64SNO+OxAIVLtMYJD8zexAxkE1
Goj8oyTIN/nW4IUZ9nWro5Mu/9hj8MyQLPFADzss3PZxE1Ire3slInHFRveBXD1ys5vtl9MwbkqO
ikcSujZqg1mPvQ9+cvQ5W/Obnib2hm8G6fZ8sV1dIj8JKVWeUN4Iwva6vPTN/9pQp44nAGTO0Vyo
IEbrf4vgctPnjKhQS+xenMkLKCmytv5gBzcJRXh0yS4eXV2tUcnvIJcgerdpawSo1Rdsm5G6wScv
/AqaqsHyg0WgF63V6WxHJh9mnbwP19kPHII0WRUz228FOoC3KVlCrnk0QB7Og+k17BiB6XrKc1Pg
b28VBd0/HA2YYxq+pRQUibp6a6xhYjYhYPCb1eBzFj8EenEb1yFw2g0LXrDDFt5rb6Pdl5n7qFFD
LQ4ab8pq3tLXhFpMM+Ljmmtf85bkvEcEkKOb0akTmyEzv+lxAZm9mYJoXgcpYe2dj2l7f+G5Bc8L
GMbQd7XojFV/ZbcLMj2DkttTKjHWDOFbrEooXCqrk+GUNCAEd1AOAq7vPp0KSrmzfKGtqKLw+QWw
0P4077p1BZC1wAZMW2MLPvUEkG+PRi+Cq48rU0tuk1YIWcrTSqXUumR0mTWwhoxFdxpki+hVXMAN
m92aoJxVYNJmMEnmHHYDSnxjjh/p3uKbD1odKnvJru+L8lrbtleWMWpMTewjycgwkDZ3zZp9gA3H
7UESCclj2CPZ4Fz8L1/RZJXdpZmcFd7HvA8bdcHAzR3/STW6930JY6b+Wi2kBb7bMZJGyK8x78ln
MnKA/SPB7cvVTAD5eONsdk1lH02aghi9D/DJbYD+QGYU9eq5myOXZIoSv4QDEiIB8g5FE/UKBn//
km4Vaf9u/AOk8DkbuainVDXaRpDGFy26VRRuQTUQNW70mRp9+5J4Ga9/x+h+8E5uIg28mz27u5Rb
gOLyJ9sDE8wTF/vAT7asY1O3vZPw0ZuutAV5hMCWV713C+qbyxbywEvOYVDowqCMhuH8RGXlqtQx
n+9Pyg+h+xhMq/Wozy0t/FQ63OnF5ph7uwDwnztU/iT6D1VHU6O/QL3LbFsHy2fkFNvb+H8C5Kr+
HDI0XCVXGxQGKTG0fBbeCnJ+zyuIYaMXa/Y5uc4F8Aa/8mBihX1JUH/RpA0DaIaYPXSoslVbq20o
mXBYAx0HMX4+88xCVN8mHv6dx+lRaHWI5GmbAsE7KVzBM5T+iu+/01LL6LWZ9lN0oc5xJ8Sr/myl
wbUD//SCNMxloRKUzYoczmguf7cyPurpujyX+x5qG1ZTh4tX9pVk1yBdQ/jipt/nkArJ+9TXjWbW
SgpkPK0R469vLGDCgtB2bOTq3p8sV0ZRnNIv8wMWv/P/8+Z1DBTeTolsAyQgOM/to0MOYm+UgmWX
85LERI+vUl3Dt1Pc6EuvDyY8vc4a+FyO2IOFttiCC/KyWTp7bs+dZxOciJ1YbQL7nEav+je/7Sdr
ZltHN1xkbT1D9iQhDOaO9TTWxhSJz3qlHfUYwRJQbmlYE9i2Gu4IsVXlhBPHZZoaXtCuyV8Mz/IF
3BPwEgWyPO0yjukzwmdqJZv/aK9drmdaLfqcZLddnLQI3BsBCD/0fOOmNQ7YdeJrgXR/QKqWwvks
Io5c0N5NuMOCI8ru2SRz+Ex5PIR0sUR418edx8FR8ozsNSAkvyqnJ9ZRKX7eXCvQpk/9wStXqCax
6Fg8EWcNvE/yIpNmoaL452VuueHXB+JqxpWqpR8mjOouhxmv2JtB7c0qYR+zOInRCN1tZN/UhqUa
sLYYwbxExqc1R8Tw3nx3nTYTormf3PPDyLIEPAD/egWBUJYN3tMIqFndSQSltEZWBwmgpBrYUAR1
v40vU0EqaOxRW7y72zNNTWfH1FFP/KUB9T5mvKVgjXn5I/4c9AH8EBULUKH+eAWwZnOL3vhpELxh
9RszFgQSvwkodRnkhV/i77U6stDgVHkJ8NoFqW1WG6B/Bo3j2kMweltpGAnnFvrcS3+PNL7K5BXa
9PUgxs0155U+ENd8kOuovMIbDC0NjGGILBCLaXXXKzH3z0+Mw7yGJvakdNHyzycJDeqVUEI74oO9
llKkz+iEMKyuUSRiSlrXj1952HWQ3u7Z0qQOQqBQo/Arz0jx+lNpZkMjMD+fng2V/FTpnPXvPHfJ
keaRFi29YWBF4Ft1SfMy1NUsUFF0kgp7C7+WoMnU1tBYvzjsy9bK6R7cslBtkOBkhPPla8/7mlO6
zCqFYz3aF+xmC+4KbNUVWe4kij5NtQ0tJjsz9xpBatQNHJ0moOcEaSq+UM/RACYz4aIA0fCwfpzb
WUIpHXcVGOcY1oRBkEN7djPXnYpZLme7f5qtebetmV5kGTFsGRe1R57OZn+EKXdoAsz8oEDVKzIm
ubKTnsOe/yYEIx05d1busrXo26/cIAFdPV3Yn8EaeCCTFRCZWxLoPmzsqpQw5frH6FB2Lizd2atK
q2TbY3SU7ON2ytEvu6fMySfsTZFmjMhKKguyBnh08FHv5f8hnE32AZJWEl8YUd6w6jT587W/7WX9
+Ap96yjvVYSNCkccB4lqtJOj0zz5/kk7hV63lPvgV1uVq0KAb+OqDk7fgbEHCuGabuEcqsWL2uto
YFj0IFsNuU37C/ycQF6u5W7FtLZi3jOfuZ44fF8jItowPMu736eWaZ9QwsmP7DXZDhytds5pK/Lm
qXehw03uRbK7vFZlkqBffAGXhGk7d9eu4N6ojpw9R84IzUUfkzxCWh8hsVTZyRcRq0F5i7lF8KmE
ED0sePeqq1dPjhT13DvvaGYL9qMXNKBdVXRcL0t/r8iXkdwOwra9AIxOQ0NdO2POWYUBb/tluIgF
a+lmjftAoqw8NHCzQStDljcj3NhjKA9DdPSfbaTxsmzHU1wA0Hfrm0Chv3AUEqgawb4tP+vjaO+0
ghtZDZZA6Rj1TjI9O8Dk/8bDwJWflhcIcDAN40rg/wPf+c7B9CH7tfEiSTYw4nKbgAJqjsodRgfa
1Yl75IxC/X4XXL3YwC+GythhhMQ/u9Igr68HznbyG4xFxRBDpKKWDY5migtBPlIbiCWiCUiLCZH5
xMlNQWSz+6fovXxiGfAlGIeS88Zz9ZONsX+DzgJBeUOf9ZddCkRu04qwL4C4vVLtfAFB/vrCWC0G
kSCFgpzDnrcmIz09maNwSeSzAeqrZ0TqK08/7Ri6qN2y99ipdH9O+TkPARiWv1Fl3iA4c1EJQHU8
X3IA2skZQWUWN7LAaolbD7vjW4LGhrB7A2+jTVlD4hgWVK9Um+YxHTMixxRRDPqtW0lejGOcWkvP
VFlexS6E0Ylr8yFCYZhUYPK/68LTEO3j8W5xiIouImswksDasfus1QW668XJq/c6P9hVkMQJebTQ
WAgIStwWl6P1B6ru6ajaspRftaFo3sOApOtSv5m0OEMSiw8LKgO83V7Wnf+sJ0TK/ZzERxvFVCYQ
0kyOvQruDkbCInTfr/Fq0nJDXFBZXTdtL4bwDt31S1W1fSx6Io8hsngbkLU2tHb744Kd5Zb2fwbg
OjywkECYzdUAZVPRUJf4FTwsukSHAooJvQQyWcqYdj9ZSf1+sCQTg6fzcdbyMMcRbF2bjZJ1xesO
0HMbtNj3Llo4N30FxpJtz5qZ/5VqZEuy4hzkcDb1Wtor+l08VRXYf3OKUfChjgkLnEm3Dm9DgMFA
rpkkVfWCm/rADeykiRfWrx1rLNJXVamvYgzQ4lT/rvNVOBRKQThUBuKZ7F7MUy0R7rXDX1Xxvs8H
xjq3J+7k3z3eQ6Z330xtoHDXm618jTHmZ5AJa3tGbUFbe4shehGJShFOLZf/e1qIIPqY0WPxXesa
mSmgZ5EwOBmOEIS+uQ1Q6n3tvBhlh9WxctkVBGJEhGhdbKWknD5XKGvFcllChREI/W2Scwn4fQQ5
1rVeHYKUbeEUAuynT6/eB3Y0QTjWs8cWbWbKI43/WlM51FghT67hgr9fb1tE+2tn0dgBOhDNH3NU
1e7V8fHNxISqj+Ujs4o8jhtmp8DKzrXlRKgGIpWoSK7Do9aqV1TukZCy7ug8OZFa6DLSC+vD7Ug3
rXfS+LYgQh0EOlmo7HPYdF+nchDQsE55QO2dpiv0dF4v3xx6kq+k0Q81fXaTMfO1RZ8O+lJixP4o
+faD/tq1SLCnFVrQN8YizANtNYTQbBZm/AW1PdKZuBqYwtU5E/KhIQy7hU1wwEQq4cws3g1lKfFp
us1Dhe+S2orUmW/KjzAHragJjDgxGmTcWRQVAr7EYvAFoEDbwzMFvqsVyF78c0F0t+4GjaiDCvrp
byoLWGMiah6/zouEubbo4JdGgF4jIUsI6xhAzXvBdmATIe9W4UQ1dUH8WoM2unwjLsX0XR3lfplU
vflbuf9l+rJ8B/E4fU5FrieiLeXgh9+e9ldeffIaIO5pt3kzk1Z4m18EzKXuo/TFe5Auk5yCXs0e
u1A/5bMa7ie8Obp5vR5sQ7NdDZMMA2GKxBwnU7KeOYM6A3mL/NbFKVZrB1gvP9PXosofdg6Tnl6w
66p0PIqKBZnvNgtWTAyuTqEyePwSVywCXSEgfJJacZIN76PswYho37XkyvmLk1P5hoefMlsGiqaD
vce1I2yLBb+Y+/+vHFotuceW1jeo5TzQ0QK6sEcwnUzplbjChd4o582gB4GdDmdHEFlAf0h3Gam8
xyavKTqtJUe4rphFXTxr12clxdZbf1gzYx/JxlxyZyhfhtB8rWxLKI7JqdIX4/rS4xCLxPIdBO8E
iC21EYbkWaFZYZg0mF5bVEF5BgUWgafg8ILL2JaRdS/hwfMIrLkvUAQ6Ry1yY9XlVc6c1JdkaaVr
ccNNCfCUfVEvKp8txhjsG75XPrmkjgzAm2/m94rw9ayMyH8GyZX/4mME9s82XHmMx/oArssxxQYa
NsOAA34A+kkKl/7bHil/u/mO6rZ/HhD/C7nX0LyLxtJpdvHw03hTdN7W0v0Xc0leND9zZzZvVkTe
4grx4r7Eunz3k3/MXjkKAG5967F+WXuLyXmp4aS7rjMvMsoGTjZklJmSOJVp6+ue0UviYljidpVW
WvXwEJbfFi20g9THMeRetVnvHmq8eEu7kJ2Whtt45hceZvG0GzO2EH1MjpeEqcJok75mr91JtT18
Q66h2Ox4WlkdCZ1eE8M+2dY4dh9Qd0CcNrrpo+kkejfrKoupqFnIX+YPNjYffmDKMspKskXjBTk6
/f5PmR3X9y7Y2JpwllDpZuFwOez1njr3nKyRlKl2GQ+i2UQLfxOKpr2424kzf3q1/PJSOCB31Sco
rasd9JprY1srxCSuP1210mUFPRt6AAdTB82gh8VLS0twCfnB9NblJXNnlxsNAhyNzi5SSLgOK+GA
J1QD71myBOR6cGU7v8X1SzU5zG0Ko19ztaag1eeJ4agoC+N6etedglDuD9r8AoB4A3NvKrA7RWH0
zHso6lcv7D8SpUAV9hvjJUGri1gP3jjbbmSpV8xVMPAwlVpXgUyOo7k3kQ+QCK1QAkaCvSAP+C/Y
NpXrJQQWvrIxRk4pzAnJ3/OfyHBceXfNIDbjeIoaz6iSjpKWiOvAQ3JG9Tf1StPniwldmlsfmPvl
umXEY9DpzJzwTrOew+yAwZ8LPGg9w2kw4ywLdu/W4W6ry/RHrN3PQckWQEx6qbX2kfjiSeXNeQ1m
bND3E7zonz4+NeccfzU1heR/P0h4JhEQ68SHlYtVt3UdX10/JWakbnbJAtkldPxqokywi2zci8Ix
uew9Svov/9S30wSZQg0wp9Zaam0RxIkyRc9EtGiCJXXEE6+j7ck4GMwLzUIa1raauswqNw/W3K3E
i4nkIJBXp+3C1JnNAwPjOgPo0vLbOKt6fHlQvlkmWC06TUjqBiRRsslm8uu7s3aoup0ZgwprLbqY
bI4WHPjZIYylvSzrS5K8t++tgm1vNw2WfcZDrvFQuaL7HPmz9Bk4MF/UiqGm3DTDPuzc+F9JeWoU
oWPdu402T2O4TbN3rxf4jSDCQK36+H8zKKoS8dr8lfLb1cs6y4OgO2IxFeBWhKFq4tu5Xf8DDDJx
r7fpvpqslTMfUM2S5D4lG+GeBkXLSCP1ZsolJT6xOZOa03GJLbhQGCdlLEJ+RqjD+SX9I1JWUMFM
Y3CN0STNNTW9S0xfur6dwA2rv2dzY1941dyspAFwKSygYYAE+zcBE+4DJpCff7i1IuXs/+gNnNEc
vZF+lU2NlclGfM5Pxe2zvhor9EYloHo/JCu/Jz2aBHaQmXRN1MIsXw2e4NOALS+0TYTiH9DDP9dt
PjCP+W8gOD6xAAodHMcKhN69QFnOP42ty1PF5VHLJQP/HR12NoYVe+WJexy2rnldwkjLyLJ1QAaq
G66TmzrrwdFJ9ExIf/fWpJGKKfKnGJbLF/veNzR+VU6O9cMQFTXsQeG8Sf4mcFcx9e6iXD/Y4saS
MeNVgPLCVd7lU4x5H9j2NNER7iMAvw8ID6yv8Qv1CtwL0U0NDgS4AL+jQe3E1LM+BWX3I6F4TsnQ
Uj3VmBfPEbmwNYbFx3X06TkMepC7LnqK5HceRl6IXN8TQ5MSE7Jbze5lJwuSel+PYkGXpqsHdtgH
Inm0/fzZWxR+074UMPRoxoXUS7nDatdCVshBxekbo9Uq4FiGfvOxcKBcpXFBtuhouaHFo93ic0hd
TPE0OsBhtInoPmn8PSAG8HYjFHIcrZVhoFrqrE3AEj3hV8ZZdi85hOeYRLNlpB9h9JtXzeAXgFJW
Y2KE4neGVql121KK0svJLC8JTJhnuK2yZlDYbons92XGVq5MKTPftxMKNSjRwMWXBPq0REjZofpN
uZchAfv4KwBLjCwTTFWWjB3yJ4ykW3OFXLVSEL6jT4QBQdT1/qFFDCgX6wa8WM24SwKY09Zi61yO
de/wAep8+wzvX78iKd8axgLcYmZOkw1cvXVarabGMnblSas8hZMKGVMNuIVYwdQm6W+rfVOOqJne
KlpHFyfWgp6Vu/sEzBi7p3Uz7C58C/LAUKV0YuVt/PLwmTChIZIxYGvVCb6/AsfU5Imo74AMDHM6
ztQuTdlHQrp0cUOIbZuOcHHSdUJwg569bqith4oWYPA8pq4lSiE1AkXhs94HhnKZDkwHSzhKEqRo
ibB+25rswfbYN3Ao23KDnaPINQMYzhYo04bpIfy5655mdtjQu68lrFm4cXBBx5FQgZvkW8KuegMI
UoSWKkvXuTIKZNlEJxVLEhFMW8Ib3CJIoFjqFKF6yFaRgZdSSP1rLpLPrtoEZwmaIH1aw2RD9vBW
lwCYkjwgeuk0Fpxitv7jlix4dJAW2NqDohtr7eXEVF8il/fuh89OJ+Wgzw4vK4NW7/s3lTv3jytH
Gfhxc/fHmSzu6yWbvkTJHJYsDDANZjNY2K0hcCnVyOVJ4h2NUnQ5eZ274Rd9XX7YGQ4uPcZYI/4X
eRiZwqhz/asc/F61qEhYuxnk3TXJGk3hX4lbINjgqCrf0J4gVMInwzNElHhWhzHK0yO63Ld8HH6P
Nt77QSNP0nNQTIYhigLtPnYDUk4S2KrRUk6BqnLUrpKUkbTm7a9OxX8E6aaiquYiMW7uK7a0sqSG
f+tRmL2I0WXY2wh9zbiUdhUwSqfm1bDUHygKEu2p2d6NNECtXwr1ecdRh6iKvG67KWJ02EDkLJ69
bnDUG657BlEGjK7rrCLNAkj+uazn3zAB3nQwxGk1pv9nUL7jIQzlluo7UMFhuZJzqr7enhO5GMgB
u1RQP+3QlLkD7Faddxkat6Ot5M2D/vH7KiwWMT7c/fdPALhOTy0em6eY7SyOxAAvQtI4s8cbf1CS
Ly1QH8Z7IACFliRyPhUunBDDI0Ti1Y+Ol8WoURIZF4rMFrXnD6eDCSB0JW09MGxMd3Fgy9uP2Zcy
xK0+YBkr4TkJC2Fghj1x7iUqJEB4e5QSbEPA6k7Dp++VX/LuI3SHn4AomEbv/joLt9Cw254Te/X+
C20/ah0/qATQxDQJxyN0HoLQicAnuommo0+fjDhtDpmAnYCs0fRz67Ro4Xa29sjKMGKO2oKu7y5O
j7bGcIX33QklCAYJcbnWh6FfyuOp+mv33nxmmVtSnx4+/736QUdmluOVnU8sS0BBe0hedW0GxFEl
ectmIxkQAXd6aPTnhynpwOP/7z84e20bRHc68HTlxiHBLF1NMDnQZTK+K+txI6knv7Z8FpiaGIac
J9ZISc1pqG+As0AuPluZNBZOpMoDGJCdURIiTGM4TV5s0VfdIkxrSywZC6Us6me11g5VjpRRCfiv
SGHzbolEsMlSStJnsg5B52LKZTcrp6Y01bKOIgjhW7Iz+oZSBMUNGmztJdhubYAOjZ6ZHVckhK82
DEDVJvkeKJwTkmtUbfyesd8zCPR4dmujtFled5Yc1I9c9J2itzpeNrS68Zw9QdBgNziGCDE1zOdC
8dZlIP+46WOSwWC/IgW11N5jDG2A2xz3kkSBQkzGB7RyGkGVdxYrXrW7qf1xCToPlH+wv7BARCv/
T9LFroZHR64PryBJYJcde69V927mHCl0yu1vxzc28Y9UjumsmqJNnmo5llhYNWpwYJrDZp2/YRh+
fwKFOH8J8OqE5NNubiDIgpzgsMFoRztZ6NRpSWWreQaBRp+Out88OpHq+hYCRsDNG7n14KBb80w/
VaB+yb2aauLlRwKli6UBn+cQwrT0hx/Ls+pEBL+X8MhtR86HTWcWfCiTnLXHrVav07HdLM7Y2Lv/
N4G2RiEWKJnCb+yewDY6Dwp8UF74KoNGeVSfoapH5WnS7zGsG4mVbdqiTL6pu6CtTd4UINYA639u
ckOuonXMbTY4SIO6vpD4Ce+NfpGTWPqKuZU10Un+PHObpaUONLPEa3iyLD3FXCp/ejRVZfGEXcq1
Z7FCakX8U9IWna8utegT4y85AsUHvblzaywunxNnU3d66Wa6yUa4TjA7VQ2AO7QAXQcBGXZoDuA5
WdnlTr1i5MRJQO3XyPLbhMjFCELrJ4pGd50hZlUt6rnhKApOsLTE0FHavC9yL6YPUME1GonGsLyH
5e7q39V65FWeFapdWkupf5cl/XEffJWCaXiDp3MczBLrKEZ7PwSw1tA3t+BsoXfDFibW3u/ghvyb
qIx/mEaI7F7hs46KmPIlIqgfE+9Y9tqC/Vfga8SHpSB6/QqlFCRHIr/2Hfu8iEeP+3q5rKhSEIYT
kIG2p4wWSoOV09tMLCO1WGJ30TA36jSr6FiH4CQ4ndwTfRv/ITAJ1TlZA1Wa5nkeWONMegqpDrPG
tgFLxJh4pomMDNU2yPJsgzSfc0mgRCsDYrnCHgXtoeImt2K1Q2onm/SaeL9JehH52FtlcnYVJL1A
wnSbNObM9qJko2tuUIlAKTickXSFoyK+zF4mwJEgI7zWfCi/MA6ut4uDEuYaSl8yjlVSF2fMatTk
gm0s2tdAs1ytXSy7KJuCyB1jh4hZyVAw5DH1yxHQ6yUW98gK7S7c82Y4Nu6cIJRjc2wjFLUkfGKu
OgZdG4lIXy4rBx4qbx/qQ2exUc28Dofxlucz0vVV+SmjLr3e0zWbgSCi1kAJ0DPNVGyRJYOrMQ6w
+6JTts+hSZPsr65BumczCTQXBTePHbtbcYw0CGmf9cniO45t05A4jNmYs5VAZYzLMvcsVJywwguw
V07yfaM9vjI8stWIqYPcQmJUWdaKJP58uY2eI/luMkN/O/FNAUw5afjjHXuhbuwQR4Ab9l1jXaeX
dtgguUOXoMbyDRRCYPEEvxnTWLw6fkkqc5E38mbpnC4XODCwVqMkQBBbDXB7XJJJ0ih4fBfg0Vqt
KI4CLd8FnPu/aeR0ypwQ9pyZ7ftUKBmLPLG3aH56Cj9BhxY6kdFgDK1czxzXZOImJlCYTNgRL92j
dI0+w8E28OLRA8SJEIofYBvcXNBgG7BwtUHDnRioMhwcwi2/NHn1dr+d9kuGtX8jlv9fpHZ66Std
JBjpVEOzA5BZGEe1YzbyW2Go/XsHSJezZzqZZOg2NRmz/MwayiIfq9Z8k0Ix5bPaj2xItwmgvyS6
leDCmMyBQEKjd+YDDWISCIOQEVmaWf/VV5R/k3k/MPCpV+qmZ+InsbJYC+Zh1bfMA6WREHlw/yps
lWbmfV2DxELfqcszoeX+L5UzplzyxyQyoWZXRnXlQBFl22UfFu+yXzqqCwRTyqwo8UssMgq4+jCG
50mEdp2AE34+X0V+Yh9JoT5g3+k3Dta3PbFDqZ3D4mwi/qmmJ8xWjYIsVwKvxUheko65DtAJiAl2
yfD9xyVdFEe80aB61u9lZz4A2SXXfYWq/6G+v4459jxfQWv/DikzpLvJhfBNrKCu4is4MMLp63ip
6IzEakn0pQ9PmMYHI8pgSp6Jc8fHUrU+frRMV2wt2hE7+yW3zZQP6WIL6vZEF65TLNUfAeiqGOXv
7dBMoRJqEXll79V/UvfxOGvr8JVkzV9O5iwx5dYNGWlS6QlcdVC5P5fMvWi5YF9IoAQoY3RObOv5
Rtuf2xdxQSArVndH6BSBYXrcm4pC+Ija2NWKKr1FWTOEVqPSB3kswNsYrb6vP/R8g6oGJPYMPyO0
UEucCEZE0cBsDJrN5LlpKLXH6MRoYnL/uVelGIoCUq/j/SAhLjAwIKQz54grtzhsRc7JNdMyEf/l
CkHBY+ry5t7S4+mCCQAeF7DiUnDuG3U4t7tsw5/rYLuj2Dr/jaVbi5l/Q1o+fdJXQHd+M1GZT/0N
+qIR+D6yKE0Uq1fP2f0WSzHYF9FvzorLfxb+7Qe7dVjnLO7KP7GlxeIsakzKFin3y8gTpCYH0PXK
npaALBz3Zt8V5BoMSS3RNQ8g9WEpm+ua5T52HLIk/vzO8MwBLRjJAVHJnDXx0iWSFoB2qmXuCAZ2
joObfeeh49PAbXNll5N5hbhRWxAF78gTKgWBMyjmCz2RNbAcNtPoO04sv8wOPElNOklhNMP5SIhE
ZnwtMFlvtbFyGRwCeupWpE3spHto0veuDxVMPYAzKr4mdpUmXDO6Ugxrk3s2ldrzfWZ1rf9BhkRp
sk0hXTjJHA/0DBgoF4l4vtsdUXYCROc7tdiLpb/537Pghzvz+rwPXHy3Sdhc7//rm7Xv4Qz2kRaG
vEF981t25LV6/FF1/nkewu5OoL8PwBzF5klnOxTStYOTckIXUM90lyN1uJX8xLBRuoBfw6hYw3ZW
SiEC+LOBMi1DUZQe4dCyewp1ZZw3QPu/+AR4+ttAsH/Lblm+3TU/1HQ1O9negnRW/GafuvwQ/+dq
sQJ7yYmPq1B8XVddwxqfO+1R06onQo5LHrEPCAvZ89yceSzJr9CGuYEb7GM4zkxJB81mPbms7RuV
9oxw6PpmIlNKTBzdceAMRJTHYmBjDex9ungnylmAhzV4EWBNhqzww3Mx6g4Hja/B03rc1lRmWm7O
UL67Q8SKIfjxigdbHACfIV3fHlvoTtSROP9n2jmI6ZU+TZ+MEfPRS3onblVtIgoKH6ACCROZwWhW
Ypp/HGjK5n7tYktLmzUJ8SSZm5cTRrZoGTYkGSvxtBPran6i73bUbzOoTbdIfbNCunwBOk6gDjAq
Q9o06hIJcBV3dKYEsEoDFeQu0Nha3cnXZGZbNeo3QMEL6VVhmSFZhL7UlbBcOhCZ/DMajFc4xKQa
tXOYzlLYSRkUX5pmHIF7a+dV6Cpzy6g0ZvPHIYQU1aY2aPG2G4nTQ5YLrrCX7jT8LPT7jeE0rYny
XYa6P7dbQ1Go/u4d5s1sOD7LE02V8tg8XGEI8qQPsOCk8VK30co+snlB4nsG74ZBbR2uuDKvT12V
/u4ahhtdlPI2zN2bHILn/VgC2oloUrbIAllEap/HEQg4G516N5t/K3ipKzoH1KdMTr8LJbyQRAQX
OoFB19MZGmZVPUw5+wGzzcUt1mHiEZi727ToMf37B/triweKfxUoFv1H9YF6WGgRtEG5ZEecCpR4
+wTDiEvsw4F6UxTYTEXydUNkUc+6XshcBzVA3qKxWQNPiBEV0YXXYXikRpuv8ZAWr8mSvm9Kabd8
AE6tMDhGxb4UDxdXtVUdSC3aSUktDgW+m0KYqZy/a8p6zTs1cwXPV6x0ucajMfLA2OprOYAnxgu7
2ofnZu3hwpDiwAzR+mtfUxoZoY4h9NVlUN8sOS9g+raWFpPptLgVa7b22WtHrVkAqHpqdtCNK7RP
s1ACz477nMrtMSXPmYT1SEQ6JFGigskvBvJ++ri/bJHGkV6SQ5vwxOHwjsslwlS4wDnh0j9leIj6
Y+vr1hPtvDvDoAPkLIfbr9Lb5lERFJPgEKsl/XqPh16qo7Mv3n9rZUuF/c+XVy2plPU0dp8xXSsI
InzzCKUknHs32V5r2E3gzb5WuiHYwS0FK2eA8Zq/61rbPDnxmbI93Xnu+oWbJf65RhG+E6hq/vE0
SLhjABfuzwHGslH4BO+UhPXDYozX0Grs3UfT/WMW7sBm3bwxBJjrTP1RK0tUwnZg8wEe46hfF9cT
slSmr3EXuMDzP77hKjusgziz7jwVmHaZxGwbzyb/plEqFcXW/8yi9ibeuknIBNd78HWeZ/akQ9Iu
v2ebDEOlPe9PXvbMc9t5/hTQoNyvUovkD0KoxKaRsISaPt1gWZxaUTtxiY3Yo6WPTIlHF3kKk6OZ
oPs0f3Otvv3t++DQj6jt3cPL1760G9GmPhpa26lGyMAJL1hXKE40SdgXZCzOiw5D93BTftnD7WkU
0TkmKAAJs6rc8fegSgnXla8yhO6PhEVHC7yuM4mnCQA97t2H6s7F0ecvLE+hPmF6W+YkAxdRddNO
L2Iknuzq1UyRmoEGpWriy2pvyKQ4KjzMohgdsh5lMJFFtF0Lex/RTo/gh7OhEMqcDT0ZyZL0xhvf
4rN5ZGT+POe1pDy4zVhI+Nh2vJsNzyk9cBrjqga/9wXomfrl4ILGd5yUaN3oyDEfFrQk1SirO6dv
/p7ybVIt6NSA9n4bnnPK+U7jZhsvBBekmjuM+V35miei633nvhm90CmQ75XS8+seX+G+1oXeANN0
cWp9053mSDo5n+pNM9pLRW/nPunOzYWyVbVbSjhoYMDPpEQmpyJW1beFw3vDxj/8rKy40wViCt8U
U5xuHJnj4mt++bCJxHdc8zSS0haV2VIoIqyKuSqs6kIo/rGDMPBe43Vf3ch/BNLJOx9eg+hnsczY
prB5oatZsqcNrCccMH1ympD704whtSZlDtLkTOPt+P6NtSeSmDCcTGRVGSgYEc/AvRjziAkMI1ZL
/DJGm0fxbp5j9S63m+wV5nUbqXGBjTZ5T19fiE3cVNmUEZEIM17Nk77Rins9J/UNxUnUF1rnO7Vv
XNcnmiQPn7lMK3/PBXGEX9GZncdFWWBcbYdPgiArWTCefV+OliAl/NCp6ulPql+sOZFL03JFFjeY
f4+zkzn+QYwO/uIpc7TLbAIngnpUQwRKr9MXexleBOi3Fcopd502ThtnpW7IaRXrNfD+sjVOIE4M
u+m1IBE8nY6qG2pU+VGAxcP0DwMPdoTqWPLDsxP5OGIhq22RYpb5McWcTIIB6BUMZh6pTLpiPIf9
kjFqXguwuhSt2ZWZxHpjpKeO7EQqkG8Di4WPBxm4KDgh7vZYnFseMf/5bgKy9EEir21SR8/71rTL
X7xKaSHuRiwlIg/BJ5mYNEeOy6VDEnTwy7GOMLtVERvc20Milhe0QGAxtLULhGlc395bTy7X/yIf
nmwbzZIOUf8URANicJ+5h7auzCrXrEnIb3i1L46+x/RwO0EApiCOqwfBU0GZItauh/zSM/E7HtRf
Fw7fgJrkFEERQJuBocwzTurBS9m+R6KPqpfNLPIiPJI/8O76PWZ2OG6ITPCU+eGqWpuTKDDshk8q
uoaD4V8hhcQZ+E9lPcegNQ/VawhUkBl4TK34LuhI8H7dX9wGMSMEmeiZWaJx6BrtaMfRfK3TlAHq
rNPKZ6fKTV8vIDGleYyTQGp1x7XG2dkgvevP1RR7v3q1FDFBN7VzzXhe8nLcCfg5cnVvN58tdYnj
s+lnuqwUM/RaoS2SUm5Ypz1XGkB0J+h7Vy4rbaD71FamksH+UKFflxbvQc4tmblVCr9Gfyyx7Dbm
bG/bROlK26wBvpXg6j2uyMIStTTeKe4uINVw5wJUwCpzpzMfpINTgXuZ7Wb+INTZnMgl7w25rOQR
Zpfqw9uhstb01mgifJsFhboY/xA2NhFk+2gULH9bgfdhyUv4IpAV0mmPOTiz5E6U9zYZw6D0RCMv
qgtxdk+AyF3wurE2A0Sy93wpz/ncBI6P/2HldOknT4Jt1kMHqL8Jk/UYabz1sTph9ksC6lVlemYA
kgjQ9n5Vqn85/FPbC3QQaVu56XpOf7Y41w3BgC4tAr8t74B/PBdQF+wnFHTREIzDidV2xOm4yoP+
PkFNzBXH9ePMdskdv+qxeQdDEoVdXCSszrK7e0c4Lj+7rUH2cx01tvjG+nTQDKMRjd3W399vhDNu
ntUU+lHVUjZuNjMP3mLgpszwKtSiX6gnsJDulQ/zozQyf2gtIswqxM8dv2Yda1l6WQ0/kWUHcQQz
vtjDB6NQorHSZ1CpqfzwG5k18s2l7J7iKeB0al+YojiUR+CUcuauhd29kWDXFsKL7IR94pBOfQnF
hv6v0gsCEtOuJOZoIwa0LwUShk5IixoMwREX4uZa9JlzmcvVsnoam1+f0LiV/kOJtDgkJAT9Y/fX
+m599QE2nyajWAKoC5NJBue4oIjSPXbfVsY9RmLTJsEERbMQGMZQsphnrsxahp0dp/3iXsxzuO8M
ajUa+JF/M41KF0zCGRQWZ/lSMVDoAa7lPp8cIzTKhiyUVbPvjLfncQxvKJNdIdiFQrICvXzOyw5K
ikT2vdBYvyrVwmliK2nVRVdnI/Ub4sbAs0dLzHlIzJBtnftLwii7OXwJrwDG4kJDJJ3Uiab+nzci
Ft6geEHPOcCx7bsTFEzvYDhUt/1BYgPcSEQv2iGrQEJw8WsKq4v8Ie0infi61dt5lgni9u/wopA2
5f/VFPBg03ez+OT7G2ZjbYXljwASiy29Nb9FbZOXGaH4/leay8k/n/TwnMB7OvQnT9iYps/nryeB
uKrTLq9CpFjIm0Zr6TqQ/0Uom2cYCksJIhiiAYxwYSIesmycQarT5lDTh6Jd5daHXKl+oJ0eBsPR
vQIQq4DNH+10y2+O551H3ayF4sLOFE1IARpI7sXdeUU/JJjKWh2ucWORAYlYMq4TwQGDK9XeSBsd
aJkwZ4J2+WkQk4CQKO4rcvd+nC0rV0Jw6215CAcCj2TZ1oCiBZv1pqmVwLdBPCDpBXTMF/b3UjrE
zBcrX6QJjnNay9bdZ3a+nJV2WKnh8Qay2WNqqDMf3ztmlNCdpRsWUXQ5lNH3o0ADTc+bv2MStF8l
GLJFCS46kfjUamIojDYYBe5Jkck3d2l89gNE6PkITwIGVJiVedFzwMCE20iXAHAMCKfmT1o1DDgS
1r/GdNy+SHYiibJClaP9UqOBsbp0rqAVhr9ywCLY4VMm3hq3uGdg7nWwpLkv5/VPobglkN1RaU1k
eidEcvBUTQfzgcaLIJ+e6Jg9wtpVHnX97bX4H1up6zKV90w6y66b0Hq2lbAvSqF5vUlo+DfEU3NX
RDSxoG+IB+uW/pnqHuP2DemxDqMpBCluoexSQO6B3HhIofocSdI7QJjFk48B3oWoHHmrweBvaPm/
guSDHDx6/KgMS4nTtzSnw4Vtry16gGGYIbSlpJVC/JG2XLV0aKHni9Szu275hJiLR9LEbDrITYbp
5aa30kboPS67hi6OQNx+I8I4WGitz067igLAVSQoJcA5eRO4PizQowUzqivavH6vJmoSXMyZ/IHa
Frb/koLIqjPFHyMB/JLE1IqdbIOAsOIWARZJo+8lsR/ZUKdLyWENAVnwMbfyMDeZwDAWH/2PMIPq
nrZjKYEHhUBiDwqz45iajF5KzfQtL5jWhRMEYECsC3cErYyNFbpceOhX7d5CPUKJ7ytS+ohNVtUu
RjBbpWPJMPPAlIdwqy5KixWjyPThpKKKa5Fc3DgLm99gLvOnqUtXsdg36JxOL5ZK6qkix6RC221j
wxmGDrnuOcDm4VuuDXrgH8IKZZ0AOQndwgm9uayC88jZQYoTA5Rk8/vDhdovf8Oam5KJHycCE3Dp
eFgcriNA58fsecK2+tuxwW0yqXPr/DO2FRlriZEq7xZxkIoQgBYIKhE98umlN9ylCmpOrx+ZBnZU
AGl8+4G/ZLHaE7YgbX/M9Z/w7lqUgs0pWKgyegDC/4PS63CknBTWRPcjVjhjvyAEKIdhMK6WEs18
LsuZpinGZ9DgAnK/Sy/d4kEfFDhHcvrMlgSUKRBS7Nk9W6Mki2e6CnBLgLpI+nsvbdDBDTYyPYoT
QJV/XxVPv1/OYw/DMLvvznWK+2WCnAhoHqOpv6Mq6ZUwV9xXKD9nXjAOthwZFFMDzPaokKhyRP6l
K0Qj0VNSAVn56ouwufQiODxJhW4qJU6mYpBaGJGJfgdb+JLDQ5Gb8WkmiXOoTDT4HrHpqmLGfYy0
nLbwNArKjI3JW7iX55QRfz3WtfOl9YFtwJhUqS3+QbnooIsWrHzs94KdzamPoyr0DJuHjUhvkEvO
bDzpa+T12gUpTWSRhsXUgoG/inYVMEXRuE4oX/O3VsJzmWYAi0xkAyOY3FG0BCS1wO5FoF4OO7ev
Kmz4A020zJKOy8Mvpl7530eJ5rVHU/8m66mV/Wn5arlgfPeFlHNOE+xsAzsg0KFQw+7BBMROvo+3
W4J/CqhtQt1Er6iyqZlxTxY8cajdHKp20/DUom/uo0T7EIPEFiA22Mu9bRnbcY6rPkESY+ifYDRi
ffwdso5pNsoPNBaYxMA8kMHXnkCmplmQLLYkY5een6tx3bud87BgSMUgsYvAB8j4q9vgDdVXbJ76
YejeFxuZT4mPloF35EyUg9o0j8uVqla+heyEHopCOOhUDwWf6AxHtWcghcTDZOk6MvLFmpscJHTL
Dkmr9p8U/yWfqWgq/yO15zca1vc3+Z0UbU5AFcW4bi/GSJrWgECBfC+w2tVJMXwSE9zIRvVisS2m
JGo+A2+DQ3eg8c/DvHN02RFK2hccLzpXi8z8t/5XNbVkQTi338Bxxx9sUU3/YYZR5MKRczQVpf1P
M36oHEs775peqQ4hkatPpDgLR3zIhxI46dodmSfrNuWX5vE7J7NFRMwBFxXrpBX5iwQXhLxDpVhD
jAuytqCkjrfYZDuHBQpPTOOL9sumuSQfkhPewev8vCWjDTC4bTGs7xYNkKn+z+MuvcPJfo7lFWNc
zguz5XrRyEoWEiv1OLNH0eKis345DQYQEvhhRNrtz5P9UJBnXtlR08/0X8Y5FzLjr2uIpUIvUXUB
C7V49z2geRdRc9C/gos1pmZYfMTt8vIlA+OQN235C/sUbROOjO5ZNg5f+pJe7h0bykNwt4uJcOBt
RW6QYsY9MUMwc10Gij7O71EPMM78wgreB/xqGMEI/oD5+dI2bjUlKdGG6I8AO+i2dvR1x45PTCgx
O2cnhdiWfOZT9UWbiP2yRTpUi/I2dcIUeZMhw/FK08A0gJqhQ04IoPywabc4uY44kZj8xHWPNlie
l5/Y8+to8yJN892+hMzvgxuWnysUotGqZ7Ak0Cu+CxKpir6vqteoTMB/0zdcr9ZrdH3U9hNWuLPQ
nrI1RH9x3Sd/ts6/xy2OWgqkZZ8MSYzcqhvksD/vM6ZNJypCLuZmP0cH1dDx8uqE0vALF2ylkaKp
cjuCHbNaPnEziXhisccB7DbyqkQm+qbOw7aTaTDD4rGA2olcyk3X5b1YjBGWgvBiUCHTLmKedLNW
1+NNgkUaxKOwMIgPtnijm6olBe+e6W7yIZNmM2ik+IpUVmXcoNpj8xIoCe0n7U8Bf7WC5S5G6KyU
qvrcQY7fPbH3FKn/zRB7WbiBfWZPgmGt862uv8+P6Dp2r4wGJRSuqbQDWSE2PyCy+/JI22bqLqAv
s4h6+BDUyK87b90ec8pHE95GgS52IuNTVqTDrePjb2D/HgKpZsum+HOwfLok2u5WA1oc+WJmt30o
rIEpTq8yrTVKAmtS4DsKsNt8m+fAW1FEeECOGq5CoTGmpLUHVw5TQe3jaGsUidukPJo2XkakjR0g
cYUJwKrNrMWW7HyepQg6vVdHaMhALszkLoLFfQ2PFLn5BgG1BT+6kcTKTj01HKOQOKQdvcP7tmou
OG0JUDN0NHMB/LXd4mFvMMjUHtBrKkLqQnTx+RhJnDuCtL0p3CVrkxbadrEBO+rpTjnIdn9wjOLO
2Ywpt+LwtZJxAqWcQRkE2Z8B5qaGSZc85yQl/kfRXIiCmqRchBxb5J8xDnXhpTgRvpbW4TdJObgP
O8tg8XuCSorw/FbD+mMxEqossINKo45SYzL98ZtvtTMtxqegVIZD4CAZsF3I07E6tcBtruLFGmU9
zpOy2xFzMebqCNxft2EO3thf/dRyKCmvCxjVJONBiVRrxouvXRU5CoYhJWweXexUGeVp8M9L0Oh7
fhr+D2nd2cHT8NSjgnvnADd4XpurxVQmGaSe+XZiW38L80+DHrAmgVLq7z601wo8Ew20qOanNLSi
Yd/9obgN4U22SxnI4fp9yEgUBnwBFzcjbpqBgudvdLfxIXF3xIdV2RRnEVlRD81uIS+FfO8ASaln
a8cuiDAZoT6VyD3FRIZglxZrG7otebGkh1O5KO1TOj9PVLoep00D59sGmksHvCO7RykvBU7xUxm3
hEM2U57wlACfT1Bxhw+w4f9VOrq1XNIy5cpb50jUEJ9mGkdn+cGjlNS8MpddOKje/lIR28HGSMxz
sMN5sTAIawstPxhyPL+jbrRTIYNWxWx29g99r4NNIL4cBXKPynaBAXCT6tUd/HE/nWwgk3+jWxmt
mlo1JOptYUCFhdd+i+BOI6qW87n/lfnAks98u1VqosjOvFOmeAH8cvzLaAL6r48ljKHd+FQTwcRz
CKsr+2RXMwv/B4BS3Er4+nOvRR3mFqd4wTuvoBDQqh2VxMQ9bHutXfyrZ350XeZQUE691mpmCJ/n
o1/WAtuc6wspdLheuPMJoa4Vm/jOsgL/qj1v8SBEFDOpaZlu3uly6vo7PcYmNB4XJbIx9Isc6Bpg
d5YplkPhaxUBFJn06cI2OuvIlNmXSwBGafrNLAnQ9fk5WNzOjt5voPBfgDStVBlXGZ0l15j6a6vc
ixxWXrvGcv4XkC8w/OygzWqXbvVX09SkUj//rb/uTknW0G9xGE22SX9dYkL3WBMhzs93g26OjmR2
H+tzUPNkuscbjS53IbMviQtKujLdeGUyVj0V92syz+8Cd0rjV2hRB6gfzAjeikJ4iSNvlygt2vYR
DKTPBqHe3eCDDS7oqOCz1BBeVlexkXzfvk3Nc3xtDmH8vdJrEKY/xZMAaf3QwcM823MmEhx2FOrj
zSuwKNc+dv3OfQgj7TOvtccHdxU7tjAnLeLLszLxp6EliT0ogbBAjUGL5LyJ4g73iRcY5+KPhxVf
PcTshQ4I7VDJckj/pPFIJxJ9jlfMS4LxsQLoyBnedwiMMTnO8Pr1r4JTxPFPB2SsP9PEpcdqmruC
V3xiCD23LZk2mi0cKeOHmbk/4KwpO4R4WylVAx03ssG02GWW3dWeJNKXvYABMjeeX3RptSnAV4kr
zf4VQSzKq140n/jQy+c9moENmJqqaJzo6I0luJdQ9pTIl1itQUMMl09uB3ufaXPd09DdIW6J4Rv1
ZiGFQ1RiVLH2Sj3ZV3U3x49GMhxU3CqvuRuX2Zs8U3f+VnJdzhci9im/kMhvPi3G24Ngp8Kt42Hj
Dt0YqsLHlw0iF6PmbUl4NMoKomcVQkf2z1LxC7buI2+pLkQ/NiJlZat5ju+KrtnI1ZgOICTX8Hc0
fa4fyFocWdt7wxB8/aS9j9xsS/Gvm9xA7yNsZl7+iGRR46d8JpGeoZnTEgat+qL2h6Ia+ho2nrQe
LvBZhaE2wqmcxY3QiSJ3qXOOz+eHNM7DolPRWCqWEZnHV+embK2MDXmPVP1SH9LBD1JE7F9kaBGL
MjEEa4Km5aoV0fAzmmZpDmgMm13QPu+hGVYJzTId+c2MGkd6vJORXS4Zp4GyKg4K2Q98xSjpC91c
y0QQjuQaHJT2hVZl9159d/74Ynppdv4cmDMdSplWZFK/6R/ChtZAnXVHb/pQOlBVqnBrOkiw4k5g
Ie1Ck39CdfITuSJBbUW4QthAnKUs4SuBqnGB6DwrO/jRJm/hSbwLMX9X5tQeMZ7XmMG/1ZWWvk/s
dnjBf5R6uUluWwIRcAkYvFLNhdt1QBieuDzqQHbiBd6YR+ZuHrIyrxAUMmN5PgHJ4kJ6wRGVk3Ln
PsDTwg/G4ULRsvQvXGEiS7IQxV73vLDrovUXs1oFl4v/5WNi7FB+JmmneYBuxC5/xSef0uKkQ46a
MFxJCn8E2gaM0Z2TxDL+bYklwvaLxP/xzlPXCnoJkObY7DGbC0ZbjBV63aMvoYhcZzRBviXJtzFX
T0qUDxxhI86IANgd67dGiquaBJiFvpjqJSPURqSbL+UJYc86yIyiJf7L7WghiixhDO8ge/0HN8t8
2kOk5M7/MDQFqjpMYTGxnlDab7bNeC9dyoDWmWNMptoEnJsfkIfFgsGcCe1cmEhNviSlfEPzONSm
fntWGCXjOmmPWG/iDaK3FpI95oWGvQrw0Ag5kpfARN22eVQIRgAvtHn4XFJn8Jqn1hoaESHq9Dnl
5DkoVheft4BBG6KSAjbvNnASMkLgGgmDKJQT8dZfuIGCvEbzS6vJjf7pKsNXvYPIWjFGkI+lc1Ug
8zsU03RADSLxPS4nAEt64qXDT3CWp3HmDxVU3YdXdGNT/sRoc6x95Poq7HaoJD5i1CY4YzPmDd2h
FVFgX0m0NeKRRsTtF1WH5eBCfuO5nEU8Y98YzezfNpqT0bi1jUygsl2yBG75C7YfXxmFt6Xd5Rz4
XogwgPj2UkPBctMaiptB98qpnTHxrYlqMXTc3n0KZcDfvsv+4OqaQ0yLNz1LSdMDvisbVCjsSnDx
rUPaoZybVVEpoveOrpRdOXAUeKStmbTr2i+yf9cDXK3rkhiDNHcSSpX80jpGVJlXXOMEz3AiDeLb
WP9PBHJLRYzdI0pj/6FlORot626p6bn52ugfmvR3eawE4GKIvzCUWl2Sr/DTbGVC1wQ1COe1Nes9
S5xGeuBl4w8aC6qWIvdIz6rP7QzYv1318W4kYxgEWgXnXgcaSBifI4NY3/P2IhdNDroJovaz+JX4
mS+66rI8EeRuhJtL3VBpLOmoTobOnLzdG7smqAAWIns62/SaMq/35a4aiIoJJq0wKIfvtvQIcCiI
O4OsmxMX/3UMZltB+lIS5vxNX6I3ujnBvF2tY+9BD+/k3ssd/aVoUZgKJs6WuoCiFx9FUg7T7Abc
1rHfIgB162F/ssJIJMJr59uasE44IkSWHiutO/HoiJ408J942MfG4fb6BABWFTTnqhv6ranO82Hh
AOvCnmfu0j5qxrlyIhcu5qD8JzsekshSiGax1LzWe4XdpzASi+AtQ467mNqf4J4BwXg1G+/LihA9
lQQBjYfjcW2H6MIt+ujf/Xbqy5TETwZ4t2DUrTHKCSzWZdrxhsUkktdwEDWMDYMbiMszwM8O51pd
WnTXhKGpFiNPyWBXlUkY3at/7GcV3WMsVEWfO1KntUfz3gqxDa6PadJnifWtlotet7tEkWqJr9hA
wDGrF7R4UtD8PG9AtNVTOgrHh4uqTTHgO9L0X/lxPTNDIaAJpOblRtcY3TZxv78zsDi4+TLiTdzT
Knv3HWa9kXYt+TnzYjNO4KV/Ou52HWFvszUF1V8QOaOClNetlPYmTMAG13cNq/QAh+nk9ryOblfi
/EXiyDGLfA0pqDn7YvcsZiK1fqe1KQ0TIVqe4bSEu7rCsei+XNpGmM22fg3Csc6iFNiow0N6TeFU
oqg0zWdNQuxIRN6Dh0ONxnITvX0jAc8NYNxNqXiEnuLTbgcVj1fp4oXPMGkOO9ZbZ/CcXrEPgI+/
MU+0vOtqsK7OgsGMGhpcuroeausuuN2sM4yYXibf0sLvQm1vVUCiRzr35CjZ9x1ImK4R/QDwYu3E
qI5fNTyKuIJ2bZGyh+pC6v5lZPNZ6zMSkbH3iWmFIrUhSL7UP0S33Rbien21Zplu6KTMW2u2V+BU
olLONhWayPPt20m1hk2AYB9c0muPArLgerO6J+gx7uySiGhogW+zxTncBMtDnw3JrMxrbezeYn7G
a09JOxlomzl0sn39o1VnpNTRw9hFDcRU7pyzKojSIu5o07rKHgc0Yn5ZF2T+xsOuut9M7Nwqc7SY
xKZG8OxFly+kWS3zFrfJy2IcGfVzRigOH/qOnd2Io+D5eULkgJfbCaYPf0a+wD8pl6BUUipyAwiP
nGfzCXrtRV7hVhxpZJsdVWROiVfQsv3shMicwQyCD8npKwDSCbwIKpua7GcFFMnqZ59yl7S83Kob
vLHTu6BKSGFDKeR9EWYVcccGyWNYuF0au3PMHCcFq+EkJR9C1A/pII+MLiHWmP5483NHccN7vr/U
2QNFhkdJ2bOXUUoBYUeG8v4RESilZ5Gy8efie3SFxea6gyW/0IPaevLVDZHFoecDCz3iVd9XDa2M
5IZD65Q/5Pr5d5C1XWA6IQQcz7LpeTa0+wV5NhYG3WjOQ/4EhfAa+FOYzhaXAEtcEkkxeAFx9giS
YwwFKMWmFLpLqd2tdlaAi0hy8lSoE8Jy7PIzDfBI3SkN3zGVdXtvJwUkZvCyNOwn9Am1Io3OuE8N
rxd/HpmHXqrwAbInZhhhBkU8N2+iJTDloO/eYr1gFpiMCgiiADValQVFfTgAZaOzXUS7jjf03gGC
WZuLSiz5QtH/psuGfjBE++BKALXY5F7RtYnOpyfmkztGrsnh89+RarcKl9XlbsfmDHG4w4YdLiJ/
TFzXml4pmru6byusvN002KRlSz71wQGrYAOqhR472cCqp7QG5F/vJJidYVLdBN1D6Ae23YP8KJBF
XluCiX+zlXuhWI45H/j0Nrw6mFMN8bvgcMd02O/D67SzY04y/Ag89vCx5INqqijqhq3R9Vqeeamc
Rref49D1Eg3lFh3GN+4k7qt8rddjIzeEFngaN88k9hTrRPB9psP7fq3e/bC8JiZauZxjZAvZnatc
jrbReBzMAn04BL1bYdzW1mPG/Ow94IZ2JVU8ZAC4AnR4JkSiX2QOP7qy05QuqJfH7Ge58P4sD5TQ
xzelzs6M8ErjXcxSmuoiD88eib3Bwu1NmQXMlX2a+meHO10NUXcvBt8K5BpSoybu0d2DUhfclzCS
9+4YY0SVJ6ORAL0k+J738UMl+xEggt+HKFd6PS1hEWh03EZX62a3H9Eykj2ydQ3BHydqxqBGDd22
/ETPQRk+QhO//xh0oKam+g24wq4+4Zq4t1Nat1rA9sPfw1esXcE9LRvIol5v8xb2AKHyDyZT/J8R
QNn0nJrGsJuMzm6mp0akDl84gUIAgYDGbx3uJDui0fHJOadcFXDjLh/V3dTZ3xMmkYzocQADcKUU
SzKLMyVW76SmU1bhVuO8/GxOYuB42I78oIjtY+jnAFa/ucM46cWVEMSKegKIA/unRXPAl1ie2N2l
TeGlf/IisOdpllRhPERd0yYM2ebTk9YkYWR+PK4o1NrW3ak5HwvZuwhGTGoHJlqNLnVYZYxOU3+6
Hyeot6C70W5974o6XJILwgbwuTu21w0Wq0Tf2m3uuCupOBEeA2XVrFPZEqPuIyh0ubYFoz4TqT7F
EPofAKPDv3eoBYZOFkLMj42L2PFpaHTQmEX0MzCrm0Fxe+Pcu6bnHevGmzpmfNXqeDXJWdl7+rt3
PAvC5ddxDdECKrFhJWd9vOWxySEekvhqsm4VuMU2NOIFv0OBoU10LffmV3vUZlwE0lSFjdmd6PTV
uVzYF81nuiKtx8QQFy+ZjA5CxwfbpNDA3owpc9dG4pXkpzuNW+4NzTDXsz2cEhi39Hf6AxkMeffX
tlN3qBesyn0JgAuaCKMVCZmR+Tp2uJ6tmG9/3SqjlwJ4MekYVFLfl+cvDoP7iWqbdoaHEDVHxThd
mapvgtDolr/2Qc9BkDrNRDqz3SI6YLb00cCvhyfolBKBUQTCdwkD4bt7zhiPNDgfe9yzJoUjYwVb
VxGKFp97KUOkiEis7eH8OcTDudvMcMJzFDgUZffMbgTgMPZZId0bamuVbtOtCHTstQj96tDtMVzc
k0m7+Tpc1tUA7nteNqFsHb/TcizYwHruyhwMWYJG4/FJ4Ua7tEsDzjd3ZhBGNbO9I+1fbHHBY0TW
rEjIsze+SbRvdt4bMDbCDYdu3LZArhtK6O/BWvB8NSe7tL9AxjIyyJMjv5OpNiAovTdnZJe9I3Xc
WaPJ7gQGpsVcVIHXvntwSCt0bkZtloP2CbHjNsWNqOQCeo/YvaKAq0BENSVr3mo4foit4GPJzkhU
XOG7bdrk4og+QosUOyQeZ/CfCrJ+eW/BA1CFbyjPxwdBNVYt+GtfTA56AzqWl/vdPyUUeEOR58EE
HOGB97dThNNDqYv5+KjAAn8BfZCYtk3Rd/Juz9FD2yMqwsBIyK7pJVxH5c2KdSSBt1VndyNHB9q+
9wInVIybIkBAPTg/pn7UGQPRgb151bXl55bqqSAEJnMEdx7v7eKztXOmEm/yntZurs9ADnLEmAOg
tvLNu7pJ9j4KMMXyQa5ZP46ReiocCnyUxep7o557GkRI/ett+sU4Nzu7KsyOAAGsq0t5vYVDEzda
c/xCT1WMq0/6PElwvh2r3ftKh5soTGo9c3FexsVSCaEOFRU67zZBh6ju+EwTb6QkouwLwOG0LL+O
qKC8G1sDL+ecq5q5H12TYxyTufZ+QldL6oDiMVfbHFku2NJ60o/YLlB5JI2c91Nu7tnoCKlnjghh
+c8LmXckIEj9Syi7CEK1u0Ys2vhfRc3BwPAPYUB2WQ58WpVpzdWmspxoPcfFthLtu+9+m40I0hft
a11a1TBaSaD6TijXWKgovwKScH8+PkLUy1aPULJiF7nE9sux3rn02lvXOSqx61clfOXoF6obVswZ
qNbf5NP97PwX7JyKhwuWfBseh20wqrZmognjx5l5aLHxCgYGoum2izKpDIwY1J34Jay3+eTXanMl
b2fMqgHEQhE/vQSUcDIde37hxu5lb1fwcNOKUKdiYtXtaROsMotnZ4LiRlbW6Br/RlR/UH0iDrQV
ikaKeNqQNMdnRHPAPTaFmRFtsbhfg9Zw1/jFVxnFMBuOvEVx7pGZgrsA9JMJ2KLobPcfDGD+qTtV
QNKuq8TLBQy+vdMXZaWPr7SvpeA2aAp6fn++NX0C+2sSUf9Wag9+Ua+qW8JbFNUZWT03UN+vjT0b
bFaLEh06BQJ7D6j9AluIhM8XApZqAGqsVFuexeIGvPapRAtaovd5Rkmp8XEalPRyRNECKoUDvPQG
jzTTLjYNKil2mG5HD5FuvaFNIo2dZZ/BMRWgk9u6hjTz/NB1JgQMQ6Wb9tIKMgreEKOVugDfYALZ
XVeL99vj69NHOga5If+M37VKUq2hUOuJUqIjGYogRqPs5m5lQkwfrxSx073loPL8yUMiJs1r4dS4
pYt38nmAT6KsBtqhbuIch0Nx14a8qfopBTvsS3gz4HS6TsnbuQ1H1zaxgPOIEruMU9L/Lr+oAsEE
GBjw89C0z3Zw4knkC1RU5oJjS9Y6lQURE38IoCrVhhqDNyX9COzx90GOtqzJSHylJup8/D+yXd6W
yafNl3lMrb3OhSvzGLR7ABaPjJ3CiKfO57kgrj3/cBJaWvlcZVPQTJKi1DAUMDLY8jNLLj+E92ro
AiX7im33r2hxUPcNjQ3BLiRAP/Afg6Fs/T2GQVMIMSHNjRUG8/gaYMxgWOmyoYZ2oh1c08bHlBsq
EOl3hxpBYeLjcIZL4Dwd3HtP+XcC1vMyAN4BbcycqDcsf0MxU2HXnLXfWQ/Sh8Ny6Xyx1BZu+QUo
94xVPtZwdxG/9NqmjahEGI8ydNO51uo5MNlGSRrY8ULCYVfhtUPhpi9CU9c0LvYjX9r9Whdki7e5
HgERXM3B+pM63AK7GPPb1vTXsQFRDQB49EYYFNdNugPFsELNjxNp0aNmCGpxhClDbjMojqNv14gq
UOGPFVJ26nrIC0rpq4hMV2wzmmg2vA3iahkZ9Gp2chk57l90G+ehXvJmMIBYTk243kqkO3E/ABjZ
vM21PLyfFiZoLKQnPcGa0W/xXcjs9kDLsZVHnUFiZk+J03XXGrr3Ze2XP3a6nIgZppsiZNQe95oM
zOd2aZbBOVQ1/iC96R7lDj1YyMqe7XygmAYQzfe18lOdY81oiAVpp6knA1q5JfinBrMrnID90p5C
dlrhULsdCVW37mo/PFc+pzA0OTlZuiJrN/ueCi/NfMUvC0PMtyUpxJZbTTXeJQUjeCZi77M5uz7L
pZpEJcJX9nCMbSC35dSwffQZHH068uUNJAEATKxhDUiaVZrK0pUqgYO1dfQYXHcT0Ex5Z5n9w6ht
0bDZ6vzrvXlJIjLWTmhykIc52+kxtb6rmuJh73YbkFiz5RLaLRexvlrBTOm7HF1OfbtkXP1qJCYW
ewcvPeoAo0ve9VhIjaVIIuyZ8md1hY+JJVhuyY2TSvjJmPMFchekvj9b832leIRY4PbZ4EkUkkZm
6OpYA/5zfii/eHXiOaoyCrx/QpLHaq6t9glRHu/Y/LUOVm+9/FtKKm+ni7HHtwAUGQ2txpeii3/S
pSmJARGF4zLubrsYhWao/28tnmsN9iqzA6J5cYD4BNDjXx6Ao/Hn1aXvFBywouCAl/R2DBQAAgBu
Zrf8wBS01JmDhi3Cpo4jX/buwshB8nTZ3peVkAICfuUUFq6cu3q+YRAM1zI+ErjV1YPLQBsDOo27
Thb6SkIqpqM56manrREsyR3Pv0gtEyMura/Y6jteO0e4U/zxJtp3UEBSsoAtx3T+0PlGv0jbXS76
spbCTJl4Dpu42DLdcKAeZPD3K57547qcCSElSd9ArX/CKcoEReYMyqtfXu2hLeJPRmieqvArv4xI
weuTmybauaGU0yhPq60QxqB9mDuOVSJTO1RuWPMICH3JmloYwfos0Yuyb8IkFqlJoHgnvk/KKlgC
WuJ6fJwnf2XXqBrUNmGavtE6o3Iu5PkYVmo/rTIrIlK5zgC0NEMFrxqPuUTjFDoN3loLgQVcZjLn
/Ea3+4aeWAQDxP04DZDV79Hj8FOOpyos9qMq763Uziq3FZfwIxSWyIzN0N8Jt+oiHK79YJsXXoSt
TpyLKuQ8m9A5yZHKk+yZA4LaiWA7ort/VrLQonALHjOZzJEsLTnTONScgC4OR7E+leUT63uFxzSZ
H9lx4WvPP0uCTr5mHPefQ6l1k8p4eTbU13rJp/osS8bSf8V/CkXhUDIGsYyRmXrFIBHtvLv0Bq8U
ENm43H4XhYFXlqgLPb3IAGmO1wEH90H9qebZSIkhWB4bzcScVWhzzN7+OfptbagySqxs6/OraH7R
iLFyK2o2Vo7PVGNrrIUJIxpsMd9oaK25AtuAnVS3YwIjI7+E/Lg9ID8uxFDHOb7kG6g+a8if2qJ9
cIQwolDHTk7nQOfBnC+Lpfwr3XW3xOiyCpC1EIlD7kxEyxKZw3Tr3g0lgcNOHfAPzD+SftUNogUO
CBtBTNf2JGLu9CiyefIdbz6eYe9bBcfVlL5GHNxRTOCYkO2tyPwL+w9i+I0dtTsMlqV4F0sRNzoK
ENLvcZSY06jMcdCtkKSoPFNQz+DEQARRgw8Su6CmyMnU4FhY/+7Ms4lUbabXZ3rJgBPBQwIC87Sx
+36s1pMwa4tI/JEMLQqOndEsE05SuOM2bp5l2xWNwnDdao1F4kIznc05aBYAL82fAqzWNBj6CA66
Yb4VyfSf0Cq3fpCEnnGvZIW00MZeKX5zadjqunA2Cn6FscO8qtMI1CVkjd6MxVMfVfO0iYZnwn2H
61y5grGxKPdb3BAqyBAKQbJ3YoO0T4VVs2jaGvP290S3GdQi6iYcDQB4DW8Zt6NDg/GNfpDerW7D
kTUQcxyLJXN3rorYD/IrJYRzeWHGLP1Bn3EMC81Xw4srfADcNg7DfztE5UwKiw9MSCqhGMdbltXd
yUt4OaPOrti5TgjB8RzJ3gtTJQVUyJ9ccmfUcWADV0sZDzo/syUVI32iStO/MSpeR/AnvKo0X6vK
xblN/IfczsDpYxUbPRmEdmUCrjJpE6QDP8EUxqYT8dSUA2OPBpTdDuSM65J1CEHOFOn3OMJMAzxF
8e/YrsS3X4fzcfV4V+MEfpJRvW8in+56ez1RIZ9cFqk39I4eJjglGBWhGUyM+mScsVKzk+DtLd+m
tvXRdLZWozMc+78Yljzb6fuvoI4MEDdpadtsklnEI/RwoVa+0n7NatJBHazWrUTBj+FNoJLyOqad
ezQuWPqNLNLPKsmJqKso+ejPSzkCCur1209CCstD88dnCiCy/IDoTajvWLsi7Aw30OCYSxvYwjkI
C9RDPSH/kegdsuuHVLAd5rmFMJAiAraNR51bxKcAqeMWcZ43+BlZQTtkH4IltYqmdLojHq8CmPOl
5tIjd9baz7VE+j3vwGHm5kWenhBlfRMVGL4dEVgiO/M+ebLWC2NVwQwxnC5BxCwg2bVgB8LRN3Mh
awi9bHCpMGdlHrlfpHmASWFnb7x4H1c8Cg8zN8ke5ZNV1gpBrYjuBGdudAK7V5v6T9cHFXfv0Saa
Fg6HlMkbHLIKSCDDNxLvZ355v3kxteEyiADs3oBaLGnvin9kCoiaux+i0Scj1fZ7zn3kLvzbKbmu
A5AdSsR/3GlJy5UI3XRRfLeEgIGAbdx8KLvv7Utswf9mUSyOEK8x2gz0cffuxqqte4MNTeJMV/ha
sp0syTLN9JOSo4rAoL5Vka4eGvlSNFg+s62nQR86bqzLFv19Wlat3wfj361kZVrAINrvMxy8OThj
54YhHHdS8ITpHNKReymthRK2H0Jz+mK5rxfLcW0pGLFKCXaQAVWy5Lm7OponCa0aabBH9hifzJIV
dmDHezAUZ1tZfcnOo5hpiFga9898q7cYl1KvQnpBvm3FtS+4/LFDTFfTvRLY7xvbWDePa6Q52QeP
ZGqsDooDaoMrlbwnofa2NcFfyrrs/xl2ZT3yb/zCX3Bkx3+giLrvsiCyVgCHHg3mzYvOVh8irnTw
Hn/7KtW/XXeMtRAYKwRiMjgYpKD4bCTIJjykQ8a0sdzSV5OKQ7jx0nH8Dhgf3ilNL4gAqBOHFLgQ
X8Zrg4fTvd4RN0ktt5ijUtPU5bD6Y1aaooWgx/SKP1FGM9FHeIboAfMgGWt3Gj1P2LVwBU2uGcw8
qGQyU5pBVyemAz/qn47prWkbde7v07Tj9kz5+xa6JSCRJnhkS+q0NMinj36nM118bVukD9a8mrqN
8wiXqRxCUAfCAyv3ngw0t3+n0Vlsk4EsOGS0SwMp5ccHPg1UGhG5aLqMn5pn9/J3BY+BArP7K76E
EruCWvjAiybJDrbsKooioLXxXypADRxVuep8WTjoFb8tzOV+yTZs1RuGsElT9O/zJtRlZyq16Z/Q
Si5tG8K4szMkDVHYRHBNS/iA9bbr/b0AlOGNZx26wg2do3RJjZdQHSAnieAWVuo4y0Ob++5v7xL+
6Rn6Vvr6UWW5E0ZzcvteP6Rvaah6BsDn3LerSxPGqyP7J4aajhyVOr8cUNEOoAFfTwgozfmNPQfD
FjtQQril2HUHd8lv9IpdGYZA3mKPOFyQ18Bev2dzrNvBpGHQQXPETMc98LIPwhnqZhBwZp7ppvHa
Pt7qXH0WNMJQqjGYSOBX9xl5fS8/c9/0NENEqdgD6m7GiSOVynZfkebzNaaCKb3grbF/7HeulJk6
aD8mKwkxPdudL7pesjPVtG+4C58Z/Im1qRYqAr24UWHimTYpPtoYsZLxiTMgU0ccGwt+TWfVqCbj
guV12vaPEWHXCJPUeYCzAESX2yYPYPSllAD0fwuDBRFSlEyyvdqEhZah9i07UcaSjN/1+BywdSQ5
/7WlpSUKt28Kvtpf1giteGSviTS8wSRtLjMyKF1yoyxXXpUUwY9FEIjFAZkm5kdjCfXiWO8Y0fdz
LKWCxSoOe484LDfV+yy3Uofc/00A+eUYG2aLuJyMwVr01rWpwoo6RkqQgTGxMwim29Ky5zVvSk55
mhQzRi5dTpvKfpTj4OnSrruvZjMCpxeZAKI9rzVwDu6SHPNXRjt3o11s19hXj+dh5V34SKcPTRHJ
SxR/+CYD54amYORjuJkhs0ao8/5DGrJZe4Kvsb5H/4pEW+QSdoz8mJSaow0dEIuanC9PrKrmyoET
9OeWJDRrGvrLMt3czugPvEtOc2/vt1fdUKiTwmoa2E9DNqK58GnYqC3+9IN5RKcgusqW+WZHtiKN
8xH65y7PqC6z/qdgg+UfxXU1suQoZK3jNA/rQIZy/BahWyvjg8paQP1gnrrlgmdP0552HV8Ie4iz
kD8MNtOPiCRKOsBxHxHZPdTYU7Xet+/sJ+DrxVNVjOFQ7Cdbrb+NJL37tDRC2r7f0NPl4yIQNA+r
hl2KaJl+YHf1PN87LdAo9lW1s4gYnGWsMpBoCsxoEGUt9mDF2EIbWxTZMqq5Qd8Q7unehNqBDH+R
CcBz244a6Ea7uAGkLph8cgpUzcBeDSALlTyf9y+Oh/MhkDrBM2YFvZTJYAG5+H1AYsacyg33SE53
zZlb1Oqi6INVY/wjJ1wfMGAqr8CQYROoM1vIdZkPgU6Usij9DA3UgsIXMB2FCiSdgj+prrHdBkPx
xweSydGfGCnlnwubJRxmsWgpOAuuntmoatQJDK6/JoHYZDZm4FS/cDG8f7GZLpvYRwMMHMoE1Ald
V+CpsFUUIRnXd29xM+E0PefoE/5CmNGZGDELsz44WcjGFGgWE4QMMIDqgy6e73Fb0FbPN4klmKoK
w094QdL1/Bb73o/+Q5Ef1O11SRkkX9HG5k0jpvWaxMa50SSCU6gyax/1MLL7G19l9/sUcFA9qhTy
FtfrP0CS72ClKpZGjr9VEfQjEr/9qz1vsd/1k6Sei+78g0kHuR/pVIKX/9QcbTIPamOcLBHY+yEy
AeKm89uRxdNcXOlXDuWd03TzIgEOuJcA3bvh6YVPEEHM1YOiBX5LDwz0N4Ok4nyeBh4b6kD8L88V
E2YJZTEqM5TeednGV2+cq3d1oHP2uDYqMiz5ZOVFH0FNhpTrK2R6q6E6Bulk+sYnyjTIY0mhi5iq
q3MBIHOOYmPTn1QiVIJwKdAv8wq7uK6vyYaMz8ALP6KwqAqU1QpJyN4oepqLChWdrvS+AAOuVAal
asqwfu5y/P/HoKKF97a0WT+uML0F1rU2cg2JoHjrGQNCavk4hZR9kKas+0DYT6ISkJcWS30yf+38
GBrBk9jsSTO297HuinD1pKyYMU++7jpzKBiBw1NV33kmvTE9JbriHxwtLGlECrwUZP6aHavF/2SC
fAvy1saIN1GgWNS+2NhejuopMDUW9KJ0599alJJ533nHf1mwxnlTpE8Lc/Uv4UJPq8cGKNcEqxzr
Ql87g9YzFt+ZsZqmzmmly1j5UQ9ZZRdb+WiZrYx4fSgJx8rIcfoE4OQFE3MT0iLENEi2LmfMB2jB
EofeRBLF/jBY/3c4Xr5Rn+bMBm9f56HM5La6EHGQqLZ+Qe/xjrFCO1WCpxmPhX0VZCTVM8lOqgKx
i1VL0m3I0a8hRo7FZTncOpEVF1M8sv7WIXjnDMCBenII6pi6KT7KoRlLMP5/HeDGC9W294PfwVaB
P7k+frfa+NPoFFmsaMAddwIJ/EpbzKQNmBwQy1DMkVsm9tIy8jsdsqvZpxVvJE5NfvUyAWAsI1h+
D7FmPF29knMXpu+3FefmBVImkNyQED9ru5grmnjJPVCSBHNrft+kcmjjoKCZZfvaE1TvBYqTruxq
2i9x7ekkj6ys4C3pCFy5uATKTfgJguPoUXzub9JuNI/VFQ+6qHW7YLt3umTejuMun3ArXbzq7jk0
sODULir/siMRIyw5SrUmcXl0jpRRg+V9Vk8HLIfu+H8dQleruVVKYrvDoBQPaI68N2kqcI7lzdkh
dWufO7b4FFXBXER/oxX+1TZGzcBEcSSZSotCNSpuKYLd3xnAe36n5IBCVwINwUeNRbVYvFJLh+BD
jT0Ua92sLeW+pKEruYtVenx/m/zEuA8O49kxdQ4CGP+IeCj6PkkPxZh/KfKBvYgvgi9yrXuGALHj
MJXwdmD6NlDase7ilH9oinLYF6Zol3bEUf78GLyU5Wt+Xh1H4/x/0+rLvQeQVPh+5Uw24d2pzzVP
tmUI5ONNwcfyK/QRZDdz4ZoU0laRSF+Y16I24DqxGxcW4qUUQqEICsxH6FGu06FnUvp4iF9ZAwHP
hpODRDgHi54JoDZ+W4iRBP+sD0lNLL+pvuJtPRzdgQMZKrz7V+tht1zeZfFBDfJ5X1wix/voWISk
Qlf8rfQpCUI4+gMmoLdwSGcbthQJzxrbeayzK+w8KU2+oveDV5xucAU6XZZ3krKzlc5h1lvd0C2v
RrTkzPXQ5kEBe6d+YJzTW/Ng+zu+oklT1CEmKPmoxwMkISJzXVbbTVOZGe7k1HduNp/HlNLJPyf7
M4RFPtTub0Mn/WeZn8lb6+f3P/ZB5FnaCWFnBELQKmy2KB63LnGGoIuBH6cDY4TTx0VlokcNO9hO
Yd6buq3iVJlBeyxHZTLtCUD8BGrTvNA2p0Sgi7MbfOTBgrSy4ZsaPy+OHHt5xBGFwHt7ca6tXzhB
3Q6EKpO3tFjnJLjS6jqb85D0LPBpGVa9oPLuGCHNRrYuZcAlv2ywTdkbzszeW5fqI7cUvQCLKJ7e
2m4NSFqnLyk8FLPixjICx22Q13WTcmPmN5K/gtVLZpLT8IWRjDH0qB1Unob73iClOfd0XvyEJteC
iWlyp2dvjY5LLIMAdx8BZBoaybMrzC6d6PIfWjSna5864zJkwK5KwKijhd4iSTVyRrClYM6Nlr+Z
ffq4BKYp80/Kqd9X52HZ2IO1i8z2lm0Qx3vLYQFoXMcmPlN4aBi7xWFbRTOnhFt45shUc6AccJrf
o1U+mBYmvKMgx2tPIrrFsc+DWI315EFbtx9d9L26QIx4EuJnZLU0UVUpKDLYMIK3d/fS3hWi2C3S
dY8rxujX8+k+NGVjVgVdnc9jKYFXRdrC9jIbPEy3A++F6996nhk3nXltAsG9bQu61IEU55KY+gIj
bDWB5W70uND1frPP5lyn56ho0Q41L9E0/v6URd/8Hp3HTlh3R+Pv0BSDH/i4rP5S1Q7eGsyIc31w
8VUKRlkxN2DIkQ5bJmgBnxBnhKDSH6cF6YaoFa5lcH5O2/NtxIE7Ej6gA2xXa3CL5ZJ4kRM0o8pq
Y1Bv5Zq0wzsF8Cc1YDftZJ53AjoLy8EZEs+kIyslcpboZ+ka5FbKW1+bodPY1E8EER0IqxYs02mD
WtwS8S0WXXCxfgVwySaMupMh334QGbSvDVlHjbgIWntYJpFlqE275YBMASUzp+h+6MhdgHWFVf5R
eBn9GOqxVGnsv6RxB/Z0YXXJ9ZSoJpMmQziHBTR5hh5fvlDqu5TjaPJvrZ8WmsE7gw03jCGxmXPV
IX5g5JpCCACPBkq+6zY/Mogn5V5Z5GzJbMw31GQ0gfw0T0EIpLICyt3Ij/RlLS3oO/rHRpgJGOyy
OUQI3zhAW9ZuaO4FF3mXkyhqzFLcs8HTWCIFfqq1B4VYk3VkEhJ2+7NWHoknn5GUJNrPcjDkjTbk
7REXS5Xu9s5YSiBOnRDlAXwKlbuqaEB6Oli/ZPcMuqCfNrun9+wiEkK9hiFmCygriG7t9b1Dl/AI
peOFHvZza2GqaWNnoP+3qucgdhxmvf42IJyhLa3aDFR+XTR21oDEJEaF6QzI+ZJt3zyGlHhMBx8d
dSLl0TgwNzuAXIhkRJsrPfHPr61ls6r680x9a7y3jsyiRHkY8Yg7ks+AB725dFPITXRJO9m1LDsV
2Jg+ig2x7LHmX4r9jUy+ELIx8FMThoXyyVsnCfCz6EzVaQZf3BZbkCiTq1SvGLit4cPIRGLuKXgZ
yXYvI+83lOmnV1Ig8qFg9Qq7eY5E5DnmVUT5Lo0PqjLC/nRywtMiO6djwJ5vjBMMTxwKWJ0cOlE4
XYeOrvYfbWrt0Jcvr69MmYgTnZ6sWXybfThC4+ggUOBeDqWuKToZYhqd+ijMdZezvcErICWSelMd
xHzu+9rW4migUQA9K2cJEYmXsGr8dS/oWUjoAHkVrTwkxUf4IkjINeZAvPX4S0f2AkfDWYw2HdOG
3Lz3lEsbc0MivTQZr7NETuCgbU9JKzEupnFjCBcv8u/NE0eDbq4ovhqV1WTZZS5tPJJjKA/KPkrC
kBra1FDmw84CSojr/4zmT7jNE1uUqU82EqLsrHeyG2GXQ0KW87ajgjPLJQkG8Cih5lKkPj5keTse
99ObKEUH5KehY2TVNY0Tnw2FHegvNwHQRYY/qZ7nwUl4NnqIVHZsVysr6b7x972hydbn3sKAum/e
ku3ZjNLphcKMUwe1JYVj2PAnI2VrBkBQOgC9pACoR/sm/B5nhCWfyTeh0Q2fWZWcwLUrsRSmK0g+
MKJHhbaX3036GPRhw4zXg1BDkTrL0Bs0gZ7ZOPBIW+F9h5CEYe9a90PsxMnAGCJn/WGyj3Smy7G8
JXak+L+X16Kk7xMEdBYL6fJ/BcrkSQHH1ppvXGv6SJLC5qrSwpHTHmxM0qOPXJNf+TYR/TtT0yk5
H7lhAFf1o+92UGhiuAooa2kBg3qCdiNiGRTULhKcmCx1o4OyfxwENVXCYR6WmdFZ6CHWAgymr+Y4
6m57EyUNTT5qpfrjgJD8Mqyw8iVaVcnXlScopzqmRYgevV81PlljcUZs4hNI3JyzXlBMa5c7nzX9
q3OIRdAuTaPYLn+20LtQwdLuVxb10AkN4+1aDeq8K0UefXV5eAT2sv6DQD+v+TOxvZyD1ZgenM7L
Ruy+kA8WUJhDAvcobWo71sfJ6eHy901hJJrdLv7YiRzz2TWiPBMN0IKvXOqJwMhWDTfbck0EVBta
XMRfB1pZqF9vJCWK/MQWv1kL5ptS8OMKl3QUDXxRJB7HUmL7RmSYPRx+7Pnv9OpnbcmLIJwuKPPf
CvHCV0Lx4MhOOOJxnVs7bZNkq4OkRACfiI0tkTzjbz9T87zvfeZVQt1vY6GjDMuCBM9eN6bkblsY
woeKeuFpZj1r90ZNM0JFE12xryT81RZDLvljpCVU58ODEv09+1SlYnda4CjT+Df0ZO/6VWmPyyKT
LpyhS6W/eU0jFRP2q83pds4DRI6X0m7hsPbB8/K+9H2hZjpNZuPluho8L5+JiMDzDEIni7egcJM6
N8n/DfjR3rLrTrcWjTIr/N3np31z25ZrXfrO8G7mmDRb8m9D8BSRevv/vhWMqGZsfQsEPuAdrKnJ
PSeORyaFUmlmGkRL2Re8IZG7wA69NF4GJaY6zXDEj0EiB6pMHXUVQcx41+ZcIvYdkc90yZiMH+wk
KrqxetAejNJBOrCe+yDuZKZpy6J0Mo1BK2EHraadlajelF5eabl481VXvxeKcXT2kaQ8oOEVOBSd
RpJH4mpPZWLPf/P1DcT62dxcJWlNJfw8R7t0lhuTg6Jl04fxqBvvYj7xJ2gjIBEEHEmOi+ubkDjh
u+FJYrlQYSt+2GfxkRZO/08wXZexmLLa9Clyq5iUOve4/wDQBiaaEucRcdmBnNxS8S3zHsTmD8q4
s340dnFHHpclD3WYvFzFnNvWh3/cVgwpSiHuQHJtJlI5vd+RQ/1cao9Yuaqq3o+/1drU5H7kjRuH
l4eHE31eTxXxfRuLhsLIk3tOMmXgr5kVxRCowha8RazAaNVap7XqRaDEWFjkPb8d/r20rrs0Bjxm
jW+sQbuBkZUE9hHq9gyQeCeXOQtwy0leIebksd+FJVBlbC2jhm9k0APAmrBjeryiiWIUWlHX65ur
Hn+Ep46y0BhEHxlQ5BbNhBa3It0h2HGJpZC8A2oh2bvsvAO0BSFfg4mu5EP+w3BNXR7rzmSkT+KE
1VsU1VnJGXWXEpzTUmKWMy1tKtKvRO/cE7FDx2fAYU8HnpDZoCTaLaS/0Joq4wvdqYrddnVMKfSA
ZARFwhxWA2duJAnTBVNQsLZmvJyVG4ew074Vms5UmwrNqz1MvnyELXPj6PHiTvqYSdhRCOHu1HLL
rWu8E8LA/t/5Mbyr0ON6gPG0JW8YZghqumdW9y9r777s0e1/o0BA/HLGfbBLglorXf7aSbhHIMyK
XtZcNXbzn2pnVTPvYEjgDTpI0Ih5vLrPeoJTSvxMY/Xs4B2eWpiNchvrfEDeBISJZK4I5fNh0QWI
CidnDJnXUORsNEbAAid+xwFKLGW5eqrNIhhFq+4X7PEy3wdrjqrmkaojXFySmq7yiHKapzstgraz
EyxpDUiXZSeuJyEyKZQjslYIysOY2vqnDoyqF0g8CqDG5osdmIDDINbCNhQYIFUXq8/qbFJq1ecv
ZuG9Z23KrwW9xsHXSYSr6a/nqxCRRmY0PRYkfGPv4yIswbjY/DDoCgQ7fxNCjgj7TNo0GZ74yftw
z8vzYDqgZZR7Mujk2xKnvmr+ORRApr3RubUuK9AHSZToTC1DLP5ul9Pz5xBxq9Ug/CO3EeNW+P2b
N+MdmYRxeApp5OfkxuKETs2l5ms00UtpVNsj8gkw5J6Y+iGZokBmvfCUUV6SBi82QhGRv198QZcD
aOEe/4/jeVIJHLcqC5jHy5dzfCWrM5RLUphocnxhk8ZNns5Q5BXkAEdE2eP7fPPO+7ujnLza6pCV
TZS917wzaRZY2Mp8qQ/nUmOmaEzTm+8Syodu8KWpnd0c21bPYGtpu42eyVxWSy3SEtYuQfRWOkFI
WPVmOyZzqXhDtPaxCd1jzAd1cDdH+S8iuV1dibbXffRgScV0PCfW7ow6wqGiMF0svOqHXC/Apfrt
SV7ZlkTmfkSA9Gq9tpJgpSa5qlq/xrpA3yHik3x05QW9qy6ZH2gVmUpkSE5FaymyD/bYGpmPXXZt
dHPDR3O9m9U2zN5QmVF3l9OTfM/iZzs9cs9mP09sdJ2thnQgp/4M3IxNkFaQdyyi1q4AVDemEIsi
YhvQGV5LL0x++WqeUsmoO9IxX6Ay5ct1gWdeerTN1mvFqUJvxRKMnPLYEkCDRfhipKiaeuEvsK+7
btgov4Q6IUTA3p1AA4HwOWyhikfyRB7ZnD0LHha6IUGjP81DsNAuKMvW8WZEz9qfA1asYHVmugqd
Vb3qd0vhuxmkqEEEQrIc7e0hxGBMRZBTJCUdBtzIoRJ68cDhr5qVikoyOBRIjCqVolJLOT9cyPN+
mH6ajAIgGdlGFUJJfzMn4pA0CaGnbyNjFiCRuURdAEGf3pxaf1QjiHOaPfDXs1NiybMQAt8fiuBs
xOqIk7gFClkB7eNdpy0xtU7Fb+tnKHTDtYTQX8RYRHsNbf8F7k0B7AfWT0qk5W1wYgxWDO6bGWuJ
VV19+HCwCy57zIyL5v7WmbR9E28d0xaRqOJkOSaqdj5lA2vNsazj93az7N+KLJTAm4xYLKk1Wa+8
Np6WmboJ+I41uUxEW028syvCTsSnX8tABYMhYn5SyQhTHA/qKpR7nrYSBkIVbhKJRkvNS8yoXrUZ
uiQOY1wIbQbOVmdrUvAbuf20HeiAOmWExY4LQWuYzWHAsRVNxEgXwxP3TvsHysUu+Z2HqV45q4yl
nM/wvWNit3Ygvn2v5J4RUe40SbC4X4CGxkalNkAcfYBGAis3hxiY+7Sh5yXILsKbyeA3lJ50nfqm
0bxnxff/SFMvA1VrYVh8E5GxZx1DBPEe0lVd6zMwqPzzWBbPLhExFYMm5ZEa4p5Myuv79up0S6pG
tZVuDAyL04ay/xK76hX6zMTSn2WBzC94UgPtQ9YCzcA38gJpYXlCpTB1I0WO6pSgeRROXTMBzz71
68Ol3S+Iy0s8Q4V7mvEE1Lpvv06tHdDnRW9odGLqUd+45mbHQrpqxY9zgio/r21uPYNh5RIy5RNe
nlugJysAPNkJgo0aKSJ21IZ3lUSklRIobrLONBo1NvkL4J2y20He/S///lNrnihzMMZRgFtA8jGA
2NB0gFK5KVM16CTCDTElw2qtTQg9kUlAA+aOyp+OQxRJASmnG6cI1SnVykpWkxixXmKYhJJZG1JO
TKeET6B0MZmynTMzguKToOkOyoMJBj6YCSPTRjapgEUsV9WkM9sXqp6ccT3642MvC5iYfuwC/q2t
TFvn/07SwN/wNs/FNfmiE8mu7FGh+qudb+DfTY0XFQruYErkOcHHXvW2Mh0n1PWOE9+dc5II7Uh0
WIIHrIlOdzybbI5+G8bgpIq6LaarUME19+VvAbeGxfWbG8iLetA/hEjyjFB1h3d9qsULbdKfngJ7
KuNi9AWSR58BxQ4WYygJZwDqJ0Q9OVFYvskzwG23YEuFSGHYW/cGidMPxjGScA2L+bxQcKZvQATu
L95nEjh1IFeX//NGyhDSBSpWeqxaktE5xu+4j588Ipxn1sTbd6b4CqiBvTgmW8EYJYOkAf5y28Va
TIHpPNBHQ9uYVwQKiyZcK+P5JpdjnRJFZCK0cCmCVe8Bp9tWK4oTe3wc+HTFkYm/MQ20jgj9WCEv
kcvI0DkkRPifJmgkx+a1wg25v9ahdCKTsiJwWa1U1UdccbS4nzKN4fbPHeF2dS5W3A+2OBDj+0vq
GCr9o4BN+8KhWNW3zludnDAN8szOjpMnkXkjinGBvtCD0ZaQdNoF7AcoRbevTjBelFYLpweq/yRp
RdG6E/PyxVRKuPK+pBvg/BFZe0ovj+4YgYTDO/J8Vn1M/82wTlhj8QTg5hP9Y8vjyBJ5vD18lYew
fGI3iSwgMde4aZ2M/bcsF5+xJjgfoETQz19PVvWQ010q76vhhAKYhiGR0KFuJSRgy7foQbi4S8iq
qf1KFxYbRNtro9t3ufgHx76tOX/vRmzKIfNLTW7zpRS4HdeXuVVHYGPZabPPpaz64h5JTa0tzfxo
7DmeAai0Y8q87zaLKGaD6HEZPSJtB+oy9ylxYFPM+0pJHncG6Xw55b1uNHS0gvP6kSpmOxGDjJBa
EagshajuP0SvazNex+mEAJfJmAbqDoTNk840uA0pjByEazMLPOUapOUVQ5IMyvh/q0+aaa6f2Hgk
8m8qZGvrC16yDeutcdxaQQvYmOzZvJqMZriq4JNVQJkA9z6nzTr2czYfT9n+jEplL8oQQbQVe2k4
M6ciTqVjdmKA2bLhhXGa2aofcV1KGJb0HOKxCZaACrmXR+ejO4gHNflDp/hg0Y5zY4F4NqANPU5n
hgQjYnua/yFGaIcLoV91t0l7um8MlUWgBnVeTmMoVCGWmBhkXKOme6gkdY6P/7iHLT4aF3zoeKLK
F9kBJp5xCUemSxVXEomgHaPDlWI7OKgCXyN4ORo9UQAEooLkdNRRec2mDGEYy6Tk2EW6LPgEx7HX
U38q2DfcbaMNs1vsXDIfQ/aLlI31TkjWcmv/XFHf4tip2GQCb+HmIs4alWUH6ymJF1+w8mZiDD53
9ZJ9iB4VlgkTjkUa4oRk2dsIIuaw2WPMIQVJ+neO0MQPhsGFPdhIBLZJUMdDgp3U02AlIKuxTk7K
kHYCUH7ZTuPM3gYXQcQ4MBFrVvTnC7gvEkk939+78XUyv45Rjp5VPILdCWVDJDPeUhbmuCkb4Z1I
kUPyslgLJ1kqvyPvc3y52Kf8103KQ0ag6emWrTAVfF5GA7I8I7gR6nxXGpg/JHfPf+KVT17e6614
dCkZVLevOs13VMPRiu2vrxeLYnLzSM3GsFX5L1PC0kk98UfcKCnmSP2sHEeEkS3EkHPssgRgTSt2
dctD1c2hRPhx0H80hCn+23JlbJLro/qWhO8yHtUGyysYniEuI6sfJ4WgbVQGLx7cMAOwin/qvNzO
Evd08lcQyYJa6JUv1BjYOzuXfyMqAlqWIBZHDGrF02mbAx82d6YJyrnYbFXmpImZ4PdCpkBFU17+
VLf8+lwoqMdS5GzlpMRmPhZpSThPAnGaDawIwmacHbk+c5KXkK0B8LUM4gaiF/6ZxreNacobTHeX
q6gMWJakaBc6Suty3iuB6MPh53XjllUpX2Wd0aet5XtEDSAvB7sdhzUkclJtcUNCz13pYsaHwLJw
Q6S7+NXYHmsQgBLHhm0EGLDtoC1Dy+Oga0WoVN1ihrgrTrHOUycfDARzbLKHNIS5MqYGPBujq8dX
vs4CHnDA5Guj9Znfs+Wg+A7UQb3/EXR5A+McDpvqwpA6pMHxeJ+do2Ak+mJzZ3d2N4IeLChqkLQ0
tIKHecPovrbnmz8SNNXIPBshiwj1qAgG9/jjyn4YFGJfPgj+B9/NJmYIR8bDqYNcYCfa/1ogtZ4L
xjIuU/2GHF0G4BwY++tvEuA9kSm3zVXfy/o8ktN1Y1zVOxEML5bqmOaex8h0FcEaLVqr0k8NQ+X/
BU/jtq0t3b9ixixl1bab3dU9Gec/OhOe1eVdf9DnUeLB5bkpVYFIYRsPqYGmOOT65t85AUYIglX/
hiYxy98PEAeCRAx385g4NkwqhKkr14k1f5V3fPadjdk2hWRTXgFfJDIak3dwIK/O7RZTW3+iZXRs
nwm/uh72Hwn4tZc2CESrwMApp091qJ1GJB/ky4L1zmeACpMEArHVhAOqTCr9JXyQZj5hYQicPZai
fepxVVmwyuqJhi6yOUH5efggBIPfcHg1UPG6t5ph5IXkow46D6mnenfN33hRA8UjhxvvYHhPr8cJ
3XiA77kre0jqmZ/MLeuVrC1HTFrevLbWSA2yg3cShBx4xBy7vCqL5TNnZakSX4aBRfHJsiOkYoDd
SXTldf15b/GhYhhIYUH/OEJkbd8D31Bgn45ijbE8dYbQr0tOfw2RmSk+7gnJS3rb5yw/kSVk0ps7
wK0YCUZrkoMsjYv2dUBR+PGJao5yofUghlZv2Xvfse/JkcbL8VJmmhZ/xhnUrn4tAyrKMq3ijBFV
hQNaCRdTkea6uNgQ8igOQrpqFXrQf4y7RuPbrl7Ixa4nozfvbx14nn7I/x0PdOqyCMR6JKkq7Gwk
j0sP9qCfGZHy0SXJHoCrwp1RAKYOjh1qWXJEC2NoRmZj8u+Us3KY1pzZ6arxuWFD/9PdKyMv6ylG
xUT7UHsJT202XKFmQXUHwx2RR2X9v3p1NtSBX7Lv+pxcSKo3fsYtIowSrIB4AAHEjfI8dmSt2LRX
S74Gcnf05QP0VSar2KShGwW4D8Km6sTxBJeJc4v+pQUCE4VorlWQGzGpLs0lH+xIpwchujdjje1d
EQ8Aj2lDz0oV1WV7BkXn3TzWUWoOOOcCCpiTVfxdmnt4A6nfO5ZwDlZg7s/BRhqe9Ok5r05GVCHu
QsLwf540ULiGv1RKD236CoQ7BrU08NZOR5TVx5LN4NKmy0jWbWxpnw5eXsjhbX0TrJQJVGJtxy9n
J2qFpIpumTWQpQa+SDv/HVZq8yUEhyfMV6YQMbTu0oBXBzgT0g84OX5KWaQJOF19IaXipM1meiFx
rB23MG5plv5/2f6X3P08q6AiCKUEb6yTCg9YRlDUESPIQqkqO/HmXatFjpyf+S4mBvpD+7i/nMeU
VoeehmY/5y9Hp3A9vtdWYwy+L5UEwMsQ+F4OkRaVXHeLvM8s4Z6u7f64P0cqVaON/y/GQ8udSDr6
qMM1r15S/t/dQzAg9NEWtIicnxSyyf0OJtGeWJpO86hYQsqthHdznKwcD1k7Fc2IsuWsXhgdSROd
z7CXuadF8JWKOuR7TDrHUvLV7XMwvZP+oGNZTfpN5P9fIxnP9MrzdaJjiaQqzSnh1DS5hqAc5Ip8
t8oemR0W/T2oRQ7eOWcewBsNWKmGRs4zXjXpMtq40cBlaqbTAveeSTT5w3N1nC5Urx5um1sMsA4h
jiwV7onhUaL/jhAPVCxBXoOWIT89jqOHhxT1xZ4Vi085xUUxwUdP45PxTDxU4Gm5yfLmYXAoZAup
n6poFKM4C1CqL00IWTH5IfGGKAZ7BU6E+xX+vmATM9I425z+qaQHve3DgV9zRg8j0ymR4JRU0Vby
JheyzFHGu2UL5fhElHwtI+ZO+sd/8x679XoF3nOEc7QULT+KnwEi3wRY5FhTyMtRQQaIk08ekOJE
OFFr3E1o02msMp2hpS2HZw3l92oZ8kn+WDa8hTABm7E/5bExFtppV7kiz4mvEr8F8nlBn4oiH1P1
RNWyO15Z4VrQFYJBQkyNHlx9SkJNWwNK+jEazgk9f9kdYFJpsmok84qFgzfFEMc0cQ5mc5Yc9LYO
gOXIdJAG5D08WPpWEC/HrRyzfML412jmkM+kApNUWT48RskQrRiYj9H9CQinReS2Lvrkw5mV5vzL
VLFsw9KDyfmoIVmu8oJ8lEqme0gkzd1VWKsMk0JlMsS6gHJoWq/gnqa9aDJsgiEvXyZEERcBtYkZ
3hvOl8nlObSpjRGJJTazhEWe9dhjBe2v7ziSzOaxNcuhb5RsuLhvRI0vnoyAww4XAYbauFdyduhf
0gg0VyAkWyh/SzvlvvrfsZn7YSUlvllD/FfzuEaOs3oLzt5P7mRnZ3yAV6K99mE65U67I29wUzWL
o9ITiuz6/Sppv5bbAdJ72JjpXLKKXv9UgHno990FdwiN48lFyalVp9p1TQ3Yy1T6DGNZkprS/hjW
N8Qq9PXOuT4zTf0hzhrZpQYkMiDafeq75GZ7XCbsfjvZPbanjLYZq6+aurXsOQQJF6gG9R8HS5h/
TX3B7sKHBZtQrisLwiHGKodBZS2h8rWCC3X9uRmBdX5YJ49mROsHl141nM/aJ+IczJe1NpVTBX9N
+LDljgTWipqYFUYBPjevpuvnxgq1wm3Pu9VJzQLB3ti8KDNnIoRX3DwkuN0utLEjWLxaGrM4lfw1
DGMMMEkB5EJqKobyEjoxV7nE+SMoTSSW5GBg7BxDWM6HG0PQsR34bvoBl5GP6HA82B0OG/6/zoKI
SMJtsYkqAdYRHx6fgvOwdpwqdgQYgUw4UYblrVWjibN/cYufcUQYPCw2A7e09gRfKWG0swU1jBFJ
J8G7iq+qM9ezdF1aHdiLg0jkVIiVbq8ia4+ErQ54zK2Rf+kgHtQsgec/FRbQCguwMejrFQZvSHGu
8/OwCZ4TsWBL2eJ4vWBusMs1slRjyySBG5/m16HWOYuG5kdn9mViPw1su0Btgho3klDm4WLBzjY1
V4Id137SzCTTdZgKaUQrQiGtSMcgPYkB/ZJ9/7LMOMKtLGYsFCppphguzsEE8DSmeJWYwTJ/0fkH
w9gBDWvWJdN+ETNnfd8Sluyc4ldgBfCtfnNz2yVlI+Oqmk8rXWhvMvQYgqXdJMFK6VUoFO5y6+3o
F8btXsYY+AR20jEo659UfTiJ/OQkGwDfiDwx6lgdK8K98Q71YSyvwnlDuH8YEQ1Zni5h3zHBk4zY
jW1oaUB+5e/hY89+VVvJUXx0fGdnRsAFAkE+I4l6Pb8vOqiHUflXLBw9dYhpaPwq+KaqZJe+MdYR
/1DvfUC7/RUfrjUpQohlkl/ZSJw2WnEvhtgYgbz5e3F1tKUBk0nBBeMIGDU9rlrtGdiM+1Hb5mns
VLUa059Oe5/ymkCdN7KbpUx6vQf7LgX5jvIObICJynQWUn/4ZA2YvD7+Rhd4fM8YVQiAjhEhTWt8
AKfR+wuLMP7+kx3RzxpnspEUthG+F0MB6bx1MaYAz/BQEKTTqhLqs9aGebAhhiMtlSUS31HdjQHC
oZFBN3+kWT3y4kKQpFF55KhBjjIt6IcjkZfHvXWKMnvAnStLcizewnxHC++JGorKxxwBagJhWMeh
Yx7Z0eYajk2EUx0jDpzuePC0zjGkCEWCjtPSdagosw5B2LvG8jBjUuaGJQGQ0T6CjWP8aPDeIkAG
HHnxtvR5PLc4t+Quq5R+V3KN8qpf10pcsg9KKZmJtilB6Mvr6izSLORzizdinQPKxVpgarbwDGy8
LmUeS3W1FB+54RdlF6cPvLW8o2LpmchBJXdTQ5+hXVV+06N6Y+hCbi41RslitZJtWHeSkpfZ+Hs1
UrtUju6fK6WKMnUjPN4zgHBYTKxC+PFwpq4kpeivv89f+UrT7d9JvhKZzdW87NWq3qpLwdEYi0Zi
36zB7ikKTS7BBO1unkV42tQJCQl6GPpIzye0HPgPXMyGM9MFWHG7cGJzYYm32sblC7dBGcmiIPus
uKnDGzj++1pkEGr2xlHh1N3abwimcjtGcH5Xa0G52/QPCeVUgs/pvX6KqqXZpfLgn/MfGapl46C/
pHU0PTdhOMLrQH9FR7SbafXQJ4snVKjFLzxWKIacGBEvn1HpaVXLQUuqvYUGu3nWVYPNP7Lh33LS
MMqCdeUxoqPEAmtDucYFtyL11/0UebO8E/0RiBN16pGBloSw9whJwYJ0eNQ3xswWIFIa+VKNW6gR
VohaChomltx22uTmN+80hh3367RfMdGaSzksGUkZt2RPFYTjbebZ0Hl9ASho6LHCEvzoTzmDm6Ci
yxZ8z6GKhgnci1twEJ4TOIOxw+J7rVnFWhlKM3DaDCOZxlx9cKJU2uVI4IaXPSLHXSuKAHQkOBQz
kpL8h66fmhqJ3Yrhw9ZxIQyXFLWvgNmMbGP1tszJmtLlaq0CgtbSAG1V3/Ik4v2Sw1aKIfszY7L4
0AEDzRdw11OJF/IE+gOXXHWiWHqEuZfI69Ga+1gPTknWMy1vfxtWvDL2eENPo/qASkKHljBUaoYl
etSOLHhYbABaWSIUbXDYWPxICMEs96ezYLa7X9wwMNPN9TnOt7NiYcUED3FtHtL61SOyXhWvuI2x
PpZX4RRbxAGW8NcypBscQUqAEKh/mUI71iyRnXDZVtKNRiSvIq+AQm7BRKhzpxcl9xf4gFY/F3kD
2GTqToFvvHx1ccbwS+s1AzzOSmxjKmKizQaA2J+y4HXp22miPSaTVa+moiOM0MGj/bi/unj5KLXC
J2llQMMgrbVV+KxnRSDrjzjeki02nfFDTO7qaXboHnG5ecV1XIdftGJMnUkb0+X92RZxqozmM92X
R6zk+nqfW4JnPjiDFmlrSTjyK2V9HdRqcVv6oWgGKVIDoJcK7EaqOnfuEzwRbT9KdSfbgZT/d4Ph
IV0z6WQ+82mWkLo3jUj6NobetEwkDs0o/W1Lntfki6kCjRAfBX0ZvcE+sTX9Q+xWIHT0nb/0oiB3
YrmxFE5sFw0nln8k2jiYFSyBydgsCHOnaYH2e+Kkgu02KYcb6k3/u8YTdvoipuBvNyn9gI/Q5f/X
thrx95+9cq93dBobkgzaW3zI3JzD/M1247TPmlrBJyWOD5S1FCuJ/j1zGm0E7wg5iv9wyOzH+OIF
wFRjmDPDyLZMl7e+Ydlr3rIrjek4JS4j5iB09yTKTb6RJ6cTO9qXKuQhj1D/OTttjbWMkv+VX5aC
PBMe/sP41Uqm2u4Tia2S/EUGKVu5gGuWJIzfZPOZYach/W7nwLSwVm3AZNfKBWWgfsaftjkw3AW+
Cb5zyFgwWar+pn25Y2t4OivBtggTwWnqDlgjUSi00qQ6/P2MDa4VUeT1H/o/Nxl+0gI2s6yJoz1g
HMvzVSlnlVFJyWdPo2g5qjnd6vy1O5BfABXTqhyp2Ctm8kQIsuPcHiXe5rXhoI34cm/RYEYXqaZV
BUJJsdkCHszkuXyJspIFmHK9oPDLzVP9o4q4RZ8z1ecDWevoxPHcduXExf7Jen8Sym5AmO8bfL5c
vV7KFwjmJmBSIfNEhp3bczPXTUd6Ys/GyDg96GFQ+/XGTrYMRirxtKeEjBoA7Sw/npg187wGp+X+
RjLrLJD9nB6PfPerFhmPxWTutEgm2GHyDoLMu+3JBM2Q2plXvxViR0wt1nFUwDuXbdFb1wMCWg1b
N18iVbaLqdd/jymRLXQx662QrSepdtNSnhTm8KlaI0eQQfn3XmKgfsHjn9cPsJ77WCRXfqEvUuQ4
IhXCp96rTZPlm5PHA9mlFdlF/a7v7TN6cl1xNVqFnGqG7l1IrBpf/VUWMSpo6LSwlGSRKhBoZqM4
EOWzvVRnGf8eetfmNMI8wqvlfAucx1SE3fsXXtyKVzzaxwova3aEiEtik/H//11XPmF+lPef8Jz9
jvfOHZabb8HGzglcfd9JohH5bJG1CtmQWo6ayLGF15uLb02RjBi6M1dXt5NsaXtwE/1VYXffSnry
KngYXqKPGCk2rHDHiEmnOOasEccWZ/F3SSoVTx12++h/+ViXi0RICb0cLb4OBT/zSR/pQtP6GL0h
Yhb7L3+odTZHTOTulQr6JncsYvylDmcnjcof3ulrtVSmZTvVEEJcc56wfgjjrR374L8Byfcr3CiY
oIXG8ZIbQAD9jeVU00STwPaejcvhPYBbkojzj3k3/11cwrsgYTbTPb8qgF6rUXSsS6PDkhIH2F/T
+czSb8/u62Y34FZwU0tsxQuBitoixAahxQnC0O+9PkobX8RRE2IfC28BsAhDcQdJRclWRbp15+Hl
jywbu6MkB0I8fvAllHxWzjIM00PDrgh/u3rsfO3ZjzyrzGwNCh8lDJId6EmMyGAveysoUoOo0S9+
bY71kHwVSzRtRe18dCikvwVe2ZIGk50HQWIUi/W00sJ06SezuTiwxGy4eV2ZVDBaj66k4osZ65nK
8lWLYnKPYiuzxoRl8mLEKTvKBdcQTKTKSMpkb4w0Qc+neeqr4mgiRSaveEVbwgxEhiGGlyr/3rtm
2staf/nufIxUKYeEluV84oKOiypz/U8BEgydom/nbLuCejMnkd1MU12DCQmgYgLrc4RFrKThOwNN
AT6w/G/qSBg0eEh8kI1VErzg4NldYlOst9s64OZYqy7cLDcdsMGE2lusuNuZW4f0wYq4tRiatRUv
ZUIRr8Eh532GSCMAJzpUZ+UQ1G85ltk3z2XnDBPBc1FhBkfcu6A2LbGuuCzGlG6JkTcUs7ThsC+F
DTohvI7rnTxR0AOq1R87U54oW9ukAkixvvPgqFO1kfRgsVoHnzZb16DNWSOkaaLXpBKFrP9h42Gw
tPFUqbB26QSmzJeQObzi+gFLcrJFjO93jDUAfao0Bcthar7+ujdYNoX6Qrc2qchNsWjGgL4ftxer
RdaTcNuMDzHLSv7e+VyR1vQYDkJKvlGg+A3FVkSiAIOtKZVDHu8J11GEDrr7D7pg5MSDS0hbJHAC
se3w/Dk5U2FN7kZU4uLWXgD3Pxz85/Eh1qulwGt7gXaYrudjMsNH9eO1vsW1AyqLohhA7go4In+J
PFW2UwYDzFbzQ/MNiM+HmeJyEevMWgSCuIFkSU2CH6rEH9bntlyFAjXRF3tjrvprJk8ISLLD2zbG
8+n65h8mc+JcGtYmEoogZ1mJHqIQ8yqRDVAMancW5LBf01EYmDwNeh8ZHEebsXGx78MrqJ7+0AJ4
Y5fT/nTe91jsKsNbZQVpYVbIqQvTu0XdgjzRjdZRxDhJjJzLemRw82JxIN+AQDK696qUBmCcn8SS
+0al2WvKGPhj4vxdSY6IWlUp1f9y+AbqNnXxRII9Wrxn0FdxIedFjUFXCY2HBe+sx789J4Lc4XN+
uMtnX+csqtLd8INL604ftHpsYoqkzcgZqJPP0sxBjxF4QP/Mki1ugwHjAUdm4SJhPextblVdY0hq
QWww/NA2B3xomWk3iT09nNXJMzHIj5McJvSsjdaYPcK9QrheU9uvPMpTbFOhJI2BtJdYX2upV2C5
2NNQ37VJ97iX4CUt1/+R+alCuMVUrt5D5U/epXn+u9xafHyvF9/Vk61joc+IBC5IO1L81HZFLypN
XS5BtkZg38piHaA8PeJpeUYzxLxKGMX+kHfTJJNHGj8FdKOEpaHa8PqbBjp/XNDQ2YQGjVPGM0K5
hdVzRotALgnpqMdnalZ2SJKgJhb79fD4x6dQPP6+2yX2R2Glj41MeIPCV/2EJnR/HRS8DvYocilW
vYO2W7Vhb8t8lAoiKCP7WEJKxTU1ehIC2ikEUmDAl7mIHhboZKUPsoqHmfnjFEGjAD+ad5Sbanax
Q86JZv6Vi98uSBEW58YD60hv29MGxLfx3agJzw43qn3rO1TsvCQvOt/bZR+cKUWNzt0DRs5+yb1/
CDmKUMWgO3F0px5Lh22znOOA21UkUCklFA73UdMz0AA9CYxCU0Y+w11olthWtvuH+ovFRzudRWiv
eSleeHVngCv/ySH0jegwbL7CgkwMrPx2pY6xdd1V9WmPtLOCP2503ETzKx8uP0xABduEzcara1Pm
zBEfbx6sSMFvoc0KMEIMFaxDP8tkumDG4zdu0B7TBSHlPrU5JZl5ttfSlkzjd6x/MWYUaVkiuPyJ
cmqCU5nNxdVSf3Zk/HRrhc54nJDLeqGMyfUNe/uOicipWKcI2ZX9gDuGCConqvpqG2gnQFpc5IG/
p51yS0GXiawLAlGx64gmOIVqTTJkn0RNXRc2ADLShWYjw7R8oAXkN6bfKBEc3OWx2REN6JhaWO1Y
znLXwob+5YYZReXdwyrSuyNwRiVdNsrNf1IdewfUEOGTLCobHk46qQJ/ePPuk7qW6sQMsvZIwv6u
DOCxqSgPo7qsmaZBGSQNLfSHQlAFQEN5AdbKAniz6bQ77MEWlzhC2b2mKGFjcVWO+ZHvQAddcHiU
tixi4jm9RnTu+MMe5b5eUKs947l9vgGOnlK20r6P68jeFyWBKVXobQExbBGu/KgC5uLk17Z1ZpcO
KI5qYI+KP/tkLTa/OoE9cS9tUXQatP5maJwPGmKWJx5bA3kIUx4YBJEgwBhOBIuPOx1o/T9M7lyH
8r4MROb9kexwnSJY4Cx1NyLa2ts5pRHF3MVvsLuqZKLzoXKUjwZu0FKqvffSD3FyxiXCgdTO/mTL
bt+74eF+KAaZT6tSBsVlXOnKFz9IUvsgoNxzdJCmALjkHs5/byctwkimcj0BXK1x+KO4poXgzpW8
6sdiAfRvsTKICIdE3HZxeBE8aR51/TrbTyE6tAm+4NDjEeci2ODaPzahkz7ZIek8OYhuIz2BKl2V
pHnllVm33NX5rplgXm4369yNimHEXLW7Cykhgazb1rEmtTnw0H7BztiP2QcN4uW51KSJhOyCkCz+
xO7qKYTqSv/uQmyAQ0lcZNijXPBUtHKqwfdNgKbVAtq57C/NJcQsIJXEslHxPlKXhF3Zylsiif6K
9ZJL9o2oW5YrrtwXNmVzs2zfZ+NomUt/girp8ohMl1gEyPIjwf5RVpUM8gigdaciuYPA/mltxiso
gdQo5ge3TRtV7Sru2ngY52AdkJfyEhTiPiIrEuQBREgPcmGGPaQDAAFOzRAxHMwBj79GOUD/Vqhx
JdmZ8YlwamsUMa6UzaSprf0eIsezJohNFGWM6WYk5Z3iWhXFZYCeaBXAb4PfmfevKmtvD8J4oLXg
tsmCTy74urWB9iHs8gNGblT5cDE2YFUs1fKmxcRtyIyFAqlQrwyZC+BShrb25/Z25HD6yF001yo/
xz7aoxDxfLXR2dlEI6Z5U/Py/bTPbhm8oxdc+HTCPruwEsH5YSPtjDCEwXtUgWPIFEUudefY1vn/
5iekWxMNyxYIW0zazwnRxHOZEByOQSXz3ooXK8cf5oVkoVKHKPS9oLLDJ2aScUZsUo77ixJ+0XMF
jKcne1j5RQmhM/yMhGYr7OfDmFCFeL1W42CGxd0iffO2eUUdss7LAzHMPBWWA/v1eEQikQXs6ORJ
XIbRCPL4MKoRrVjrrZVULyTaiuDkkx7DyxxkIaafwuKtsJxK7sP/24dG2n5rOiPW7k9vN+zWE/JT
rE6E5QNyXwgdfuzkc4woV4Q7kaEIzStwAgup++1UYee4KcIZmNvSpTntcdiwk7FLbjxK9Rx0UlkG
hFBprEo+Qa8HrFDsf7DHZcEpLkwMsZT/aEGwuPyKEKFfzKX2u7U3h+LZrUEhBvQRutK54JsNETNb
3TUXkRSkXlxY9sE2FRvoGVrcM9U8TLT5swGGfRkfx5ZqPeNq2gBxBVugwb9NU3XesGUmbYRViedV
VhaqX2cf4Z5BZmM2QxTlo+ungEmOArG9DPAHvAgXtEh+RnDz6hKuDPofG2SUHbDuLLPtccjIvU8M
8MbHQVGkjEHf8ZvAbETA1U7/KzE4kYzm1y5ZoSLNk++Kah4xIm0GhYGA04evGi6xc7dMnLjvHVkp
jbi+HpMTHfRuTshcRTgxGPCc6bkxBzUcLoPFRqX2GW6bR2wpYZWAtnxdkDl4WcVd12bng//w1NlJ
OXkKO3zduVNf4gWDBQkggEQE5DM0hLut138XFKVyM2BJ5nIlEvaZSf06t1EVT28kesmJMqJ5rmGX
VLi9U5jUNyImtbZmcwW/7ir4pXJGo/3cU3/L6iwOrrLDloxSPrO+Hvqe7wy2ReMLheIKBwqQ7YVB
fuTyjtnLBoeaqo9vVXDWf7s17A/sCjAxOLVKSLcWJtAuezBk9YXJpQtusxd/XPUrhK9s0o1x0rF0
VwufwynPmnYVvbwK18gm4sUhzzZVSR1LaDCG/FtplahUtmim0ttgtT5+p1LrEaMFZZH0Wj2xtX/b
fWTzOKRaJ8bnXU81r4d6jXXzuBQFsEE/vmDVbuTjVvrrBje0RyqPoED6ZEgPvl182HZpiZU2R/gA
0TbwHlHulWuCUvKIGA2NH5gRSsGP4JbFr0BXeFu5laVUBULvHKuUTYqJpAHUo7MZy4EXk33R+scw
/RzBYpAEcp8Xmtc05ChrYUg8vsBk6mlZvsvT/U65D4RyWkuMEyKLE1iswBGtkWtFFgm+sKWHhyzW
o/tDbBsPF3TT4M1PLBV+hpjB9zx2UGQMSryYisU4+XbhuVdwjPYWBZkj/tDgxl2MsuV7e6IrAQR8
J1bOQ+ZCdZI8wSLmyXmVNiywZ933iQlRTn7LciNBbWcyPuFiB0z/YSbxa/EpwDIIAx7CYPHRQAC3
44eeDPKjVaiBsSLHsXciIFkUxqnrz9YNcdiQ1D5FR9tjhr5NrpaGKzTG7cOQfJ7pbobJuc6HHdac
D75HFk6deX9MzlkDZpWgwsIASL5q7bNOKYRmfS9ZzxRfkI1MWXaZp0ToR3ZnkD4IF6SKePvlTyLg
Ah2YtdGFYJ+zIPnXvoshuLovbRTnysbUcmt3+MtboSFi+GnbIDhTfoTY5xWqwALO6BLHFJ15eTv0
VTu1tET0P1DGZmH78FsbgcwLtsnuQc5WKDyPvoUtvpMs+jnB3GwXpavPdPQwxI8IAHMcuGHOB3kF
fKeIrjWptefulG7Fvk1Y43qVz73iRRmQdsEnpJoeZcCk1jjY95x4WTklUpmIMNSLGpTlSgyCSMrL
hcb8wL4EePQIm7XfH1nBl6hiNaTQ1LN43wEMP98zm2c8qJUOqVoA6mXyuA4ysmaQh/2TJ3aWCqCT
87d3WbCaFBrc9onvp8ZvZSGn0Ra4IOCch7vpKtUaJbPQw5UPRie1BV1MSDy85O7FozeoLjICbXDP
tQxSnwlTvWNcJPaxxrDqyM26k111TO/ZaeEMcAe6hxABw7ZL+q7fwM89jggtFpY6q28oZQjq8YMt
BI3/D1bRs84+snwDbyLxwmJcRL3GuAbQ10XYRb+ic0N8Z9b7gLn1r6dGNXtQc491flnzRvt0xlDd
npMRXAGo8le2Ta73Jyah9ovXTgItOcx7Dig1j4Oca1AW6TRpuHPI5kOaOzXTyVsMOkYx+x/qpTbr
nYEx+GWNu8BOiWs+oQ9tIBBt4hzRjTGvz/OZTzUwLfEguMdxn0eTle2uWRrYWqqRi9KXZ2UF3omZ
2kr4271lJBvnExLXXrsI4Si5LAE9J6NcHbudg1Ng3UKZaoZnYA2mdQAVfIUQ5fbax6I5eJM1o6Js
wPszfYXksCr9Z0qthCNh0N51iGIrK3eRcpfem1K1yO+6iwv+/1d0bhIIregt06Adjd4vvlReHhzK
nfTlCvOfz/HzY8fM1LGbhpULTlM16w6VFTGVb0caBTaN3zaT2Yimdlwi7Z/cnJ5CEisjjzBSHjV+
jIe25tNbYaQXewb2CIdW9CBd4vtjfaftQzU8r4yY2Q4FEbXhfEJWQYyWEThzDB/nqYvG2pzRkARU
AOD/NKuqYJE7uTsTUbc8YRYlpc5o1LcWdsCxaom+LGVxPib0JaEc69ofXgGsnzzTO8ggPT2p4RQp
QK7GhOvzZGQE1Ir/QirGRP/FudWrstbv0KPEGpvHorAUGF70iOA6pUDTbLUDGVCdY/PPH6rL+ISA
8oZdbnbLQXs3Zpk8oHBqLiJdDxS4PHtCWB066G1JTYBAUG7/QMCTaN+JG8LXdkvfW/3pLFl7e8j/
YsAXkomwFyvAuxtnIyFIKodmPE2rUUuV2wg312INcyAr+Ee93NAWVBSHlDZLGzD/pXWoXIS5UF/P
CNI1nKOErYeBkAw//mnjkbn0ZB2TUkjT6x4KPli2wuOIRCpauvK5UDTBr3fUQODtvFJLfBKYSdeD
g6WDohUZJ4bPtWBOwH26RwNQyZz+2xdy5FIx9DM7aRz7UaYy2Xrm6nrRmwoiRppbUE5VGEu+kTog
eps0UGDoBF/hWDKhDhuXuXHt/xwSlKMtIIBt1977jWglllvulJyxRxRIBVjg4iOmvi/gELQ6Taya
woem0LhWZqpcqziG9HvDeY/Ho85JRMdV8ohoWeTja6cl3jYsM0WpzU1FVUDWv9fjEOsQwCF7Zj6x
TLtQDlpMDnzOECxLOWpXqzKHTDk9D0tnnFW3PuxZ0yV34GmKCpFkdE+mEJGXyeDKQADtFVkED5vL
cWxQeWK1c7dvQ5IrfVGwzzHwRaS7XJrvqlkJAHP8iRxD5cvakwoge0m4jvpuamgKF9HuxatgTpBd
u5DO6cOKiFQ0pvuuLqEpzREoR2rU5w1BKIaUAz/yh3zOJZ/ALlWszeKswNupKqNm9KiH365QMH9j
60daygqtggKiBE28yNlZYmX9U8qzdVPwnkqKW130LNRebLvOlA/CTi+5Dp/Oqsv1ackfnpIy09fJ
TyMXwnd/GHX+xtnGIlQAw/HJc3Ysswdgd95qgtBD0HCFoi9JXlUWVOkDgXrA7rFHMZ6OejsAElJd
Y5hdm3P1jANIvGW0St2zayDZgYlWmgaf9PXh6hJJKiEFpJq22N4j6rSkVPM96dL6tYrVHF0wIAZ4
uvKH5+KEz5ooLvs6nz/o+uZxxJOYUr6/4NALeaPqYXN+D8pX5ZhWTCRpvgAAzszR1rs606SLfo3d
pKsHvcLIslZ/8jvs0Kw+dBY/A4YUZqQD/QkfIjClcEQDzujZMEdVS0dLIsLp/nikMZjY6eU6hpAK
5+AtjUF6giXTDcPk9GHtBUE9zCutR+BULWrYMkOLEzuw0HP7zXwExReBznarRSTSEIWqoYaxrqiM
TzpIV3yGl12ohU2OzcyxK3nN1H8JOWUao5Xv5UwJ+F2VeyvPnK/7j1TbQzd+UGwli1qY8wIM74XU
qaI2LJI9y4LZKKKa0dvM6KzFWPRo9jz4LfsdVbzYATb3id+L99bhm0EXPTrvF5FLMWYpWkL8pTl0
E0VHh8SXzNBAXOr0oXzBlxHaW0T0JCbdUJGwYUA3U6VcyXFNngDMMHDq1EvWoXydJm4h3SKJ4Ojo
eiNadRUrRE6dHTpb/jzP2hQnyAJM9PGwwnUUPsJFgkU2D1wzfPGiS29xWSiRf46wgRmH2BY7WDJi
SKCUWTk5zmgSS4BtcH2573/WIdeBZu69+tfDd9q6qh9csoOOxTAizFINKj/cZre42WwvxjGN6ks6
puG21be45Zn1TPSjOTebeSdw4WUWTAvMJoHIx25GnqrXU1iH1ZEBAHK7wQiHY1bO9HcVyWPSU6Cw
5MuEdug7Sis4UPg/JQu28jTlHkrUx71XISzh/rdKWsgDPR0ECNzWBTyYmW2+Q9d6TxNoMLhmxtSC
w640dEz41L4JrHPoaN0QITkzH7Ay/JuJH+jXTQO1OE+HENhMcoLr4oq6ww13mNTpYOB9GUfHSUrk
wmqL5NPISwzv8wuJIsNq1qv9rmqdNEf0Gmx0/1Nt4HveS6VwpZsRNi1iwCs+4X3uPMq7lvf1CTE1
k2p5qvpTMD2bZk/iUdTooBImjzelIl+U4D2HUSV2/arNoGmhzamjtJQJb+mgJ8svlmni+sNJGtra
mDJsLNoMc0NeAIlHJKjr5ns4u2aTOVbvPhmsLMZxGED3JqNg0Y1pYbs8lEFse+L+ppuMwuVIlACd
Kbkz+Eo0ugSmlo8VDjot/im/sOrnF2YMj32X4Uw/nl+MPsvbS7duGEyJ1c+JLxaw5JUJyq+5/hLg
gE3AOjZBjMbBV+H1qr+B40A6UU7t9ZZZZqUvdnY4C7QcO5mNr8VEHWw94ksOT8zPoJtXRpqPzRSv
2A08s+faTnDhdiBYLY2B7dauA8HXGv0FstjE33QuPI5na7nnjQCPcnLo8MB0QHZ/rGQM8/iNHxBq
g4RQo1h1Rf6yy+ZHnsrNEqbbkrgEDbZ9zDbqYw9TeErfbfDFBZm2ePr3fDllRh+9T9/hAxhuwanp
6/EcqMdoh5hiLw90CNaezFFtvPOJJBmKGNLdke/zKaf8RSngH71fFb5b1XgM4Cvsx85kmNIb0lRi
tspTSBg7iXaV0rQeW4ftw8JaASeSD6q3nAgQWRz1mAJWRloiAcT6/fo0nPsf0AGLnWi+Kz5IsxGm
jjSBkXuQKkIueLsMCkPI3AdGKBmIAHGKjfzDcpdUu4c3Q6OBt7K2x7OoQtaJmAhkNu2ICJwyPt/P
AQ7Ak/R7Ounf1L69oTg2nPQNHl7OyNWAn7MHoWx3wZ69WJPgBmI2Rmft13bbVM5iuMyul5fvKSn2
aOBxBlWgkF7kpGIcoQ4zwS6kuAZEMawWNlt4sy5t6fKZhQMlPycX78v658nxaOVF8nrnamxdorUl
EcKgZPT+U2Xt8exbtCyuOMZRi7zKHGdyg4cLyCom1LoBxSlG0179WDUU9OC7HONjG8fOB0SnshWZ
2JCxb02vPa0N6NzoEBoji74jOuTFBUHXfDqCyoR23zc5x2o0cM7+Xm5ZWDyRA3VHxyun/19E8H9m
ZNzfSsibnqcuYxm4UpKSa8Pd8B5krEFwDzZ364L+aegga0xBJ58tydw3YmCcVgsmOux0pVkJDnwj
bAtR2yTdrs06FcR3WKJXzessaCsHLlafnkS5TnxWf3xyaL6IYXJ2i/FR63/pOYc2FcXsbUQqVwoz
yn6QqFRA8MdIfe9jrwtdr8Mo9LJM8F0VhXTDoOB2Fge6RvUMuOOiyLFoPU/wt0VKgB4tO/kqxFXY
UandEDT/PN5bR/geghv5OLm+u7ht8tWf2w8+gXv91r0oSX9rMPQZup7MCqR9HRxlkSuZeQG8tEao
1+XS/9J5ndv7xy6FAsIT2E4swvBGK0p6LwIdP4HgAV0GVYFDiuA8Pcgj/PdWFRQpoeDAm/0vQfJN
ORvX4yurY+/oupRESBaGHL455wgcDQA/4Rzt4tTb9/3v2WhkLU3jbFfJGAsNRBuIYv6nwHU+Vjdr
YdNjaF5TS4gV6C4v7m+FsbKeHDM0b90mF2mOcU+35YQe9175yffaE71qsH2W4mwfvAEkZxyGg3AP
sbJdk/wTMyM+fv0mV9zfn6XStvd2mD69uNqy2/gxMQFR7GwlDctUayPTdurOmDAMJ4+NkyjzBDR3
KqBoTFJO4Eg7KRCgJ/aOxIqune0jO4TBS9fYQ6k3i3A9T49lNikHQw1Dj7Oqx+x5SpFqXxw0BdKb
Z4qAJ9tOpjG+WINejjpWj9Ln3093VdBfDRWzJ67HR5Iyqm098wODvaRvxYaRY+kKt341to/nf+D/
Nz/fSV6OGGR28yP13z0jH9DLjf1HLBmk1NHeItiQKa1cnGQHtjA/IAx5czRoAYGmM+KGSuj1jfM9
JaXqjZ+YjTiRKPcL/WRT1XrnH81QTEQwibUlEpNUpvCqMzFmPxXJQ1C0T9hbfCZgvzrx2u8LVEk+
8Sz3iiABhz/hcrTAbnzKuZa8AkT52wZ1UGSZJv9tY14sZ4vXFJLhgkg5aqdeTQKqTmYnYGe0oLum
iFbHu8yxAACT0iShtbrbcyzYMkGorMdJZmcJLyREWVqKRj/3DxCPUxqM2uJ6B1PKzNvZey34HCNn
B8T+AVp5jhpbJcBKR4WfxxhIDjWgDIG49GWIkSnmn7UHoa0tbOUyGfdn0f2yoMacfKy2W3K+s5Fm
osQzv8HsXI9oXDPh84tXWJ5MS3+rK2WXFPmcxgLJyP7ne9q4rcmddCi0BWbRUdRXvVA8HMRCLnwt
J9IwFsxyd3shnQEkpU7YD3MZEfpCydgdGvqgvkuEXyu0pEK1eltOZ5XFT8lhPTHGzWvtp4S/gHNj
LnUOsHbNi5Kh8fqmN0eunRb9fHtJdVhrCyItoIp9W4Z6epqkSqFWR7dMQqEV5vFkw44599BN5qoa
LU8x5FF5R6xxyaKvVH+uYcNZvM0CTbnbnBeo0OvYV4UjYVCw2gSAsFI3L1BEUmL31wVPAJF9lGzB
6SwpYaM+/16OV55K+fceHN7xfGWHKTuvs3VnC4Ars7E0mrOzBRs0IbA595n8IOGUaPtz/K7RdIDm
pwoEik0fY7EltuWCIkgPZKcH2r4bkW8ExN6rJj0DZdFIOlCddhNnbOThHe49dTT3YIm3AEsUAttl
y4vwCDFWf186evlpAGlWBGHqTXk6Suq/zcR8QQDonFjSOmc9e6ylccAWTIHATAQIxil9k+dso6uu
btTlWOe1OcS1XfMbylunYK/XM09tpghF/6GeTkBOWKsTIvY0u/a+5H+3nxEBj2Q+ZmwN72gvv2bD
4Kvk87jSydssBtZC7Fzwmvh9Nyv5fey1l06jWTA/wvDHa2Bw6Koa3rs6k4DCnHyOSGTQtI3ZMHzx
qNZx1mPXZN5BTI0l7SjUvq4bLZ+soAVyKx6XsmrEHy7iXuWjeUTK0VjEWW+FjukCmr5he0ovuj59
zC+Twu9dYzBG+ZVt09CbDVgQ0euM2Ejl23sXjnBOURmaNDUOO6sTPT8QKbxdrLsjVr/YXXnxRn/0
jqf140/6n19rCofTrlswrY7JoGlf3Jdfw7Pr752RySLsuLRKb1hEvP3DuIaoo4LgZBBQL4Dityi+
de7yVgtxM13FzefaG/n+nF/uDWCjy3ld5yIXjUupCpeppm8Ppm3wvDeQJN26Z3Zr/zRZ0AxQa5ri
fuKT9jJA/b5ZUiBZd/3Cr+6xdMF1YnXUY1YSVP9dDO1HqI9DtiBQkO2YaTMXFx2ClPxij3ZDINSP
GS1N61m/4v/0s6MMAsNa/+dLJd3p9vXWv42GQjnQIs9w3SMTxBxw92XRkzali0E2SJRQLJo0//7/
QxwwYuHVYcAUhavu2niyMrmY+HiYNNaXvkGMrYAAiN5NFhROILgVbm6ADgWfwbDgEcfQGGHlX7IH
YnsJOLgFW0Z4G+VDpQGAIGU6OGQUi1Qji9oWogYXpcjhP7xniFDlD3m2LPCoKLwMrO5zaU+J26gs
HkytGZ+AqX9uV4V1KjboIasL5Ycoer0z0ScY1LCoGvQe8sYpSsXy5Ez0rY9/s0KA9zeMpzyhbgBv
eCeDpiLsDCyxCA3O2C0LahDdBQSVTrD5Qm1YrHr10ueSUHT5zrH3TICiIbA9YLoGb6MOuEAE1U5V
zH9535mdpz+zxARiDrdRf5dwbzmoKcBoqirKMZT/rkqDfrcozH9cpi+pFA5csuIkdi8l7HMC/+4h
FRqccQsw+4kD7aA+qjy0pkEW0e2iFxGdWBn0A41fd3aJlrnkcceNjkXAAkWrVIIUSf/4y6yl2SOO
sbKVcO6iii/c2tEQVPSgZFQ0mgD0WOn3qY8LTNcTq50q/a9U3apWFuDtdDVlbdUSP7EvYDjdYfgy
CSxm8rkt+EXnurYdL0c12cGL1p/UlCFc+5Y8s0euuvkRNZqLfdJKuUNO0AQQfcZIjarE2/vXj6V1
EOZsW0G8JUIqDljI5T7bVCkySqtkSHYCZmLcbghbQ3s5RRcAlUW+OsHR2jB8aod0gwEalRfDWSme
joWwbULtE6Qkqvyb1D1v4vOR6HLT7lbmkcyoYo0bTF4q13R2XqozXIPnuQ+um0keS7q81Nv0TtY4
DhWCgwKD5xRKBucmB+CFb65mi1TR7zqmy8Mnh+ZUToKoqW7+jJisAenb7P5HjnOSB2jDxilphvMX
x8d9Hc5ngYYRLLjH6CNX7SYJWuvR3SH6aAnxedr7aMVgDNZcUAVOMz3ytsYZiofsQJTYNDImnNno
Dw+ZqMze5UUuYl/PhbSb4hjF5kG0Hbk0dMZPdrACfbxrTbgd3l0/HWmLR2VhMsIZfsAnbJtlZJxH
S8nRMJfJxroU3PP6zLoUScgAtpcxh4kNSkpwuTH6uu3edqys7ofoi42UXoFqFoxDmc8LLEzprHwZ
Ehi6RCmnZ0h9lKBTUV20B5dwK1Ow/b89jzACH6A6B3dgkzwC0yi0qMBL0zwJEXp8L0BFx69aLK4c
FREOwIlQDyGRLpieAQ2D7VjyXeTsKF4+3fhGFaM7D9gO9ba0RnmkIW2PYChX14+G1hIildu38O3O
IQWE4lSQT2UQc08jJHhvirmeGfcsNEkfbtUxciI75DpuGcMM4xUvRs3SYp4l49msZOVEQLp+ILZW
ybjZ9+fEiTYdWnTHJl6X1vYvNdej9M1OmZN90xdgdCLVv51jYNqlpc8SSh7sWwgcOGGTW7+3+l67
y8qz9Ah9wlWHvi3wMol6lKV4Bc6q/n425PEgtp8sDyD7mIUD0mUUaEJHQywfUpI4Tov0xazG4Cqv
48D/QHIkMIpyeMG1e1HRQ4TCL/Cf3WbXO4UJZ9O6wcm6N6PnK2i8gr5aqYp4v5T+0SaDu73Tf5+8
V+S+q0JuV9gK5n3cdROeLTzI0AuXKEcBs/Vzv/+AmzDklTegXUOLdf98nJ7VX4SbrCwARNCyzRbY
vzHG4PDOe+MFp2FlPX59k1lxb8xX0vLTk+sJRe1CsBmYDmEG0tChzLlu9M/wlGtEP2xE2ioLSqC1
6n9VS4MsKi2UmZg3WMAuz3jRNQO0AdOHFteZmMJpVJjjZZthNF/9N4xPSbxqVbV49B6QaT5k8TFF
3FCfXVsfyv2CwpFC0v6VwmubopoVZI8CwYsOrB4wyKJIfGVcRXwbmhZ+yCLMxFpVsyuZwUXvOlZD
6UChGiYyVSmk25cbZ599Rv1oKo+e88tlTrTUyGN5XyIJM6an8/NhpgUizawcXteuQzb7x8FgTnDZ
TMpN+ualR8Hbt/a+GREsyqBvtIIF7lNiS0WYhyH3xGtdU9cy2NsL/kU9dRoSwgyUj00Dyc1VW9zD
XRxfabimtr69chhZPd6DZSnlRDWh6jd1WCiIap5nvblJ9hXU7FvCZgGH0CK81Ygc9jOXtU2URtwY
79kxgPTSEGw4Iw28Wy2aRUi24SyBGGYG/NosvBxM7rCo4HlSlLVki+xO/UMocytGXAhBG68JLVqR
bWN3nA2r7GRcy7DKAqNsF6tj/kBUwaFJumHPC6RPKOZ1yYcVbq+Z0o4tcHq54U6uZwm0w5vOeZ8l
65iih44ygPfMCUOYZypOOBy/QX0ioKHqWWsvj1GjiIloCLYfvWk7tcso3KzQhghyivV3ZR62tbIO
aduEAFGQ3upmbCqPcjKBGuKGW93g/0AVmlz77x07FYAEJSBmPZq6k7bHDB883tBbJH8OgOPE0sQ+
sZ5QR6dqUHwwWO24msZmt7TEnLvGwYy/kL+C+eSFha7hb4PKHyYNfCMgTG9YFynp94irlvg+axUP
dC9Thw+RqCAyfpgSx98gbXKxLHT+RMFb4M6kov4RH2eKsI9hat7sdv7BUtTfXRDe4Be+gopA4FPy
+77y8a0xMac/D3qSwoaWjWipNwLTS1NWhZMmGgYTpnF+ankmbCeYCBa/rhZLz6ap+bonrEjOzq1x
HGmGa029iCvCid/SRIyiCM60tgRYLpMhwMrNjE8SWMr2Cs+x1lZMyQehf26mVZhAdWq3uBhUuDdN
EZ319oHx/zICRaobkgHftFhUsq4Y8cchOKoZfaKy4v9Zjp43T0vYYR8x7DBj45PDCo8VuRCQ4Jz4
SczCTwLS6AjiJ1khNXtV7AW2cfjCs19GKIQwauQuc0cLoNmIV/IjR0UVhVSeixkYYKbnVxPzaltQ
8odgrWfl1AuUTy0SKEbNOVIjbBQNTKLEP/d2vLpSAkZ2vTs4LAZ9KWYP4l9g5ZgTDnIhvfRxSxGI
fBzwMKR0TG4mso6aW/WKlhOuzZlc0/MH0WnPr3VbS3ep+EgbAr2W3Yx/OI9WDwC7iUYD/0/Ei4zy
MNWUojBV9p05gYYXC8bRpp0EgpPxsWl0dJ0846M5WwI8JoQGC+/uPOODS4X27hXgnt5HhY3qvtmz
n3DJSk0/u/w/xEEslvZUun4NaSsmwriKuAd9G735V33uxZTStz9KH201fZRKgyKIYXK2Kt6kWBrh
Xg9dgrbYeBiUD7TUhl4qdTfYrilfZ8EmlEbl5m+lMqXR9CcWHFVejgfIXRsF9gJsEn7TYoJfvA8U
LnVmvPh9Rr2yN5EMAOTx4mpulwmgnZ3ot0l5WF5VhQ64WZML/SgcTjJvwM43GxD2v+d8pxfjuXov
pIOUFMc2HlFV3w0yvvI3JwkOWRxdMiAaMWDeTu1FBTYREktfkmrg1ipit8JCC0oSH14qHHgqoEjC
ouvMbr6XyqVTRFTbcY3/Y7jOS0Jic+kfcyGkhmQdcouEkXKyeRya9jqHe2VZYO1d41szf42aCgCJ
dzh+hFNAt4e6Nx77fLr2MN0VT1Nu6P3AbteesglS4928jMY34du7oZz9kWFu16cXIU9ySqK0sOHJ
4PerT0g3wja074OhUEYpH5ybI+QLxya0YnOneoiV9tfY3LMzKPh3pf7LMC7gNt9ip7dMXtkOWV0f
xKcNWltZtecOrWF7IISbnnKN9H+AmQ+V22mDH5PcmQQQPQLIIpocVjfrA+1zPp2WBRzf3ZDBgzUB
1o+apCbqPKkqsXeEqQYLJ7bFG+9De/vNNkwOZPIQsuMkX5JWuPpibMyeXk6tGFAcmxkQRgxxW1TS
81qr7gUnRr6cHzu6O6DLt0ciAZFClSjc47gUieJ1Tdjsc2NCmo7wqKjb3bsDIWucQlrWA5FlL8Xu
rffU26iA0mmeosHocDMZylaoaI/CJ1Lo2Ua6pLnJu7uNJMH9mjvn84pg92HQha93crsLmdnnyZmx
fH7c/ee/tccMMv24CyLd6am9skWYNcyWEuzQHxI59JCdUsfabqMrdUQESZAFSMGmGOp/bojgQyo+
o+tCuI1S+F09rqV9ousCcT4tfTNXwBKRjrqOHj1I/HeMe7xe4EQNeh9erskuSVYhDmrgULxQELxk
CfKLui3rEQAQlB9LYVoI/MhEVNQ2Jt8qSuxjN1cZDocjUefyGNK5rzQN0Vb2UugvBa2UXR/UFKXB
MKyFS1j5PMIrbj8cVnMnNSff7zh37QkKDZRdIsB4EwJSsWcfjZHYV9SDd3twmQTgSaxdfutT2c9B
GeKbOxrifbz3Zov8A9hYpNAh6GQ2UHKtvWOHONyf45EPzl5jj1pNTC/FTXtm9IOeeE1m05fvlw/w
fi8uBEHkRIgg8r3bwNhEyEsj4HAiFwE3DsTWIwt7/rg+lTgqoLQHGwCvBuy8W0AIRVNvhgiXTtcL
0IXswUrYXssO8DLQg0w9qFY3YUgExiAy/U0Uo8sOOVBkUHbmB9DE7pfY0lJP+ulIbvZsDEFlAaLT
smS/+cP8rNAdkHUoWqxhVFYzMpz23Jp/fLbZgnAcZz2T9Y1kAmulFRr0XvFF04alNsNLfxg5g/+I
mNmKOlEhTAM0gbUQbwS2aiWce6cVrHxBiZIrWsBbhCrkT8TR7IfQ62qFPzLTbWLCmdX4Bow238a0
Pck1kkhXn6lQJnS9kmNntoHsqtq5L5eKorDFOmJkxy8QpONUQdxOZRC34NQymE8+IFUuFgAkvPiM
JiVSClNY1lNcIGJxnYrm9Mf5zUnby0v8CDvvWGi3ux/bazubD4Bhe3O7f4Z4jeTDGB6CU+d5S4Na
PUHvbf6RLS0Yv29+f2PZJ9ywZA3v9KClNF/BAH32mkWByD/kIYwEwkgsOQCOgnGDiVMAnL4aK3Tx
ibVYkn9kcOHAeT20SeHvb1f7OFslTDlloErEB2313atlKREkMasSxoBhYWyhlAWUlCP5lfaOmA2Q
ztb3vbK67N5qv9CbIQ7Zn1N+qHSsfvyUUY9GakGHRrQFtMJG7xEG/bxx5polj+RYdRs/ThZ4OBHU
Dti5WRRYRQcnTMGmCvgV44zueCUoCRuHldHnc/8gFzqmYaqNYj4450iprSNYrF5J+WbFplIwb61y
sj1sSaKFGjRfNGUcKZOAp5gG4gqV2Dj5DuU2NnwcoeWQwqMQFaWiY3+fp/twH6QQxzNXaVCxz1Kl
TV5lmfve88uZglFx5YXx/wDJm+CK4sqmgT8/tTp6aK9NWhq0W2tK004/7arf2+VTG+bNARUoSwn4
HdZ+noPu4e05C+vWONzuCmr+2flEUFCZz2tRFKD3iJjwYgLsSOkvXI5D/2Y/VwMxng1C7CBBAJte
NXK39caGdQd8GVYb3hRvG0HWQn5fSPoCLMZx6VUMAiWPSI/cIiGJ7UXu4lQoFtgXsJdnGByEepGA
xs4u+k7OIUaveGXd0RS7jC9W4ZV2yHaaYJ6CVB6wLYaUUiuR67H/PRsv7xm46TSX+WuHovsaOiv5
x17Oa43NKZrbAKZWmv7a6YF9nol31GkJ/5RLyOAA8YN74oKtFb0k9nz12Jrd389sjOur2URrYMdy
aUjv/houwNXTTeCSUo5y9Ogk4iTTH4f4LhNNrntHqS7fxj+hptFmo3Q2uB0Ks9E0iJNiAtWaoc/4
+dKGnGgOUnRpmukea04QnGfq7aCfes/e8Ek0g2XfOXF4clg+cMxznzuxpPen46+79hV/koMTrRrn
IIfyWHudpuguCk5FiIWQGbJhVSZ3+Qp7G9XlTGfqMgTlCoVHC2kpleYqsLuQt/6I5R/jD8Ovjvz6
IZ/oclAsXeZQPu5XHaeTpTqirfRoMIX/qX5VxtzML/dIyDYXBkCi2Z5DfYeC8X5RE+frF6/gF4Ww
C7fqz2DfrrDJ4qKbl3+xbgkTOshwQgWDXvhHOzDZQdOokhl3l5O9WTJdzzox8/0lYPc8B7VMg4lY
B+y1P+n7IA41DU1GiO4lkeRSHcmCVnlb/bmaYTodEXz88uUQDQSuev30awpUdSNv7dcKLl1ZcEku
ReFJB/5pN+86p+1Q4CipcbpC3nu9EZSTDVHC68hpzO7YkIaKtxyHdqojWbuDFf+TJhnC2gfgg3wa
Ux8Io8UJNbBL6bo0hOHgaFhiS9kUf/fuYYc6HrRuIJpQxCh12DZ+6EczSVdJhxUr+wfXJLFzW0Uq
3TQ5mdlWeMCAG2NpBh9WCpd9iWr3v2I2/DxCknQItVt+W2mN5BixKcVmyPYEytgINPTznCrNFrmC
hjboi0DhZ3JeEK41afRsbC+iJi4/y8ujxbJLSf2270ufVdi6foq0SpHd05RTkIOjpa1wrA3Eoa/o
pw1OXEQFIj4hpCsGLho3Le+5R1gSveMmOLovUY7omkSfL0BohyCqDRUXxnuJ/NUsFMDbcPd+XAuH
i+GSp7OOT+bfVKQ9lxlmL71XL9lXSReVeCrskrVgoS1P3lOTCX2G6W3sFZMw4t2EenDrsaIT1I1k
absJ6+p4p2K1gru/h2snZL3hWZsLYZOAODEP8rg6Be+4EQqtuxTvNcCH9W8M8ToxW7U7ftEkw2Ai
BYadXuFuJDbkuA81lW9nc4r1rBExR0ih0e00ZnCRcZWwGe/q0sTN2TACqiUb5jPVzvcomZSIoAry
lLcASAjXPLrqTU5m8FYW1KPNFoFWY1QikakKhuki1DYZPNYCOsrp8Tn8EF1ZTm9WRq52L4GnNM01
ZWbk1MQLrW/k+Ii8X1VkLhRiA2mQzYpVMzsQV0T1DWKwDQV4j/pCvuwGk7bfKhg0sKP1iLXfXyI4
Lnv1Qoylk7fdrx8Vp4kj9YCkF85Rq9egizQUoE+kllX2YwfjK+D9mW0xdaFCfCzvYKbjgDZjSnXv
XmD6RpiP91Ljh0FfV4rf9m2B6qJtQeZIblLhINvWwBUliGRl2Sgy/H/wmeOVtPyTSvRKw0o19427
x5+/Hkg5sxTjjXi03MyvbNe6QFCjf4YKp6XRmGeJ8jIJ+UwuNS+v6f0nGj5EbhtJbXFFl9G/H2K3
8SBBeHM5B7HeElvx4dwvF3Km/KIBJ/ZTLPqSqaVUFoPSCmUuo5dUlDAj475Z3NJaMLq07z3BeHQL
QGnfwydDsowCBDqT5QCutSx13q+ouCngYD1jdh9n7vL4ls0sYZ6BN+lX7K0sRknZ2prOnicEVxvE
2tTdXov6B8qa5WFX2+jHhVZVvHcl950vfflbK3oIDkxJCHkEX4mVu7kNXHtwGQ1UWk2+qdo/VWxS
9mBorkTaP5tW/28IBMCXWnNeGvf9Lu3niKyk6bdMFb9drUReq13C6kLdJ5ETHPkGpzpp5PvXuR56
xPY/D+6DX0DM6rF3xGLo6Te96tg4wv6Nimx2AvOyVe7FkmadcRClgzhIbsBFb6B7yBCFmnoGAY8o
xsedr/TUIUVgGmEy+QkhX2XPUrF5Vgl+sJByrMKbYYJC9KdHEm4WQjI3o+BJgONhZwpvrusAzGes
6HNx+q//MyDaHcIx5zqIC4eZjTzWmhQPELy8G0A51FVV8rP6P5Ao5JoWKV/zOHnum71tmJ0YuQLZ
RKPpU9BY34RlQdeN/Gs0+s4QkdyJTDg+WcUMw0dhxMVKqdunUcHyLW7off/VQMdTDUZ4OI8got6v
DBWH5uhnDqH51lvug3As0ZVU+bRskf7fLSrIJQjdsHChcQ2KulpmyIWx8slopJhO/zWgnes3dpdM
O+hCr/DOthYwhXfMc7kkQ9CnOgnUMlY38YV2VBwE47rMU+yUMXL2y6z8cCmv7auQ4WSr21lvYJeL
+UxjYqqOzAbEMQRDw71kolaGxPlTMH0+nnooA/8yHYnjsAQSyMwvMrVnuAuJTAIMAHpZtRckUlmd
xeDSMVHQqFKqajijRarIKh71yXO0pPeoRaUcqTUHEGo2ZmS793IPTdzXCZ81vjZELC6DFMorT7OW
TxRYtpFK2LqVeGOYZ/OF2doZ3krQXby+EC8XWDdFVmOB+tB/W2g7kpGGzL/xFi16CEfpnLCSq2l6
xTnvmmiyg4C3nQNaAEEB05HyIc4WTJ4xO1pUtuUJTxlr+UeWV7JKX/LJIOYA3wYXk/e3vZw8Zwnb
GAvOgsdOqn7g02t+C1Af5PfCHR2Pz7Vq7zynMiO7WV5+ex0Pfu7nbkhpg7z2XeAnbVYPVRfoJHKJ
hR9NJLQgSx6Qm2aubRDSgVQx3BTiL2UTGy6kLY1QMzcjjd9FzIFL2cGnqfC33oxzJqSbpD3ZIGQM
R8n38gv+Q9N/o/2yWwy4lB28SF5KMZ0AvFoa4+B1ZPFYpqdzk5774Za4ToueuiYcqMe0FvXg0MgX
Ahmgf+UJs4HrCkANx/JuHtrBtjWkguI0wpYI+Jm9B894Yrs0ERDrPmFVA61L2s/SNNGaIgXMtiZm
Ac4XS0gKftgAVEB4Pmt/Lyl434ZR0ZidqPz3N2BcLLXE2cKgMTdeFLJEEmbThEoVG6BfjqshsQAf
bdDdNpBYKiIYLTqaviwR/hOIB/e4BQsZyW44Ox18m3JZErCQl+/Gi++hZmIg9eKS5cHDMiY+8jeV
2Y3j5MVWbFXnmg9NENXbPEKiGF3Fo8XC8t0mNv8YOJTKq2I7lHEMoYaOTsc+PeE2qt7L5c0wVOeP
g/b5QL7jsXlvektkuQ6Uxnd2WsfiwwiK3LHoE7OkiAsV3t+NRAd7FPGbOjJT0SmrIYxtBXc3KPEm
30Nmow9JLcnmslZTaiK7OuDV1GHVy0E6209NTSCcG4P6qzEnrGDKTBOR9RlNzSwf45qjOy9Ni5JQ
75EfAQXjYxxki5R9+h8o4V5uDiWKoc61Mz2qBU9izoRPEnon1cT6r0PQ3reSckx4qsPzmddAHBu/
UgRuKchFL+8kvyzYC4z/DUJDUyrxRR4BWjM9A/p51NarPRwuoOjjDeb+ZfQJmChmHbQ659miYvRX
XscQ40IdarOQw8ycVLPjq84OItrjrYKYJse2JyT7/Ve+Emmp09996OnzwKR+AcDpdtjASDLMloQW
JZQZv6EwwqTCJa8ZoUXZQAOM3iRLk6eB66VfGG2Pi5ZmatR5qTVAtoepi+dtJ0xuwFwgIEvi5Dr6
lBtCX/B8PZyMfyuqRTQXykgkQy0FK6mSsiCRhRdB5oslt05Qgxb8CYRNE/YkqPdh0ldb/qLDcysE
YdLvdsJ0QYCYLqqx0TePGCPZsjpEEWXO379oV9by3v1YL3x/PRE6wWW5h+NbFiNnNnbl4Qbkh7Dt
Uqm6MgIWTPEBfr+VNVqC4ZWRzl9B6ZrcjzZ3lS5ZfZMLkLRWa1tw21zVQBz681pS3vPy5ByWoXMt
Mteb8vQj3rLWBGuVqVMcCWz6XRz6DdQ/hD3pKVMB8xkD9VUkFJNSlpRradlkfBH6MhCilu9vBXjF
A8InFQxQqUfRV86mGLAaObBpGqibFVoYh4SFg88GQncNunDb2AeyOEkwQ2JdQTSa/e8U8WFlUMEc
MLCh/3I9A+tX8VM6KmmwOw2vnYPI4dL3hxoc5dwn+1B/L6edlSJKHfBovaIeNQZ8nsLNHdyh81Pn
k+Llzy/9ijqkN9GjK0X0D1telPhEEukpi9JcKDtvE5d1fyDuTfYQgAU3dnx7K5lZernA890m/4zQ
ADuYfGfwCF9s1bYOzqOUZvLdoSfeDsR/IWfM4e2ThFe+A0a5NKMniFnVRMHnPioIExfqHtiucMb7
km0gT6XQoDtkOF31CNXSwGRIVFzaIHbNmAq0S52f4xwDLRD0H1c/PS5SRaA1HKrdvm9gV0vKTn4W
SLOEt6t76UIn1FzXlXGC0ofKuAI+XFLeZUI/z/uvsnnmF+N8rADgjXQzrIgdjiCrua7IH5fovw9h
sBhYFtYIOIvF1vBHqCaVs7dn27EuLIBqh2UiXzmabRi00v/8notfju/KRQ1jpzwgtX1rjsx7SYnt
h8berZupKZoCnqKi3tgNS1a41WD+nV2R3GjRgV//mw5Jz5MW6b9FGoL17mgu0iiTNBb9VSs+Uuha
6fuYDthu8TF32VaWb7Ew2/7KeS0vkoRFcAJTSRLHHEOAysLuVxeZc6zZ8ZElxGbX+CgSP1lgHI7/
tw/NOO6u7jb2R2vYVwPNIs5sjPCJgjloOHmHAJAKQlZis0fdhuUsuQ1dyzQUHr+Qx1jX5hop9Zwq
pTZIzZN9R7sf7Y3jym08olli7JayozamsGtpEw3tn+NGgPH3D9ckgKaB1HFQ0sdMP4ey9BFJHotC
YacXmTAE3fhKhEpc3R1LHu+eFV7PiFSvT0ZzLtN1AatLYpGi7eF86YV74mBLQwnbbntjrn04bEH0
RieDqdLUlnyBJLpzoIy90jBQ5l+moLC+9FNawCUip8Nf+CWBXCod2ur5ZQuj81CA3e07uwsEih4Y
EsqPgW5dME+e6hQ+t5QvNBLQVYkhKC1AHKJsBvfmQ+xixQa4ltzNSC3l6pRKYinXqAzvsBUkCJoj
ggWX6m3AcfVBCD3bfaj+LkQDijj7UL7eL6N9+dbGCus7xf4MYtQGndEgR5KG4XiVvCgOA9W2ndrs
xxRd2RNpd584o3gPX5dM2qORdeML/R82QaBV09fMeD5KpykAQJhl7Ufb4RIdtXLnyrrKILwb3t+v
8nS531NZpqpcfmHZrWAWkY7U+a5h+l6SESA+ZHIssMF5xHYDstaNTX80FxxlbammYZUT2KX+OuZF
bj0GiGWzFGCEd+YfKM9yx6nqmj3eOuIlvMsHjnVb6ppvsTu7dAD6UxJKEeYFYi0aCZpp8lkPhaC0
5UZaZaIf2p1iPGCy3eUqNxSFD4OR4IEfaBOTJ7PYARvYjK155Z1kDtz6dzP/Yfvv8R0/ZYb5w50Y
Q8Q/hJ41gEVsErtzhVbyb5SEnTFV0xJMA9mK4mlgaq+a/3DJFVc6A7UA+iiwSU/l7uy9V6oMmdaw
WQNAGF84X++PjLn91WcSpRIBdQPgd2wyzTo9N7eCs945UFMKKxjd9job9it6gYa25pF4bvAWDsEu
3O/b+sPAnzS5iaPaJLdtdOU8ifeJ8mqJ4KXoFkIqcbgb64+f6R2Fd6/4yIqZ1B7xyCAKF9eZGf3a
IkMzjurpxJZ+m808zd2kAouYBpAo/ALoYDDwq77qO+jIyDZK5Aqi13/Uu9EzGwsejpoTchXKqkwp
8qHIgD2tAGDFWIgVTlNeJIUD4R55AZt7e2iOD56nY3tHCs1pYFmkvwaZJ/98Fv/D3v0SfGJucekd
+1uYCkxHDpvzYzN/N2HFFtR4vb+35P19NfZvz/RKlGKtbgZii8iAbJABuXSXb41L7pKoqVS2DLq0
7/C3qJtpO1g5cMDfaNnQLJkwq429Xi5AWQZ3PI8KhulkgvPgK3zT7bRBFkjn9NvhlltNEETRZoOT
3PLhbXLcvHFSE9iwXd3ZZEMqCN285AgC0M/7ps/cat0RJrmulTeNsFVPvxP4cS6pP7b5fM1k/i6S
zThAuL3Xtt+FV7QUR+W9tZYZVAJ7kp8wP57Mh2qVUrbBQ3BsXVb7frF7BzuMWAe1LcXf51hBA3+N
FmxVSsKJxxaA3ldrcEoShWLDrbv3sYkHTTspqL6OBzIgpXTk9SC3ypFe4ZZHLagAussoH6UVc+JU
eNZW7CerjTuuijg5+26V9IX8ee8o2ejFcJatbUdfh13K4070iCthKn2w/5A7ezPiO1MS06vNC7dP
lgJpmsY8DWM+rsP8kiDAiYmt7dMRiErFhRX4ZH8d17XnYYAOi6RwVgSYq5eBTzGcmR1cDM7Gdsmf
bKMPVQ65z6SDhz1zsnY3L7uH2ZL+LrxGV+tYjYdwHdT6CokewsTEK9dTzk/l5RDevZ6QCbmJqhJ3
p/l2FDBp9hT4P1h9sdArWx2H/BSpfv9nqsewMsRpOSY/15u67s78eZ+lYrA7vTmw3cO6ZpdFfPBc
m2Fw/pagOzKh/NO6bUm8fkRC4ym+ITBZwoNVzKVgfKAX1QRNOsSpn76nTFgKMWw12vjMm3T1z6jN
HTzH41hQSW+ia/EnbB3n51KRiPbMNG6T+lpBrwlBFOr+DNuZn4ZCyalvFEg6w4h4kL0CZZRZLsrD
w1ggp/sNx5aoax2RTh8p/i3v9sdv08iELTdpwNB74OAsl7sJ9yz1HF9jxHZRCmAQ00MLSU2DuHhh
ZWODMiWr2fIgc3HAdOoGW5hACjcVgIzoqDpKiFqTwrGXpwiQMMx/j6j7Kx92Z/Cg2A07RVK2PJ8Y
dT5dVBVnD+pzIhj8dQeqrEfwVcLlEo8lXH2guPXwljivuPXXtzzlEEQBxhrBWxbo/4jXmX6NZjL/
X2aTADymZIBPphSdXzKx2N2xJI20NRu6lown01w6QiIwYBld4loITwet4uer72Z/KkZ7bMtXkDIi
Y57X4zfi7xkUxT87msm5VM6Ckrdq5XuTDMkBFa4DchmC2YWzvgIAk+aM0R65Bl9u10McP7tmKe8T
DY5ZPmP01DMm16HrXWCuUTrsyqwVZExBNv8gr1oCM4O8IqAy4eeyFN2qGHb7Q9j8TUzCaQf3Snm9
fK9KdSge8//Se7FkrT2fd29RlMgyx8xHR6weLwOC9VlRxsc9aGw7DmJ7DPE+LkxO14TSzl+cwBvX
QwGZctqTQ+by6a4PDc0dfOPMQWLpTO0+imxmCvuaBuU4AkZ2J41/CMhA2Y+I5DZFMH1n2txYWn1l
XeJRDt05S4C2wpQZd4m6wAvMid2cHkosL0DWozDKJGE0rXL/1h8JogimIxZEAyk1BcB9Gm2ygFpB
wgCmBY4qOQoVJYX31dZWWQUPmVRkqPcpehZtChqHbkGiDKaohG67d4oxNn6yK6vOX3yc2bQo3OB9
QqvNJXYR2jwG8d/Gy+P1JGGqcdcwwpi0D3lIdyOANMcEpfWqMKPRl+Jsh153fL0wfIJLQPGdYrRM
Tbx7zbD0WdwflnDyU1r74doh19HIfX4KSUaaGvAZ91iq+y2OweISt1ihjHs5f0UCGPXBZeB/nFNX
fKf4nlvutYVFDt8ap8cAEulkvMQeg7P59nTlMqjUpwmP5GG+61k1s8ihsWn38xIsDCcbUVnTmP03
fi44ryPfT9cEEjEOUTFa6CQ5LB5qI3/sn8mgpiti4S5Hbu84Rfx94uJNdJ/TLG3yI+e/sfpJFw3f
EHg81iCQinZMMVFpBG9152VtwDgUWtNvpNBTiPRTJ469TqqipHZ8ufengN+R/SwOqoyAtHLfUcSu
nysR7RAUv1pEkNOxwhSdAavRtBwevBlCrcdjGRnuJ2b+Co+sS+hAIlsnrFaxGT/+1YZE9gu8nW1F
hJe4Um87GlrvV38+vnjVG//rPBAbxmo+HVPPjS5zWoxWW5361MA1EJBLvkDUoYKMGpKbvjv5uwWt
QV4+q6UXXUG034ulKsqQBT5y7wF4QRP0oE8M/MgMUGtufh8lLfni5kwXWQlVXCmPz1IAjeVuF73J
2mJ8T85Nr7e2VG8ZGZYVJ6vzm1aWgKGdYtW52bslfUbEHb3TLzhiDbP5sjKDvEhq7U6iIb6avMsq
EfoRDpMVz7Geu33Hl3Xz21dJeQS3UK8cUCzl430GgCgvCqgSkVjhoYLyi8wPWzcoI8os1rVBoHXm
5VdvhoARmmnB67b3I5K8lAducP1tnK8XJwJRMbjmOBe+YSsYVd3deuYRrq0Uyhgomcx0W4mEyJ49
91WJpiplcPIIbz6e6JAJPsNo3O/iuPK0GmzICNWH31PhBYrWKEhWjw7wwHVW1VrXmPs9ESzhpo1Y
mqV7ca3Y7qjTFDW5EL5+0OkNohh/CUGLWlfiyj6SkwoG3wfMEH2dQcYZUCxzA+85VJdnPbwH20jk
Tp1UofLoFFa6lGAz64BVHGmoqSMwB/0RyLTM8nyqwfFZ9zHgiHZAXibq6rkQxVA5WmPcGMcTOPS8
3ONV7qWWy0EJJhgCd1+9h6Bk8TEAd/ptv2Um0OdXXzjzEQY1xV/EhPxh/IdBMuyjQM1YbMZ70IGL
8lTk/99talspwnmbHpOu7BQrPFEl9EuL5JshBIRDldMSB5kC9QVGQ6YSpsjoEuXsh5zowUKVeRD2
/lQv5QAYh/dNdRKeVG8cW0Wip3zoC/SUtqpJNeyflNfcvmrfA8nRC/KIDvwIJDU9JnQbQZCPoK8P
Lxoehj438rynoITsm/CN2tpq1trHNPpwrB99b+AcKwJrWe6V67wQXo1xlfCIv5kxOUT6XKgMntqF
vXt1dqLSk/8/bGB51VSc0mIaWRwCwIsgLWrUEjvAxgDvX6YJxhuIjMIKs+uuCN/wVl8adp3Iv7Fp
Kjgp1/ziL7dp39nC3RI53ksZAeuxJBBhcFBYL7cLZF6uDT3rnr1p4AX6BAZJto4e4orRIlyFLwt2
xU3+EbFUJRfZqnTKVqSNDFJQkujhtatrHjmywLicosQnRkKS5QdAa7lN0XUozhHiphbanuk+4/Mr
o/PgYu/+tycxdOjGhlLUZJYV9EEvZ3NQVaCW8HDx2E17QrIl6KoRx1encfxjFhEGPZnlpCTpqv8X
G6jmMO0JyJiyOnVgGa0vIgPBkCq8eX56n4QMXKDPxeAG0q7K2VOlXJnMO2ZW86CNZNW9LzGu1JM9
WWNSNp4uOLTXqIcWKU9OesQP9PMwFgNkV3AHiccnZX7c+1ntSUQy6RauFjJ3pkaUkDDanfY2tbVa
4b7RcQ/Q5Zmi2lI5AvtM9t+YncNXlzEKzUp0oh9z/qVlbfuwp2eDqYbQ5JLN+Pr3uOTZMGKWDGlT
9/W7S7QdVgHYGzawRK24ZkfBnB0Wu+F/4cOeSxL2Qmn+WEu5tPmDXcz6ksKHzTKbLfAyujl+7b1I
knKFW+1vNvUNWjyYWvZcl8V6hyNdGGixY99uOUDHxrlWfozasxtU/ZgOcx5iSKcjw0s4rCoyDcUR
sXkKdZvwjWZnr5wuIf3tVLL2g1lrJ5KfEUGQAdxgnwhPzNpSJB2Too5ndbzRwgVCgQXRrT5Fqan9
SVTVQ6Taz1sclqLkbivupEyqhMGNmG3UHJ+r45GpMsVl4nutWotlYoWgq2+Nle8pQOAo+XzSB1CW
frVKo7d4SdLjVR2CWlvGYI7/yYztQfp9mFR7Rke36ctYerOZQS1mhwUOk1vOHmWTvAbM8Jm6DSty
ssW80HEeM3zX/oa8+EZd4BvanDNgq657bDTQSd4sMSUr1eXpNJ2+NO9hPUr3wtaaKf3IDqKnkYLL
SRk/JvqhBNK+LpZV3GohvARGik4UdqC+AXUJ2xTy20wiOyT36S74YDQ9XrndVRokZjUJbLGNC4sz
2OYDbg9hy0eiM9Q7eWYvmnJ+y4D7BG6oJBxsaH09M89SWmnbaJ+Owgtj8SNz2Y/oLyzQ/QqeNaHM
D4EYoklXio/b1yUIV8uYWPpSkK2I1T5vOABMOwjnQahQHnz5RuF2fUISVPwcd0L5WT1q2BPTrv+P
NTDWsQh4OP/SQYSVYlOZMAGInxwaXX2pyCSzJ6HkVm4GTiP4Juy0UIYm+ENy5/4+aMAO9eJQXGCN
5xFSsLC6i0VmPmlzKz/0mGpe9ShytqVjdN3F4lTTvKWd9pcK0Rkw3+1jes+D/JsVRZqAlbMrDbwV
u8NCAO2Tnht8e0MsVsQAw0egGWTAyhmmMJ8px8AxMBI2ZnT+l6nm8shIk0yI0qXKr54FmbaRGEaH
HOL5cxnfaCLxex2x6Aus6bEDMl41tIbl3XtTIRxhJTiq4D69MViNu4eqkxR29lLLGzjwqKm7oOk3
sjDV4UNmBovnJ9JYZEY5JRgF42e9joQU7b7H61twqk4OJKQi0NVluuMMke7mcn+bOkMNew4svwuG
VybkDLpJjnOMi5UJDBqbGX7EbfVz6Zty+unmBpZr6NZSiqWtzziIZkMW8+LTfVPHgNX+5neRs8OQ
LZjcE0EABtLVUYM498VXc3mM9FXBfjIeBgLKIA83AveUGLwGQQuhsXazQB7HGE0SwW1RE/GbMSuh
ks+9WrQcgzK/BC01ptbO9bTFjyIcw5nNzYFDx4QFrkvdsdQ7jaQwaMFvNEE7pqgkEgTZqRyf/U9d
ewtvYqHQP5DLrw0WYzUWp0tr6898RpBvYx2PSl3lex3dXkTFElMQmQ/RqoEqtzAA8XxTACvPIQUb
KhLSFEgqdHBCy9BHI79cmPez6CPh2Gmz2gd37jRcuAG7KlYJCg4Fyqm+BK1kFeJke+z0bMnSJuUx
9wh2EC1YdJQbc/65tAT3qukjDLEK0vTV8Fi548HCP96O328dsGL1ZU/OUqjuAJ7w71+iLY4irZwW
tAGSNOswrS2EXfIKz2jG6S+ts8g/SmQ1OdxrWjPGQZvTpC8jmO9zTsh1zU7PJkZZIILS/FLtt1fU
aE01+0QlJkqTcfyNpMejzH7M/ovxdBsonSXavonFF0wmro0ugPlG3F6106sbDYlCAZKFiZrDPadM
zGVHci4LHITHbfpDzOAEhT8CrA0gkh5t2sR46CzT/UDlF9rsmJL46RH54X8+dRmtF/mZO+Tukaf8
1fCzeDPVsKIPu7dtO0SdfYsI+4Y2nD69cdFxhjT4CPxhadKIOpBe+ES5z/LZR9bnI3ne0fuWKUEW
LcsfWmSKtoZdNxz2TfxKeloT1S7XMKl3RHeZF4yREtH8hODWxQ7V4/pu/sIn1d2cI42EdwzANEHa
iV4a7NhvtLvZZfhWTitQL6K5hq+g1dUj/eMFVXoccdk1/sLGwj9DxqV+p7Ra5QzlDSQ8riObGnBT
ICvoNP2ZjGXUQ5EGvd44qkd8PKBvyQD8XR32Eqxn5bPAWzMXawZIqDL0A+Q7gkgGbtJnm7KKLwv1
mvqtUZx7Ks1eSnms45qdqapkw8f1C5hRWOkF/ScT4gvaDQG9XQvh8JF55VOAQiuv4YOuO2Fe4US9
YsGPZnOEzpSmUu4HC40IzW+3fDnzS373XN1ApqLZTZwcoVhmD5q3Tdr6hH7VbFIMSWNEfOb0Bxax
doIniVz8HgTovXq4f0iiayA3bAqs6G2CyTT8RIWwPB4qOePsCMOKoeleyUefgmI3EmWVPaDywhMl
+tJgk1LGmuaBV2NKNV4llVONGPp/GCAtGR7UNcG2C4jbRRQtZ68qYBM9YgMVPHI1g7XJi0ajUXg1
2uwY/Xp0+h/s9NmNj/ida/g/EiNnB1nhSLfp1Phw2/Tx2TRYJCaQN71qPle2x9efHX9St6nD5xc0
Rsxu/zIUotT1GcShm+TRGC7Fj0Ss/Np72JFs6QmefS23fQmto1yJxrXJH15S2ZOqKWdRXbL/nxjz
HUG/EZYHs+DKml259uUTbVRY6ufvOi5RuHRyZmr/8/t83C/BJ8FlyI99OfmHILJ+6OBZl3/2j7t4
OnYXWUMJxxZIUZbAQCjbGc3REgBhszWuAFaeDFf9JYJ/xlsjmm2LxuB0K2XNFzsacZllQwdgIwfH
dxN50bKNFZDM1OLgAhpWf4eKOaKZpiNtStvj8RiUhMTT5YM4ef2FLDz2ftEX59epkdFcsLGbUHsG
LDjLyIKnm2eMc223f1i5madfTqWxL17zgmCdAT7nX9DMG8unoHI+zlpALkkQ1QPiTcoR+wNNDErA
1kl/EgYQ9HMK3VBiCcpJigcIbQX+ESC52QSPGHaxyb8TXlYzLdvoRenlHwIa+M0fYuNMGBMaeS6x
opIvX+kweY0JDej5MSoGDxVrY/mbzeLgKDKSTvbtb8B7ijzizV0VYotQ+oqUpsd6GBELJYYZ4GUn
4vO3+Fg5jFb7GjgJNJdb+e/IPFXsAkqr2OJLaefY4xmDg5b9p/dM/59NaM9fFA9T7h6NT2ZYL1cF
Fs1yJNswTUbr3JZZNpW6kxCD5XpQzypE1iRBaOHSRfj4NAQr0Oof8pAgtW/IVi7cS4XIiRGyjs35
HIaFcDPoO1AyKBZ5EokpCj+TdqOawmvYRl5PYovgfD9jGs+HxnrcNyZ/gCNMFMKqUSsqfs1f6QAO
XxKyhvhw08lTFRFQiqtCqGXI6HTeLKPHHWIynn7V4wPFMn0Em2I/oMyWwov+1ZqQ17b0nW3I9aaX
usdMKxFMizQg/xEYFiwTwSiXIc5p/KlsK1m8U6VF6nxC5+uaVnxbpeY19rpkJqIvGZf6hQBN8T4j
+nVxkLKM5n15sFn0LEomG6ebQoGpuqoFPsDRVmNTWqxxKdjSvu/df+dUO7jy0DE4KR72WUvQ4VXq
1ip8nHU+RsFRyZ79535w90DdtfL02J32UmNRs8nATu+Qnq6cB9QBJKuOejD++hJ6Gemi7QhFkEgy
1XaFuiY2JOLh+EfDxPJMaQX9n4xHymiyQUd3KJn0B7K9+KRzfkQIVyFO55urG2iCYxcgC3hPajqJ
7tBhwSob+v//HoIuTbUz/7t+5q/+YImYc57fsapNUoFw58cemDSeZRTcpa6vQIbBgxZLZITX32Mg
maX9b3LHD7YRX4LeQ5pxkv47EFoJ8RXpTeUnq3tkzN8pFSlAu5bf1AOJMUew8b/WVgKjEeZ/jbQZ
LOT6YgbUHPDgfzoW9/uJkWzXZ12QPG3KxqGVa9p7FPrHhVlKWP1YH1uuvQWBmaVuPU2grs58MTi5
6mDPS4u4Jm+UgnQooD2X+dyWEhrGoIQiRgurH42TroQElwlSIEDaxzMA4eZVbe0NBi4qLPnYoqyT
xasqY/upu2z2BUMAemqTmNPn4nuauYeivDQub56CoiuNH4IrsH/40mpPX+jJ9ZWsTVtAdQbUysEH
66jHShLFz+AGo7uOzD+seSuzamaTDd1I7qFiEk/SkQ6xNqeOfTxOX/4404LiDA/KE7T6OKarIlU2
rUmKXWtpc0oBYGrkMmKAehV/dadM7xiHeI4j6iIuGpqRZKFoJ381LtCbwnyQ2fAN+MSdgJ9zGnF0
xSY9hvoAKAnElNnr3xTDR09ltfnxgErEXxdFCayugMWZyO5IdYrNf1PmrI6SNZKlv/COgvFnbv9Q
dU42nGxdacd4luiEDxcZa1lSye/ed6JsROWw3O7glax7IjxoubF8UKtAN+07+SBjcUBjsbRTrpgo
+JawrulYmh/IqFpIv67n9l21tCFgSO8zUU6rLZZjDGhRebke+XUxetBTH78Y5t5J1A9lqaCr/6l+
nYLmxRqvOZGMszYoe2FbdQoFGcK6uIpEkS/ODqmjO2hzGVCf4F9yRuCGB4hQZeY9H+zazDe8EWLw
95G5wZTs8cZTA0HazyQx5tRjSowhYVoCRtSMKr/h2dOsNSGoB4U6Lp9nhkf7OFDHrGE4TrzvMcMO
ldkjKTfHg3KuQpQK7Nlz+7or5n8Aa3pddjN90S/XTlaQGRI8vGGepvUXglTcUxjCWHnmkwBEthrh
Voul3TMjOqv7BkYI7qZNbC/9NBLq2MB9bOqa9uOdhJZokE7i4mtJE+98kQAfXO2+nEu7CZtjGi+J
gg3c7o3JQEOx5nZdl08WDmiroDwFc06BVmF7WqmmEbhjDu7z855u2K5Lv/w9ebNQh6AiXJKjo57L
9Rrq49jFG1HKZ06GneZMUDMudLfNPEZj67f5vCdYTlA5uEqN7U2iMnGoSibPGMqwRg2gooV3aeFz
HlGqixDJSxQuOHPrR/K+nN884fpt64AWLlMHMa2+ovQ3zDxG21zvOs17VVZANoF5s2pYHHjF1LvS
y44qFYhKFQSJA1317kFaGN6i7t8X9layrexB71KBVF8fV6fkxxGs+d7OODEz+Nwg6LCW04PnBN2h
ydi3VRxTYeKkUEBTiKOu/GU99jsW8t+B6fX/qMm5c47nSS+OB27bfyxOMtzXNVgZ+Y1DxuTBK6vv
Y8CLKB75105gRKVtyl0lj1ApeqQfIu61kXk+yel6uNqx7jqjDeZdozRIm5m6d2VYzhP8E3DsRdoq
0ItNubFY3AXB+I/SDS6xcdJPRkEBCLJVfVTXEzRiJVMMFevT484B0i+8UhvGIB0PMweZ2KbGw1D9
0lmxs95jqmw2BZTF3BD23SHsdlGuue2L60ecLBFf+hNcUCtcNBhDGUppAd93gjz16YdYQX9DH2vD
ll8swQEaXEmMZIQif726nd25Udmdb6R9cL/oZHwudMuE+YluXn/9fcrJKPJLRPnIGPhNO8Gyz+Ex
1+kGS5+bE7S5J2MMJX39iuQePErSMLIUsb/66Y05oP4LcSDMeOACXV6IBrUYwSi+sAQ+tdHnqNWh
OD6fSKDjEcfhwCBM59cowcqgS8L4hsXHlyzdUMilfeaVHsiPzru9CM4up++lKSpmazg0Fbih1RRQ
F1JM9NW65N+9PWHuV0Uj3zl2Yw4L7JQLh753u1/QGaeEexmQWw2l9G6Tha/cKdIOeuaaitaMf/D6
yau1LTJ+UHlwLafb/e57cp8bJHx4mkfCuwrDeIkqgHiRTTTJ7OqrEw180T4unKSSn7ONR+3NhV6l
+5sUOAncars6CqneYhiOZE7ZGAVMG9mSJe6bnKf3gQVLn0KHW9L/1do2XGPLMaitz1qCsAZf8no0
rFbvgQmJ/x4HnqRUKRLqFXb88RQX8+qsDUJp4CQ7DR4gbm/y0iO/Gkzw7ZoI7PcMKcq+vV5wfmwi
jYf6aw00pKcd5mCZI8yIKjfOwprDaZX28IxTO7yuusoZt9RxUNow+uJsdEKAQ6NY2VecUGq4o0kU
oE8PXsUWAT5WDmzLaHSwUEmzmoHbJCwWDHBeyVJ8xZJQnT5IXs1GdBw8nFWjeNGs0GDv9VD7DMPP
qsA4YJNmd/+rM2CeoPRwLAyVY3tLais18MVIXKLQ9qN+Ertjo2IzEgXAtTigtT0FIeVpe5MhhPgr
PzGcfAXhcQRzn9Cu6t/PAvzq/xC+MMlu4lkmzNTXl94FaivwWcnTnij5xdotRHBegcrgr1QpuQt7
umhYoc+mqPDYXJN4U7iHCurYdfnWr9rSk+Mxfl9CTTa9xT85ZNskPlRE+WKSDjUX3S8RoOqm5ayQ
3chbE7vc53UavF1KzCH00nCl/KaIa/B8UL3ZBlcjGSxT3SSvRyAJF7rr55zwEkZDoXwdcoa/6XC9
SNAxNIPWbLJWqaLfhe50K7YanaobyOrZty9xz2E1fVk8Zuv3f/BQz2OWhNA6G5AnFB0pMUI4CgXf
qOt/MO8VFI4IsGPyEoKAzECXm9iyjjEPdUR+tnsGcKKLVoHrYJzCTykWbNls3p3gHGGj9+6Hm4Ij
GWTGBpm/Om2hI1zIS/pImEmyvU4h6GlKvU3GXHpfh7jkfNH5Ih2DWwtHCHGn64QZdvqS65nrdEbo
v46TjZshnqcLTPBbfKTDNBhZK60azyfdQuVvXDWrFYjcO0XHAEnHYKMjfPo/zRtEy9Ije9lPavEf
OGqRHBpWXq0DyM0P5C3A7R5xzj3S1q/5Ynm52ikz3evP4UKeBXxnlJyIcePBcslcSVanEx6Tp+pd
emHyWxGkeTd1O0107kXF0erv4pr6WTFbbu4RaH+psjv54fAUbT9qoTisr7BqqxVLw7X2zmlm1BXZ
hwyHyAEJtbLiw5UCfwQPNbs06KAVdQm+bvRZ7Syyz8RtkPEcal3kiBMdHHQZ3+LGnrZQrUu9acgq
KHiKupt5wsnpe0f3PrOXWl7Lho85/x/cLvWCN9XK4jLOy0lDW21TsXC9N1metbzGUfPwHM0Ti2ua
QZS3pz1i0yeWpH2MbShOKut2+HqjCnP6maczU29Stayblg5q2EaH5fvg+5Ch06UMnjkHyBSsGVG5
XPV/Y0USYZA+9/lFty6JW0NddhJyd+Fg1ZwvMKoGk/Henvz/aasyAQXPSkXu/Kt5IUr1RTZp3aMS
hOuUPRVH656karqhL8M8rD3wd/HXuZ1hjUO5dGs9smwvZP2AOeHGKtANQkcaYAlujuhKZKMKZvZz
eMIMD2GPJNgVknuiSWlB4pINtbVjiNgXwDU/hiXE+z4COH+bkoEIzCWKCwxwofaaO66Khi/5yfQQ
Bh+K582FfQSmFEo7Dp+AL3EpFI29O6VXVq6KxzewHYJNYyFrKzRIQScHg8UYER8T8sRwjl8/izON
mvuNaxsJCOQz5lYZa7sXsZSpC5PJGdlqjixoyvby+Jivi8usdphKtRUPBa9aA0Zvh3YnriAUwJTI
Hn7tDSyF3cjHyg7fKHdsg7EkyG3R/FPFidVHE5yMgrv6PmW/pfHFn82czl/j5e1+5StElJFg1fG2
VR8ZSILGiEUPfN3WlILYnLvdNd3rMzj93D9L3Ec0Ylw04ndNBVh6WLIHbAcJYgxPDsoYMK0Afe1b
plITP5uLiJEcae6fHINv6VL1wtNbGKrKULWQgHbnC9UYqCesj86pVPGTS5SblwXokLVLiUae/cR1
efXb+T3rCL6YMZRuaQo6rZYsAfphEnDz9DhAKJqbSrHYZV4kLYccDKKDubiB6lQRlqPrdQcIe330
ZQ/BezNcYijndKx1KU30J+T3nm08keiAH1vPxJoODpN7OLe+QetFoMFRTRpS5yk2R7lU7jXAKEC2
IJVWZuZ+WsVo6Vp+9vAd/J3EmmgwK3pn2njUwQ9YzmkWBq5rCYv59ierg3ayPv91YfrFtykipb+/
BnBic2R1LL2gmGVTcKEmq4WS4XV76Y6pgvhifLxkZOiGoSlgtg8W5yZlJ/TWOkVcgqanie4H0Hw1
ymRijeiH2fOrd6IpiOowEBk7mYSYKe6HjvnKU+KNWu/HI084m32PRfo0tN2zamwIvNWuozwhjt/9
uX+OkHw8YEnqkX1yMNk5s/74Qf763D6TFFbZwVnFOXgem5oK09D+mH/qx5rTpj24bgUlURl+SqDG
sKzFShvMHM5LjbgO+VP860I9VyMTV26+Adhqpz+zLoxBgo32ieEZWever/bmXxNQc7L3SPXfKdNK
3qkEa0xK84l5BiiVxJv4bfwmwSWjwKloy3Ei8MUKQHevv3qCjfsfl/z6ZLHwsgqbjQ/5gufvjwFd
dHvhryXMbT7Ya/I+Ula8fnZ3nmL8tjWa534HVYlPM7ibbwTR251EQQGyihTBxQgjUV0DBTLlODka
T2v/FjI3iNAoTbSlTFM0hH6siT74cTVBDQrKd1XxqJjVY9HuZRHLNyEoSpHVrMJI8nxaKTyuBppS
i27qRpf8GKxBD3JuwCKpQfM0j5cDOud7nKFVXhrkLrLXbTcoensfYYHO43hoVSYWk/1EJTln0+Do
EpYY6Jyu3zSOUSq0w46N6MvA70VL1e023czaHmKmWtM0C+Mgd2XIru5epQbzFiaPAv9lA+i/vZL3
fCMDrTJkEMDE2YJcLTxufl5H9ZyiamRTRlKHoU6ukd3re7pDlE1RF+UmJnU99fYFJgBg91plqWGr
mzRsJXzw9pL5izIMPBuZ4BuYxDN+hkvqYd/kcNN7XED32mQKyhLCdpErJdvsSL4uzkj7vB46YaF6
QoTMXXjGrWL5Mwuxv6EQpB8xNHUfJTuJQVy5uJpA24C17azid871bV7n64zbl2n8zq0QDo6qrQ0b
0tsgLpDdoExaT7pPRXl2o4ehQmG/o8k+29T1Sz6qvMsGEkRrDEgyknIUlt+iDip8o1I3inIyKRCq
RuQHGCnOZhlKcI7JASJURqm/qkw5UrqsZxEh1YZRpky2LVuIuRq63YHKMjUd3qprwse6H7dP2BQP
xal461D8J4GJ8pSQ3QtRZaEsEFwZEda1EVusFioS3aN18KNy2HVP8Iu/UBVUdLsF8Vkua2qKCXUF
crp7gh/dIH2FLA5lrmHEbjyLeeOBO4zWL0z5vL2PxEmmon/yfEmKleDD/cgBUqKl420uWuQre7Zr
+j1BB+PJni4TRREEbNFtW+aQ2sJSbY4f8BaAgHXsZHFwZ6EnHTDuncz5QpIsPR35bC1pt7b3EG2l
5b4rjzb4jDw/D1mOelW++ReG7lJQT2cIc690Gyn4T9iwJRrDrVyWGIP0CDvEboAAzk1evUlRlViW
horCiFzao1sfvh41iw1hrFhxfzC/n4ri8rSjbKqQRsD4Vkiqoo2jBidpIJLk3p04wC6cBOX93Ygq
ldnurjK2TGRzukeQa1T9YhH48kjX7/cWJbNyua1Ga1fqvjIl+d6ClkENf4reLpa5rZPNdLKi0fIN
g5tNrot2+qljUo9zL+vRQ/EOTYYiGkB3B6KejNDj9Ah9F6+Bu0dwe5aM3v1maUa79YIeN5ESI26m
JHc7qkfQn8FTw6IvbdGGFMmEO/a127IT6XEx9s0+Swg5YGMXT7aQ17wKqUx0Qq2MB5hA9dIKEZjH
2mX4AIy3/BPRTHX1i7ElNUainizwEewPE5+hsHodm0jGk4fM3ZVokK6lKsXXr1sDiCFu5ESM4qeb
INCXPeaN8qgBjHwtbzHDssOhT9bAjDTcipEPY3fJgNC14hUuhiJpbVhSKbJsWs7r3xFPt16BcoBj
SQL3V62UXBDz2Kzadq0yMiDi8jAYZD9qvhaZQ5FrFk9m4ux4duVGhEbX6b/LIWO7RvS57+qv1Kn6
4ILrmmKYB+f9R4Dk6IBkHkds+2oHnMrVCJ2ePZ+k9e+82mPs8IQeVKSbqnabCrtXXccl8RoIlyUa
gq1H4dW3RYcscKbsOyAbNUmb5+VKu2TjvEgNVL4WB0BjbTZmEgNCIrAAsH4Sh3Mvoak0sRfSJJUi
/NLvbqORvhNl7JnqllOtaIQb06/8lw/PoHJTKCHORNuLvAeTxjIx5glytFdlvYnN2PxQZld6R4yj
7JIbqv5kEp2FucoKIpz8fVawoJju0B55Ij1K3fdVFrD2mDSTVO3ahiyZjfKRWJGsS4u7xojIclQg
YwS6oDZnA3bIs9ik4jNiWIGW/C2XeOxorLBXa3SEtWBCJkx22edJhkQVxJzTFrnM+VXbFXYnfYe6
DhxBmSlEH9tSS3AZQEtNfMEy8sYGlEHd8QywjMTyXAOStq6UdcDycY3JTodeYYPAcmvbMJ9++1b1
BnXUFah7+ghJjA3LFbq1INrZlqoat8aMEyTQj28+IQkxWmQrKwH8/vQBhSFkIX4q6Ws4c7TcHZU+
XLtPnvmFtFSewot5HLPiWS+owXVhYkKJaKuRoL3BgiS2NMUT8u9fY8rlUmSMbiMPIpuGKwUdiOh7
o7bXJWlryduO2ZlHsrzKNV6SuC0FAqF9wblZtPRyADkh91XgDP4rS5ZYGEIy5aAV8fN/Yx8pLF2l
md7X5aTXQ31wRqkG8wtP8xm7FpMV2BX4ShI8SFNIxfSEbykGA8QidADKYQnx2BzrtHmGhwE2h5yN
efM0uLYiPLREgdYiU8rEjvox/2SfmeNozdhtMJRQqgApIDghgWqj46agoFjcPO9m1IOwGWCncpMO
Hwl34X4+/i0ROsWgEbwT/lS1d0Ysz+mk23OQfnnXRMqha29SzO4OlyJ1AvheBIZjoWMk+sb1IMd5
acZPhQgU1G2TvedIiYr5x/5r1V+wwJFpcoLhQQiRTpbwAHqEfDowusLNQAjSR/NWXq5+4G0cyMNq
zZQ2hPccUMIQIOCF0/RKaQt5pOv7Huf+WE9+IBRoPPlr45Er6tBCJkh4DWWeFBER6NrjDobpME1b
XfaN6Y/6Ik9YYIvetginJIusqSWw0RiJmVJzsAq4mN4mdM3OadzUdoThov1HgcGYpjFr6oO+WCTy
eoJYCHsZ55S0QclvWiBFwvu8sL9ztVw9/U7ll6zSwW2NgfgI/PJBzGdYd2qYtBkimpM4pRYBxaW9
oAAdWodReBIctjqF9h+ahGYNp1QA9/edpj/4Lco8LO++y5hGL5C4eRjCLokjfZQP2era6aF88E+R
OgPL81F7fyhTSIur7uMysk7PIoF0fNWpo/LD0HH7unlDoJL7hpxjKGkQsN24vzVe2ABGNuybOGI8
o9I8nCrGlAgK2IbGy2XqxeIs976oVxQaLDuy9089R107GbztUO3hICdtAT7y04bVlRe2XmBZK7Ee
5HZRVvaH7JCVnwxUm9COXkxKRhyi6VWl7uJAmuM4rXaUAv1gYWXecJ/AHWlpjYUeUqCpQ8CTT8Zn
ESkobgYDdunau9mgsDS1pVhSb6ou+KdoNPBaoY+e9mNnRWZ6lE8EOF5Ckak0ogkdqGqk4AG+nm9n
iG382fKJm3tvLaLnny+hyT+3ANRUgFEDPinWKnhbxTpfRTof6CErxoXGIEy9Uxu1bzIEaGQ2p8eH
ohKgM63a/C766FRK27Gj/jQc7iejR2QifJL093ygfzztLvzrDHsaonLjRl0Iw3cnVVC7tcUQd+QE
bXqRHmxv99IOCBDocGA/qHJ/svpCkI/+L7QgdQhbxO7b9lhPlyEnVwuU+Sbn8F65txBOxQew1iDr
HJvK+1sUwgnJW7K7MkmpqWYJPmjdpwe9c+mdT2/F7B8dVDrrUBR4UYL/B7/1dhkUyHHiEZsyL/Z1
27ZwDgwpiKYMP9buZdUTVyNreK3L7IFa4mc5txaSwC4K0DMEjOFfOd3fXsnjH3fQ14JHe9ZMo72z
C6lmVugjHQt5iw6kguK2xfAQSpbgVzquISEYScMRBhOLGzjEBlNTDJEPGSLhGT+XBqfNkaJaAa/k
4n0cID/GXaDhGfIyKJ5wlCOGK65ytvqmw+AFtqCk/nyV2olJgkBmUbudvcSLJQa8IKaizADcdGAO
uo9VwxL7fchY5wv0neRS32sgbKdrvz0o53YjVJN2nAz9fWXzg6EThJtoiykd3Fvr0fuXPAFtVR+j
eGPDyCvsQPF4j3BtRQAslbGXuGGwCTxtzVd6M45rlojd9dQkeIK6Pn5DpMjI2jhxFoemS5RullL4
B6qE1ndrXkhcX1dvDt7VMRzdUj55X1zIiQFVs8/JQpssJIlXxOw8YygbudZC3DJyGiu3sRVlMqET
+DOlKqj4X53/AAEpss5qaui7rzym9ahiO2vlyqV+sJ2fp4q6J7WIqx9A8vYmaD1iaeiUEerArcc2
Sku9QyKlwR8xahyTUurGcpWKThjiTKN3+PcYu+I8dBdXVC6VYn46CGzNRGtO4ZCXShAtiV+mfXH/
QBwV4+8XqMA32YmPbhNZBtRianUGYzREO8aGgTY7HPdnesE5iYXMV7g3e/JP+y98VsDVmqLZJ1Kt
TB6ARXLJ0q9DPtOxyCTyVjiLXFGJPVsfDlOmlkasqWwa+pUmAjYxLeHNREv3rOn54lhM05yimBb0
STNnXz/NXWZB2++xI6syuwCxEcooHYzqyvVj5ctyXFwfQcVk3fhudnhZpl1v3a0d2IIqtqhSDEEI
zY0KK7BKKhlPGFIp+tkq2FgJS7UQetDPAsPDhGypWhuQNoHDxS+LwFn4E+NIysiHSIxIdkVZER9G
p1QRZWd/oR8x7CgDjVA1dKjPgqgskdL6UE/rbVXMofajZCXjps0VQMfD6MUDR7YPihQ95SJbUL+T
oscQAU+ihL7mmJQEcebxR7cnikHDoC0idzVUIVkJXXtJmNDCPUabMoInvGI+pks+R21wE3iWyjk0
k5LWV5sJ5CTdA0eLrqkd8klpXNSxYyTdsGgoTsi6adraorqTFBHmyX89Zc6o81VujF97EO2S4RHB
LsL0yLuSr63W3jdcbt3pmC5qCu64XTwvF37MCP1nqrDNB2MxvzHjPBJMaLp1QHDJcRaHsby61Jm4
IrXWiFGp5VCxdYO1Olv+xK7pcB4Gh6icNNNWWAsL6m/MiFOPlcOVg2lxZTHd9xEkldqzgU0ombQo
DlsAxSMMFR9dRiyPBLgzGNZfTkRSpI4VQmASIVnlVJX7XWgtqGpV10m8A2w7gkaeqQZ0M+2//D68
yU1OTaiJWFXeby5MuYwmQIWnqwkg5sol3qxcDuz584wEcPFipSX/u/YSBA4gPDKrFAIH2po791kl
4grUMUqvHKb2gE4EcbeM6aB7ACTiomt9UkNnOX+e5RbKHb/anVaqTBCmd8S2RjgH3gafCBX4w0C9
SI/Tv2zASVKYRQMPnZGNCVVxZJ0yrquazV+gko9NwRNkJNp5iNq23HDVqIg7mYawudrSdGUvKNA5
rmNBkoAjO+CGVN8fLDF+WkPVwFOgnvoL9TJ/S5xcvZ+JsiK2mAO+NskXaTEP0LW7ZoF072ZiQN0z
i3aIimul+Xlnk/n1FMIoEdt8dPHfaTHTMOCyctngfdqtX9l1roCwSVkp2a+K/qC2QioMlsVdEKo+
5u3v14CD1t2Ac7F65lJun9GuhkQk8olrG6Swd7qm9uHntRyADvWOKXvLPUPSLXT5UvKMlkBF9Dhb
S4UBxsX9K5XwtOcqUM5zTvNEvn9BWJdAw8MgVVQ6Kzg36Sd8d7epM2RwxO98kZ6nsC1owKK/EPDC
MwqSLfgbTIYaSrgDy51wZ2F8fGQc0Bqds08vAhUCXfRQqP9amRwniCfK476U2SORf2q27lJKxsom
o4nVstQ+B58UkWY2K4pNsLTRA5CNVa/qbIkMCcy7pQ3/H7GD99lMjgrdQSNWqFLGJM78w1z2fcPk
TQ/33fwwEIUl08KX2jU8xtgKmaJqo23rmOo3iZQsleAFFxWFhaO9Qmp5c+4uixqpa1lJALBojyQI
I+5ADw/AOmiyKyLqpIwuQaLCR83gpz051MMT8oFZRFIVWyCfFimazuLM6IH2QtMyVdxPeieG0p3J
IxUEqSJpbOUXw6SqUzdTTXMS7PRO/rGQWuuf9cMgNJOQ7ej8Xs43P46Vg7k8el6V5Z553vDf1A4y
5Yw+5YKrjrahRZab7AUm5V9Okvr48HKiKz4uW36SlrkeHQ5UMY0+bTpYwYz4vmCoDztJY6lMhQM8
cW7WlOB9+comytqkB9XUfpA7PgrIuAXnIuTx9zWwqp19TBvK7MVg2UEK75wThlvtkiICZO84B4ZJ
WOzAcsM2yTr35MXOSrpmwxuAWpCsShWt6AUZPxJSJqnVhjYYVdUkCn6ZEM3PqkebuTHjc0khaYFe
hclutvfELjBtIn2ieUU6dJTY0biNOWRpXFki66uOMsyA06+L9fXg37vsg7P3EdECXyOhiLUR9Cvb
EOEDjcEslGutyfm09phTa7vjOlXWuLgRr4J6iMpJLXe9E9O01KVKdhdx6+AYr1+/qGT1QMlAxMpf
jgZC8BH/BSl3XkXw6lUixeUhZjxVSSqocMabt0jF56ZWSDCGWNwIdFTii7HVnCxnkt8XAOy+V5LA
ACrtD5T1QPbFRM8rI7JNHA5Ph0eGZHsvLm4bYgwIhSNdWT14hRNINBnHC5yUMvmtlxsP1ofqCKeS
NriXn//KXt3w6/CkvXINJukRdevpbhekD7AK6ro4+i2ZpLmQxJ/txqbxFjmnrq73dlU4Iae8fe2C
/OPO2m3XTzHoPB24Ynuax9PBTHZvylfkJ0Pch5DvRQJv8ah3ciV2B90O61z0Tw7jjJIBe9Kui2hI
xx3GTEndOgKV/arv3+5193yMS4YFlbXLQJcrUK59H8CZEUklYn+e9fI+GmAA9zJMN8BD+fvpM+un
pkoqSwkvo+CtgSBej9W6hiJKoS17LQHyPYsZOqSRW+V1U5/5/hiXuxgLzm62aAhECOimNmJ4YD7O
+mMbHEXWEXhWAigD/1uYzFASQWCZm4IPStAC4xqNR+z+dQ+NsIPqSKhVdhvNGUaO6YJs5xovLhvd
ngrSyx2XIBV7yHWtidbulE8PBPZDX18l6muKXYqdSFIU0RZkytzIlXcFcGxJYFsSUWiNSfEUhL97
HX0PN8PABBozzslvZNVHYoVWO7Z/LYktRzdoey6v5QbJFXRqkgCvppTC6hEFD6xOvcFqmO9PYOjF
WkVx88d2XpKeoWdJ6YcHIiVBBmsgN5Q4+wjm69H4nqVxc3JVP24BYyPM79/+XUTngAfQgB2fSdeB
jtakNvcbXbcAeEn7y1T/ZhXSqbiSjmeq0YBAaSSTkbrcdRjAb7ZBbpv/Xup6idjHNLq4l4tOvf+0
5b0IcKDPBkrARWi+7ldYUHs0uGBrq431IHgXTJuDrnmsJOmXguHgCm5VM48xGcptJN7lN9V6FdCy
vEiU9x7bjY6BcXUxYX31jXrkTy0WJTc9Qef+36pT6WzbRdR+Our/d/asIhHB66hSWxFyhlcAg7g4
x4Bm2YnivzuPEgykSKvyDf0xVW+eXKz486knRcZ1EaT6nvWEd0GSOWEvJ64FJqGhYF9iG0ZsynFL
eVx7fZNKehMZJuByqKGuhFZ3tM9ZzTGfmMiQmekThsDfhtJkPI5A5WmL4EcILCm1QQV3/rV/su9Y
K9P7x93X3UFXC33uI7Y49XPBcUiqbX5m3/uDxjeiIMySEf1xRAoBq99yP+wOaKs7buH9Azo/SYZK
1aoRRIqyuBI3a0uPLRkDt7O9iGeXVhe0eM1nKAtGNFpSF0B+iaZ2rfj/tdtz/YPtQFLEx4YltUrA
jo02putmXwQ5QYnb1OvpEBaLiKImsjv2hjQ1/Z/EWTHK4P7W83UJlyXR3bZ2rENqWVtGQhQiVa4P
UpXSQ9CFRQV+koD9PNgT3t6+Ppn3sVjMUBiTR2j1OYilny6xLoQqL0LZw9FzWYNtoc9U48NynijK
4PSWXpTf9qnxMDG9CEK373o8TArpvPWzXuStzFOD6MpLiX3k1NSadL/oOl0OAKlVksmW7CrSY+PR
e47bY0AWDxJexcsv1xMRxBBEzzItimejv3+/CQd1RYahqN/a1yj2cd+Gc1ieFxmqvhW6vG1tHbTy
XIxfIwTxBBhD/7aKZOzisdtdjD2aCfcL2+S173TZE9wgvbbpjUmUARdRGzwNmhx4QUhHBKuD1/AD
ZrRzVd8PYLhXJGQ5zbcSN13zJt0EPrZRvnc9mCEf5ELbLT8ZIbcRBFWD7FlUl1bKgHV1roeqqA7y
NxbaBt4YkdKBuqUWa6WbX7dAwhoOWsmQ5UQ0RiwSNo0YB45AA5KkyT5i502EUt1SC1FZpuRRXGt3
8b4vXwnDXEQ6DQH9wSD4h1+4RFmtY6IKnIBV0JgdLUjegQz7a3il+kSCfgO4LJuaT9qxi0p8jRxX
ca2RJsr8oss8PZIeK4eCFnynVK/yWSTt6i/zDO9Sxua9D7wVRjZ+830GQaaSaTswpcvSNlsv7U80
BkTn5voEpQNffz1155yAZoloRRF7Du/hB8t00UWKEwMb9RN/CzNVQwPXRZyQIb6ZPevqY+I03mOl
YWnPMCcCLjSHF+6LW9kSmaznT2QR9jD+gwknAgK5nZh8yYZBycIX1DHT8LU1cJO+NCJwD3PKR4mc
swXfP9ifd0CA+dGB6plfP+nagVcwpEmANZxG1mPWDeAgtgh/YRLv2ml/nsWhj0oKpEup07FGcWcZ
Vn+XVDpC5w9vvCfbQ4Q84FRQ/v3EhpLhKHcixzmR0gH/Mus2Hi5B+yVTl2FspDZGNzvOSGmbZZbZ
ScEeouD+lxFn8hEhLkvxw7XrWfTyBRtj5ngSuWmJPGC1HHiLb1yHNB7mpSBdkDwDoG1e0hDak5qZ
YKV8ch8CJ8OtsHP+p+LCDQXsDvTGMdSUZRBfnw5Hqrl2vrFVU5MfKD9/6PlGJPrfJ3NEDDEYfEMl
bAq9GiRVGnfB1rlR5A4zbnHLNuROiGnySuYMqOqsbCITsmEG4m7+qwfFieI5aOj4NX8ufyLqu3rB
UieMiWBoNGs+EKmTt3LNUmBtyxrXo5uEilAq3MLRF2HKTJW+ZK6/e5A/t8nlszEyz/EPQloRM9aC
2YuC/0+aWRakS9OnOCIaHbasWEusajdMkxHGpcwrn53FmUNT89DBze9GtdaXCcWt2g7USPxA9KZL
ooyefP/dfqaNfCGkkDLjCHj+i8Ais+N8iQnVt0JcSAq7BhmtNssp4cGPyoSP9ooczrZYQlnVkpaY
kZAMbb260F+mjxTFJKL/dm3o6Zeejzh55dB9DNRCCf6hh39B0wUk8nuciIbag82wYNwi8wvdNIw4
xUnAnONd5xqV9aB+J0vZUI0kuzykomylfKdxyfl/uIlHqbSohreFa4+x9ZVcMyHVOVmGLVZvVG5A
oAlhlQgbHJ9m//oneSYWDNbuR9J8HDLVHVu+JLFyIK3SoSRhLxjqU+w/iZMHcsXslwKkv+mlZ2CY
QaVrWamA2cEzWLgDQjxd5ShM90NflQ10vhsSUrgWIT3JCezYT0g0FaIlU3UIyR/rNZXqkWD77oDi
oi7f6OGFyBPluahiVykjTRPWELkXBcRdCtTAcNUfoLsGv4t2zDZxBRQqZLmDoFHsU8G4VU6iyA4B
KvtGDFTy4ckbT5wzjaJxIkdz94ySJA8eqFQVJxN6E3uVNYu1a+SS1HrANe9DJbeUtctMqwuiL1n6
cZ2P8NO36lVHAvxKCLIRt4Z0d8e+AhBjgm87HDGu6umTxS/Gha3mPgzjAVkO+n4FJS4AEtezs0lT
2P9/4Qef349OEzzFElpAbD9BawQ8sgGCEH/COwEU/hM1hP/wZJFreaY91QqtKUsexDH7PEGdIU7m
2C/SykeBJQICErzKiyhPpjUgC58/m9Fje5Da95QyIZvdRMosUmiFBqORg5PzY25Ku0LY52VlkoUl
pKZTfb+3e2rBwiZlfuu3h8+o9BbC2DSsC81MiNjTPrQCvv8wSc0p/Ue7Gow+SdoAoC5CJW09sfPn
szV23NHKXn2zRzqWqYz8z8RpSw1kZvjCVhUbFMhROJz1NIloL+pR81Z3gjopmciPrIqffZisNFcg
emhvJgyzJRWOpXEShFqWNFUxMu3gTaQYFVS9a2//mi5hOovHs66baqkFtwAr3mhEEK2eZmVYdixE
f6JmNOEnQcr1/yXtD4Pqvw0cqRIdMsV9gTe9uuXu0VUNYu5Am3uCJJ307l5O8w+JJQyWVMDuc5kd
AwVO1TBo5iIi0V10pNnXZ0pnrLxhZ/brqZUUJsIw29EZwoCSZ+ul1f2U4tSBehqz1QlnoGcFhaWM
KEydW7uBA+jatKhcD/iRxOTROAppMDsKPUp75n28pxshHjxpX2inVmpnw2JZqpBwAjXQVodpA9+c
AXtvlMe8UlPQk+bbm1AxlxSMzRG8WWO4VjUfIL7QDlVSReEPdBKai0IR+9wmuUZt1IXLHser7eMj
3kxSyM/AufvBt1Cwx9uqtJW3ZTQeeqLV1l7No+aioaY0HWkIaxvniI8RzO/wC95CnHIGDVh6mmqt
r8dC7baOL6sFq3ysXIxr9rLwPyoYA8+PsRy+z7jWT2rlsMelpKaDkceq4PYwMv5PtmOlqj+ZxvYH
tTAE6uLMwqs1aFVSsquxc8hEUR1eXH3yIg/AAhktQ+tjgxaTajIt3T7C+10IcootBOawL0mdG2qQ
tw0Rw8bij+tkPYWuV9rPmypCK5W2CJhBpIH5KsRRzsPzX2LdlRA85zWm+2/lYuE+B+HtgjB9dund
Y7PdufsIB6wA5bKkIgBF4PojiCLIWKC/M+LShKfXjahKheIKclKAJXnwx4qDZCXuy2ZrrqB3YmEq
IDhJqZmLiB/51mXW4RafdPnuTGHXcm9H4iKW+FLwt/dINh2yoxu4PBVkTCVUxxgWhvDLkqz6QJH3
tdZz0nOA0OHOT4mTS817tVF3BnquMn4YmWcJPahga+nOvgHcVymkHMMlMPDouALaxCmyISlNe1vy
CAzz6JJ9vXROg9oL1wNQvR9V6uatbb0tTv8MYC9f0rx17StcNLDCx4jftN/Hxed2FDV0LjLEXkjS
j3HGmyarUxfZDDSycD2MjmxWTxw/8pW4SLGOMuSY19pV91hB934AzTPI/dQJkwyl8yWCkCJMCu8L
5nDRYNdpOTX/l1MW5WaGMgFChnziTSC8Ola4VPUh0CgeIkEv1xiazkxL0xQ2Au6O+WO6Bf+nXQDn
c/YAN7pKyW3i1UWrLqdXg1SP26P0MPz4HwKb3MAn98KKLu/23Ow0A7oTAL1Yp4Fju6xYNI52O62A
ZZa3xTLyDBCEzXZb0y9yIwSQZr/tQJaWA5wv6+yE0GsgtS/8mQgfsYObbYWKbhMDRAv7ZRJLnps4
EKw5pJEdMY7UaO0KKAkNtPF2vo0syDAAsj1WMAxoGYLISBkqZjhgI0y39vZdeNK/D7UWsosHG+JZ
FyfE3GcnKHLjJjADzDpFwcssKjasHibrZDF3Y1nhW9IbuQKwHzYLca9MDyckcetKAcviEmW9LBu8
0+n2K+xDtRNcXUClb2N7uPs8LLHe44C2O8f9jPQ7eDLxAp4Yyuirzl4yWg5lqCWwj4Ov4lkwOmTH
lGQZyxy3txWEEBNIp+mvbrjPiB52fycwMdhdgQZJFz1JImFIqmQB4UIAn1YYiTv9wbNExvq2sjKN
dDrJYIF4N2VvIaAAvQdnBtK8E0+x76vFBpWOre9XNVOUYABA6enuqYRYy3q4dWHAt2+LNjoGAFV/
OJbWOJPalvEN1RPhGYVJRkTMeJfXMm4BozaEM4HCH0Y58c7wmDHEapCxNCTjIJEldn2nwdA5HzSY
6XmGr94JYfb+RWk1C9QH46UAGPq841syd7eDWDKbpYvs9k6Wh3OUcNT4WlSTSpVaB9KWePiXUmtD
TPHmvPnswKz0PL1b6tbov/cKVywEvU98Oz4qY0pWxnZK4u5BmQcv+b03SevgFHmx8Qfw/x+KihIS
pGz9PlRDS/bzE4EGAelfmpdzK62LObcxMAUwOzi8jPNCA8ti7yX8uCn9STrEgYcKxExTMMAOazKK
s99bxBuehk4M9Ca/ETFU9bGd5kK8G0VQkuf7va9vKldtJtGLVYQrRdfjejMuJU+P4R9sDiZ6qkd5
Nz1cSi8Le1qKDnmeU6ny2jJ5crg/nKyWloxo1kiaZTwTpaUqpA6ByYOXgokX0BAVxqA+npWFJCiW
A3FRyw2yfjMRQSDbR71PZpqlu9cTpG0JLyiOgBfaeBttRu2sbiljRZRHAudGFh4XkAhbKmkGTGxA
5/WcaZ0QAKi+xPSp4m6H65cxJGnNhMB71DtK/eJxMUjgUqrTqfFD20i5XTHAL++QGH2uiJzpEZfi
56FpC1xAKXCT4/EfHA9R4xf2+BOFoKRX/wMYriMdTQxGohk2QZlKznqTx2A+sWUktQMtqZ3YZFt/
6KzaDY0Ckx6iwNXjjuReeW2eTxTnAwG0Rs/0iFOD6hOixKjYJIbHCBDI1mxF1aqnvC5Nh51QCFWj
hMtfsLb8lw51Fh+FjN2jgdKcYRg/fR2yTDWb+VTQuBN2EvsyvEVPRJRYDXGk25RIbzAkK9dOoTZm
M3pYriJKpg4gYtFPeL96IxhptZgFg1toMsuFZYEiH3Wg3DrE5y2rolXIIeUCdUqhvFsxHjUHUkGJ
kxOxQ6R19pM719TPOEpbDq82lFoDlTfb8UpHwkGC4ZsT8zZE1kWVt4FGzL2clcJtkbzGKtK24L0O
YkfZhmT6KsQy3sxNdhbqxdG4RsW29YuleWC08qHd5XvMsflROV1ZD0ImB6F3nAah1QRWqVcbSUEq
mftKz2yQlwpNgrpIZoodbkQUhhGEIY2qIKnp6rCGD7rrtLsQZtYiDdTTwqmt5jXFf406h8f/2jba
01VxsFlXZZBNbLn2gM4Mg0brlChnMiWTt9jju0FITf/GJqwQWx7NgthOvIFgFfIDWKXXLAIRFD3w
3POoRJ3JAAHBAF1Wi18xAbURbMC6PA+t1yKAoKN5sSWL1cGr71Ohtw3mDDllUyMmQZOU4LeoXd0c
sejieSDp/xnsd8joMz65Qpih8mBZxWuKqzzVPQN4xYLRmE4WFW3Oeozrq/oTXWHVvwkzMr5jvM5z
RJ+hyYqG84hCtXhLlgnk3KEC1iFB+RSxjDFcRLvZe6CXb8EX3PS+kGuGqFUsxxIB20mCZd8Gc9y1
T8C+17kRQBy0PjB/ohDrwSDm84q6R7tu3eVFlRY8SNJGIn6OAdNOWtnTq5ZA8E3TubNQcDGkO/bO
Mge2fK3m1skt4fQhcUfYuebPAMoNdEEunpZaLQQglyJEDblePhfBDzL+u24/xSPMNvJXrMpNDBGv
fcBzHOx+GQLOttVuTBcrEmmdGjSCLdtd3S1i7n8lsexxSv0AbzMWXjJJIa4fadNjNZLYDiW3YRfT
nvZ/s3/ltbo4GYaSu9c/i1BaQcstWEeWxJcxo9DEY+ZPciA77VKOkpaCuawEfSKiAe0jGjMRy6r1
DL5cLQTs2/24TrcaP0dSIesZWpuRh2YeiYR8EpIDL+2E5W6LryiWgUJDlYEFK5z40hbAVp8B7Plq
oxscnG3OSVBXxlOppyIBCC0Xx8QmnxoUttqiUIWzqwoWLxnp8QrkZP/33QhWxx3REBtB1LpNO72h
zaUNQT1uEqlM0NRheBl+RiA0JDQGtPAR+yLcpuTz1Ht8Re1yD88UesnJo91Suki4vUXvJdEghPRB
/wtzSIN2p1p0PdOn9Mb8OJX2PSXTfkhCR3A2Cd4TSRlTqAy2bkE+cJXeztqc0/dFKXFDf0Fra1bN
bZ8PfLNx78QBtjbb47LdFxX9uQMVPSN92DEmcgr1Q0mCFpztfQWf5/PtYvK/DpTBDL9c0k88JunX
21JqeErVQxSaYaIz/DPBzQdY+lY0VXJMSs4sUFKhJgWG0W+2JF6sBlC1W+Q1SxPWFwUaIe+93yfT
VWrqj8kqpUzL8/DLvS/S6o0awKYmVXiShmHyPox85x216CpGHwnIuG+qXu6QyGOig4XML7NkropY
XDYtKfapmRg3TdQ64lhbbhfV8jAVfhvtfqqJPqU0L0vgJ7tIc9JZa4Cg8H4M9mi2RWsbKlwVFNKJ
m6i+k5EL5WVsgXix8mceesuu9mDqDZ2YAis1WDO+18vuxvTsBfUYpDwmXaokrVrXKQEdu44ct8J6
PSotUunxkwYdTZDuBJLHJe6Ww7TzN5gaoTLnoFl7F5ZRAWUagCucTzZkeyKn9wXCJT+0R6NlTNKI
QXHtOVLIqM7b9CfAWt5eI9hVefBCnmFbn5YawDrSK4ZR9ELMY23JtoazsK1xpiB/N3Hcv9BKD7fK
3IE71PIX4jjTgoVLKpcIyp/LHVRyDY2oqf5+dn3B4Rf0NliFZqqyT+eJd96tfF8YIDi03x4TUX/g
ApjOyk7JEDfazCW8Hzy6VpUf9QI53dnOzlDjqnVCh+AIQFTpQShPM3rvan0IEmJSPz9bQZDz9I+L
NImi/CyfqqcUm2xVCCyM6qZd3eex7o9aa21IB92vZRRtxAXpg+2U6cY01ZeCmEVLHB91zCrIdhoQ
1sAtvGOJkW+L2yyf2ggg8B0KJT5PFlyH4LAuqLWvfje21qAJt8UTJH2Ipciu5HqQQ0B8i1kdo+jo
FiBZmb3VLiS77hex56r2QpEiVlqsEfHVEwSAh9T1bbu9z8Z6Du47oOUJlKiIE6XdNmtoTuOu5liG
HyFGe/ZnWl1YdEvX8AKFaLhOqDLxmFF47cP+RGqjArGrTexTHEOYOzVNjq0EHU8LktVUlKCdNCOI
h/New0Db7EjJa8hBSk3/hhtowU5dk1FL49FZaAuqG7FVxIxo594PQdKSYCV9z/oxzOvoz4Bh+mKI
U/4b01bWQl4NogSf8QGfTBmrnpIcXbCHhYv2pf6R8vAfLhLVNX/Hgh3CMZvSDuATqHP7x593AOu6
h7jiBGDaUjOO0chnb5lLwxPS1S33Bt4OIopijflm+/2TV7SF/+E07z3mQLJ814DNCmKF+/84veXF
6sgGi9qN0A6QARe83GsHrHV0Gw81tWeVv2wzsjay8mnz7lGieKZiiWAAd8KMoKvJjfcsImgkaW+P
C/62dlF6l9bRzuL3HUCSgjK4qewOwkoN5ueUmh7CEiAuMzQOIV4rMXPLuL0hfaXPy74+JDkRpTDB
dRheybl4ChfYdmG6xa210ibaqfqQ/wgj4bZCaiPz0eGqy4wCFmxSrYF0+IULjLfUuIcU7tjPCTYF
+eHUALhmrAUrVxY4HXzdlwqdvvdlVLx9TATcYQXl9WriERVKmKqHfl5QFQt1lDuL7D3e8HBQjqhc
ko6y30bcX0unpHMnp3dCCx7duj3doMydAFPWgH5cfjBsL9ds1bZaBQWXSP/FvJ7r+99SdruYZ9JS
l+J1KQdZT0nR560d8Q6gQYrXFyNEfHF8mY/f25GihgBgGh7fOnjY+YggGM0FXLxEu7uOEIgeb0EL
w3C4P1pjA6u56/FCvs63bN7YrQ3gYO3U1kzDSTkOesSK6GQCNNOGcF1I0ziGrhwdFi0e0iGLj/V4
yaUjwHj5Zgx/6gS+AY3B/t13IAYOcOXQT4WVLnlhmczuOMB5NxbW5DgNKuSWurp/Br+46Tx5uJrK
nrH7m0OotoSipIp29nEziEEonq7zq06u9zM1QUQFPwTOFmz6jtkjyZyXZFFDU2xhuF5IdsGVF/H9
9NPdgFWXF5Iw883SE/62AdWFhqQl5lY/5xIOnvcZ+6iG6VXoqN+h3UYixX6DkrXw3OMOGyS9zkSY
iTlLjEaybFDaRLiAHkezFeAD3rlDr4g8+bP1jVFRkhcAHkR7wsnW3/tnfdgEMXZpR+D7LaF6qUYG
uSyCQWzggVHCsxVVuzZkQgAOYA8gAts9SLGWZtR9JKlamm1oGxCdgMRjajNe/qhf5aKBy5PzKVOT
Oscdh6bVjbbmHjU5Cv5rvh0LyNoBYzukugofyf0pymIF6ccppglrHXjFOREiwER6ubxsOnGtqGVT
0iivq5KLIMRy8TpQGF0+axap45mhLJLbwib3P8vb0+/cxkZoM5PEYJzveIIzbOOHZlAy4IS/MFup
3ppWfBXKbDNxX8B6lHmdKi9mbiccOdtoTDDI79bGTNMItli93HpDyAa4E9xzFmyx/xAJcQD31s2y
1gHcQOFklg8EL3LsG5LC1sI5MpWMG712ub7sMcT5lI8+ZYGyzAvJhDlH+1of7wVR2JiBuAiTbsKM
yFhUdO1RW7lN5ZaRyGg6tpdhWgTAEAmWQjajGUYLKkwFs6eo3h746+4PqoZET+BakVjasIPYHHlZ
NXBpO8TE7ArNCAZmy7LxLse34Y9MhXn3Cikunx1qIhiLPg2dGbtCmpFqcu2ySYbVPVXBtx0FVzL+
laoCVt6hM47YRka4ToT4x0k8FRKQSSkX/29txxHecuhqbiv/NguY7MoMRH+K/6CiuxkzpNpafkPs
6dES9r+an6rwIloC7QhS/ukRl2o56ZAyDqeILhBlQgApIfe1Lu/CnWAwzxlzahociNHsGr7vhHw1
u/edeYIutamZIFN2UlDoREjJRYPmEfWfdAPu+puy91AHeUTStSTgGoen+ZmEAcOD+TXe9TgeBQqt
V+Pk72qdIvKi8zS7R+ZECuGscpDaAaQhbvkY+sANzBlxWAYrQ5oL7SO/1aBA+GI53BRM2WCaq+PA
ldB1r9mi9lxw9cTUvYPy/rN4DqbocEgVY2yMHmuks/EDSkxEz4nrytfuD7ujaUqHI4piRUzJ1iaE
uRjVzaBVdjQibWUBoxJtJ726en2bJ91fMAApiz0ENakK0YzUvanM6Sa2LE6qLjKsW2NKW5B+CsIs
8tfS+9AzRE/jnVpTaiM/ytv9gfniapFhT16cz4vT2u5wSgNo7ZJrDsITYJY4gQjdvG0x1z03reSF
Q3C7mraxaWRYOg13lJpmoQSogJpLr/JzzQAFDx7W36Z+RS7DKm5v9c9p0p7GfL3+wTTGyLBYqNMz
hugxJMTld7JU23K3TfZCPr8SyjIMa1Zo0Ip7YqTNe2rx8mSmk7w12Jlk2Sm8m9G9CAkcQV9C1Gtj
yyqZoA0avjyMFsI4fxPl9JApYivchTAyfchEMK+Fb9zvOExvvmd3wMHXM+D11i1W79yILlVNh1z3
eLpwzhoow+SQw1c5mTP/zg/lrz/4gn4ouOs/Q8mma+/9kYHT45aYZoyZLNvTh7kGf5HNfJzYFn5/
aJEM92uo3Jp6TDyd6COLN5+BkvRxCSLFvfVapW37F+R+MDMukF/Qerb46a5z5URrqTFkWV+Pznk+
8SbTMs+aPS8EO4x6PmrMgxLTig6ypajfHEkeAzbdO7rmqbGYUksIkr44bOkO9Y5iaqqLmGtjotR4
kkke59ngeIuX+N9ZiStcr72QSzZ6EKn412t1DA8DYMmwSQa+Pc1f5vVBsNwLypQe2cC4qjVevfa9
gC2p2pivaW92ZSU6I9uCWNKxVWKQq+nWUlkSYaT8lBxTrQHnwGK71AjPnRUjWLzHDvJ6gN+yixJL
2CZR8/vLcMdY1JlI8XOLIG0araNhPFdAsffNFqEpiBc59m5QgA4vJW36cLjQFPGaLvk5DiPcafhB
JoQcfSLcCjvkxLz71dc4kwsMONoFneRcmTac44zxlvmN42SfnZy5nR/jIwF9p3V3lU6zqveBwPrP
jMHN74q/sXoGQpbfrPZRn5zuz8QdF3SrYWMu2jTZt58iGOUl5WWK18QnMXonVhvzdc/ovIOWcpo/
a6MB712w1JLRUnNOIVD27bTQja5u5Mq21TWkDPqupqJoxhXuCx+dBAXTBUEhefUttd/7zidxT4FJ
mOy92nWBoojjbesxry5DlimGtQxLHo95OQcfUzl18w5JhSH8rTBIOr1GNXzTB6TqCRJ1te7h47H4
IZYQfqjrESj3akZuRVKTYaPdIsVEfL0LYQqGaSAwWgSyuQyfz/TSWFZQpXZ1uF3TWaVyYQAsWUJS
LzzUfW4BPLjihz3FPzr8zlD5CQTd5eukMwXt6gmkEewP05TgfAxqEaW4xRURdHlpkI7iHwqy/pzH
vuXDMc040t91hqgPZHl40lrls4JrS6TZe4hL3npyoP1uzzdgwQse0HPb+MXWEBGNXYOGMsefKyjM
+vy9QhszkCm+ddHCkSruMKNADYDmZKwVNjujToVYszrrfMS2DFdjqMTaKyP7DndnwY4o5yJ9Sx9Y
PVot0+qN7//wehPfHH9BT61iaTVg16nNDe5CyR8mB88rPkEvRNEDLlwcCWG2e7OKr4ZIFSDtGiZV
ca/u/D5dLYo6c5RvoiBtuJSmItVi6ZyjTrXmuFoBornthAnH8El3jba5hH/uY/wVUyR6urhhhLxn
aLEkk2rLNrFa09jDKO7bdR8S7SEllMAYg4hIQcuq0q2zdizX5tVSPNp46AgXRK+Y14/1AwmRpz8t
6AbLM0+Wn/ZnGag58pRWwJoVn/xhcIbh+ZCd55SIsx6mWmxs4UJDWVNpMcPzzD8wzn2ZkMvwFsBK
jgk2H2XkByiYynC1zWNwxAKTczJMhOx062mmbcJ5u5vqfxSKCslNYQIgcpby/QPsGD5poyMgG6Nl
UMo8O0gKvAwLd2/wwWpvO372r3r8QeUrTI4XvMHVm/tzcti/AT3aw8b8bX3hkbOIHOS3uWmg8zvP
g0aiuWmWhv32VvCig/I00zbL2nvAjtov3jdjLlZrl4osXZVX4Lb8d1E8w8ufvAFYIwGplcP8/FhQ
gpNLu60zJzmOLgXRymkfhPOPqqQ+qj1YZOEtPG/FAkbZP9VNyaEgx0V1O05uk4oUx/gN4NAhWZOP
pt0p9i8mF2JoqYFtqvcLEabxcbyVNLf1o7AaWkDpFRNEsnvzRTDXv7BLGdFOrNPdUb0U8OR1+j2Y
oKPDbsKKQ85NnmprSGg8KpHgJDGU0NJMOxHAiQKEL6UljRuRgIj+m9H9GJSNqf/Vp9tRZF1Avi3l
o9VOz1DfAcK2QIqlHlFrKqnih8rvujEaj71EypANLX+FDdS/atl1fm6hKkcPQGsRZpJ0/zzjb6ks
0qBtd+i3viQvzbMDFniq5GRWkci/0sBlyikYZXuNkbm+R7oFAr72gF06NNyX+gOPCeDDRegWN3In
tgXEU/79huIUhFmkiEIS8goGg5oEcfBk2K8lhW/xD/ke615Erxdqk3sqFd4FiWSjral0mipjuWUE
iVULxma8jWxdxDsyAEkK3Y1PhEf/uoV4Nve0VruRLLf+wK3eotkG62mgp0SNatgNVhD7RtlQpEQt
iFSKX+8tu74DFe31H8eA5LetLYrH5PT+mdbmI6dSu6RkWwzvbnCX2AJB9lL0clZ43AORVl3S6aXC
Os1wo2Avz8qTM4Lr7yU4szeZNeRQWmyeMrpyAuQwEx3bZHGCCuSfkohInNDjHuIS1pZh1/vC5Qmm
UlrA7PvAX+oBAd0uzdYkV/jX9ZSEMilV6gS9OjJdDlO/rBYc4j132r2m46PUFoz8x6uhMcRo/67F
/sfATkEjTqLajuIPZlcrTI+oasQUzdhiXKfwJOHe9GHVKtaWiEYQ2Fm46JNq4031nfglAcdRdjKP
52msKqRwqzj92hMqoSGr2xAx+34M97h6OHDBMHVC2K02owEQN3EK2W5QcK/qG9PI3IohkEjecyQx
U6qSNMtyFFxO89HTHoUpxw6ma6GbSgzNjqR7wSqehtt8sPi6b9kCcSrEEj6yCOfuEcKUv+FYw6je
o46P7PkAKCotCBpu8okECT3LYXHq59PYjrgPkeguUMT+pszzPI6kVf9A7kTwsCiJGjvXPAjOT+lf
0M0BBogIVdop3lL9QLmLFGcTHfiHPUrDeDkmt9j7Dz1evzd5SUADAxIsiNtWRB4Snmz2yqbRIOBK
ayzVM07Xg5nivoSzqGLl3YFqKNGgs0S5bV9UmoGbr5qo0pQAO8gx/TH3sbLhHXOsJbWS8zBA8LP5
TumDP++3iV7/O472PTkZ8ybO7pL0r8Xx8saVRTmL6731PCRyx01gO8+DIO/u8An0mU5CrMmOLyWW
iJ66PSYzCcbIiHjTPGevGFmvNPCBtHxEIHV9hE96DJ/uBxte8kKLzeuXtbTXT3Rh/n6s/pZN4pxy
bVfPd+kZy9mdXOIELJPMvWMYZKJkluYdW3A/b34PnBJPxVKPQhvVlW9j/hwnU3xNNjwyLi8+h1eQ
YK4l4rFagO4r26HzxEhU6IXgYK70H2GJ9tz+Tt83cJU4qEI2k0xPawCGn4HRX/RdfWaDO0TgJ+9e
VVUcaOzLMzUbmrc5uFKrGqWnHgDjIj7+Jz0z+ZPJkE6/OxAF9Vj2XEPTIfw4t4xzIq8ASdk+1wtJ
1+tdwzJE0PoFAyV+oL/+HV0Nq4oBxKnxNUtW8VWU++d8T6wgUaBOJnAh3vPRqfjrhYpfp45Is3Zh
Hunc36dR6K6IfpzpdlUbThDuRC9F3da4sKTI2c2iwLuJhR93lJjguw6E8o0RucW9GwCzesA/zE1d
QVFYsgE9anPZbegYrxaipE02WQMj+hBzL8uQTGhnmCEyMMIrIGa3QWyZgT43XGqe0xb7FH6HD8SF
g2hfhVIBf9Bb5hI2M3oBKMa6AgGSewX7+EAdorirPmhMo1244QsptVFBtCWTiZhDQ/dhe4m7zBZC
zPhK1UqBgSHQkz4cDixf5VbYcmuOTmEYynVgKa/8laBfPKG0dRDeXF0Ub1iX4/N+KtgUokk0+Ywp
prNef4a59ybjZugxe734v59bW3PSk7iNc0X+aiV2xIifzGiF7A5tvFN5BqsGkEWZyCrUjDl6PAXh
8Qu4yh2SQ9zyPWDzpMzfFvXVyDc9tcGG8PYE8QUhhiTXOVeV/2Fw3VcalfkcHWHLG8bFPPu8ePY5
ybUgdNVa+NJixORh94jEzCmPER10QDgXOHPXX6O9Ajqy134yx0UO+kueDe2Ilrbk8e1Fr38nQcxx
81gLK/+BjmYWRBzyJpM6/gBt+3zB2kjHijs2ph0O0vAgGe1fEKhjKWdKk9q6x1AzOwwGMg4CfvQt
lrrnW+RyVYIDS6mM7160qX+dnpe2GkVsg9yKSH+GI6bZ0Riegpl4hPNt6y/+wDYME7wP6Z2u1kE6
RmA+Gwcj6TtwTcRYllq0X9by+BkDUyqP2ICHJSrgD7RUd9meD9Ct9S/ySjNapuq/VQXXMSBaJeMn
AkWWt8Zs7Wgo7rVTCZMf+B2TvLu0MtrUqBsH0bgAWPF1pj2cK9c1iENdk/z1Tn40w6j4AN7w6KBU
XwqVg26jxXBBkUW7KE0ClPf8vOgAup+pbTXl4JxhGCBNMMUEKGvg+j0q9FKHaZOMZiPrVPUGLcN7
Icjd8CFUvWp8imLBui/wWr3JL/V2SkKmf8h52oCpfWpUOQKdNyscbxx3sLY6EKzi2SH2KIY41jSJ
ARM7M4kVUJQ/Kdb3PXXHKmI4TmKGJF5G0NYUcj1MNyNfSW8H+EICP/1aPuamlBnn8wTmRDY6jPyE
zu4N5JRP6UF4v9JGPNXlv0RdrBqNoUJIwu1L1Giwdtt/8OULxLlFXCU2g2AZoBBu+Y7qYswjI+SS
uIDh7v+N4cZ8/6bu9An2s9TozDt6HKsc3Bb4Oc6g0w6jvghRGbXunA2zP0mCU8YEWNfMnpVSi/aH
ab1/Du2UDJ0h+Utpj7/1sluAD1ripN392p/6WT4KP8B/qukxU2G411bILuFqP4HRJ8PwZYbi7A8l
LLoXCjRHm5rI7TjHjBbJH3Nt7e4Aqy7BuC01EzYXzCrIJQQd5KLZ6yZ6oIzXi5rPLlmfzbnpAh/v
Cqr/A7mNi+tf2dbTPfMU/I8L2ZE5gG+DRRjiu3P6B8h/UaoDx59REe0iGCniUhvlE5hCkEiPyJAp
JOo0/uZX22W/cYoayBk66YccwPycDjtLhQV/rAXFE3097V/DbGPvglUbDbnVK5X29BLLXqTTuqin
kkUxABZBnwgyZeP6faPB5N/ciryBYPXjnX6iNi2iHeTQ2A0UXt6yi53iKrsYWnMSFX6LhKuJQSBU
3Q3R/x7yaeXrB/TJjNVhpqs++fxYl3I+1GW/9SjPU99FnqgDSVzLdJCIMQWYNz0Y11kWgeROoSB4
d4gicsb4/atJITUYPkiSmraEXj9CGuJIAG7UAqxYYTTI1EwGVaEd1Aji1TuhYiWh4Zd3WBrThlPV
ba5rc5J3lRJw+dz6InLRl6F6WqzXdN4FtJPzHmcsRPC1gJ1c9CHGXnXjibtiykR2rfDJWJf8Pcco
+MUxlifCecbP5yQbmE8hiaE8/Mc0ypec6Q9IRMGS+o0uoFfc1TqIurCOOFFhnr8s790oR1qavUH4
3HezvssEiAxXrFgKW7ZIsIT02Uc1rVObtfIOlIz0l2on6j42HxTgj5UDnP6OuLQ9h69xaGfqUQJ4
LQMLdFkZOGLe+usBW1FlZvnKJ6o1AMoecAwOwlkuZNfTTPExqlHPb50DEjOAEBaPQSI/cppkpLg1
D++YxuGBC01gzJ8bazcUQ8b8aBZwh8Mj3aL7ZP9GJznyOXXoBoN5TMYvmofVJifzKtMSTecJZVi6
Z3Gj2VxGapyrxecjV5CM0mRV8HAd3l9Lm9Kv0jI+dfCD5xBqObUFG+8+hML73iGW0yQCwez1maMS
as/BiLGboYcJ/Oay/OyLxKRcuRtMS4NWCPQxOCO028S4KHVbtW+ZxqoWudL7/HJcfBAfHngd9RbT
skSLeR+CsO+KCwkUwZDsu+S1kb2DvPlc32f6flzw8tA10uOKBmTQPasstyO/GFMqC9UNEJL83Amn
hD0Q9gI2nJiat/1Lh1GbfzUvdknpw8fTicKCM3pgKucSu2Y4pOH/xtE0qg1wGTbQPa/1agxFnYwa
krmRSOuDEC1uexLg2wciT1L6MF8FirB3yWkVPrwSS2jxF9weVCUsfqLISpOH6UPmcWzWdCDd+mw4
wL59QtLItN5k3I99PwuooT2Kz+8zYsEXrAS2HTWlHhLyffAZKVkanHk6kOqxaET9GVGxaVf+dbBn
ZREwLwdXHmdTxzEcahHfgRBfJUF+r3bCuZpHSoPEab1Gm59S1TO3MLe8dWLS4YRi0MuGefn4wd8W
cpHWrw/cDrcqK4tkNPnrvC/GoiMqgybcZndi9j3650Jw0oLHlMD1choCX6yzbObEMGN890CvvKHg
+wk4M9WwXAre3/PMpSGDs2ddZI/f+by1M+ZD1PdE6WadiATmUYbfevTUS4gxsiW9HuAKzF3fQMRb
O9a1n2Y6QmdstgcO4NjCIP4QUzw1QX/HXay9tr8N+JaVXM1Sx+0asySrYl8VngkdbCUN5s/QNuS3
DFrvJOJuVw48c+0AkkzD1AGrOWzJksrgMgOjuDLu84Indpx1s0+WytRH74Tpj6L0nab9MQGtwJF2
0eiYarECkXgTypl3tYyrV6yNDmaEA5KYrPy/MuTakGOcJO8af7BY/hvAU8Q67j5pH1wsfmg6Ka9K
wCCUxNb4rayTnUyaCVxUqSUnzQMGvOQtxyV1kN/TvC/O1XOLar/d1tvgKSCddVOvzpmUalqFALAC
q6gi+GF13sTGrVYXPbg+ajRSwcIUQARIOR8gTTgFZx1HceoeRKRyVIgJNddOxEH28l3MfZJaOaH6
hLFam9Sh6mQ+lV+pc9Z1saADUxHf2FLvlnTICDPyvY/DIFEwZc+0lQ/cWRMf0bbW7YMT+i5swhGm
w9ypIDpegzi6w6SxW2gBgQivgLN6fvDnxuric4P+XsbdHXGwd3wSRUslvgb9cTjwtFt1EptBvf+W
HNFuFCJaZkPUzGaAbiNs/O/RueaNaKfn+a24PovYs5MaZ4dR05FhPhDVAGsIAyg3oiyYVQE5OAY9
/6L509qBjNTAjuUUiPLWMZhRsOZF+tYBjvshp99KasJC3N8HqZQ09vRjVFhMGV2GcSt1Ho4POhnZ
z+EugGp4gYNfrw86rr7pkv5EjwZIwzVbr6sSfslSc9WprQwg6MKdAaNLsO/ZYBhx3NxoCtXbBVuk
ChiwFB4l43ys5ifS6AR877t7UdYkdpe18B1GvLyYVu3U27M1PFrsh7Fk/0fE6Fxwq/kbcQyOhYyk
7Ew4Ej02gLANBJyw3uYzBtPYK8WEHeZtNk+8tBNzBiIRjDDf1Jo/TuSOdbGEuBJ2II3aI/yUQJ5k
YU3vrJkh+I8xsOY56tKtuud1ulvn+uF2/udDotXvH8zT7wRiB1qJ0RM5AhX+pTqXa5TOKthJCWyk
5fpcNHb5JlZclO9g2vDbbA432kdA9Lt7TBhNH6gm5JARyVgBmzAgU46QIjkJCzyaoabUqOaE3D0S
A89Z+8MA4qMmY/gMhtzlm0vqYSiNXFbdNqOXGLldsIlP8mlXLL1Gs78eIObM46M0BeY5DyPz/aMn
VxBMGSKUiCopv63abR+/fkl8GrVWkPlxxS+/SCFM5n634yKo82WqavK0QhbKznjyDs3B+m/9VP0i
MzWMwy/dsWpXhf/C3UecuAeqZWGTaKX9eMKJoWlGEdpWkS8/R8OwOPVRe2mGqUN4M3zsrIg/V/nn
Juk+z5wgSt+PZoSStYib22eWOMKmzSvm8CDypjPMO0bT4HYx+XlhThzfOmG69Xy/Bb+/Bmycldv/
M2GEnVF71+/cD7+Ugqx2jh7FY85r429wDjiwc2Pw4tNiXhsyOzA6WdWxp2IZTxp9cPQJ6MOsCCqD
uyGd/QwFj0C28o6zyDdM5qx9E2aBTEOhXWWpziuMgodyk3gC28byJ8dwd5mlG652KioiYXVr1PBW
2JO6+SMvcnQfe7oAsLXLHZFJwbkz7tyZf79xu6wylAr8/nEtzJbpZS4Zj8skfr8MAtQ2C5LIsBR5
CZLvljD4d6PFa7ST79AgcEx1FVakgokQs1tTDCa9EV2ii1ML429nWkI2shPb+gU+KTHrOeCGijcf
0vuaHDxhLjUYdg3wzR5WTh6q/ftZcrCgFZxbPCGAvNCF56WFImMW6PssBQ9eAng5gHQpYjU2+YUd
4OeeioFhoyCediKC4q/5UEWDDCK4pmXOsFhOvL/YXfvexVpSrThaRgYaQBUQPtZWymSwYdWg9Vh5
xI794SoTRuNxp5BP1FE10wS+D8dysqoEJr1QrY8KuSHmjyW0ZdN+LKQI6sybA6/yniju2v5TYtqa
Cgw1NzhW7xrg8Fy6mOGsfTK7oG68AroJHwmxmj49IJoLoSwg5NiXGCXGnC6xFd76sBJu791edHOU
ESyW3cWPdVDIILUe2ptvx5solNaPDpahkXMuk1ayQ6zk9OwiDZh8OtpLAjabUmbiDItl3T4hPOD0
fOOpBskK76aJPPwg/XaJftZsyOwFJVlCozCxRj3lxEj+z0kZI7Ay/vANbF/61KiLOulLHGTjH3C0
tlz9zxUhKgcWCJEjVt7lcqVsCB6lGHMd65KaELPuGM1C02tFxQmSTqZ3dlc/cwl78XkzfdwNifiN
O/5JQgcvz0XFYb6t4nProFFyrY1jV6VOlDFZTh1IRdHfhRXrfLYmatCvkF2lJJkMGhaT7IX8pzLO
JXjrYjuSEFrIZeBo6SRvBsj27futOoR/2f7Qqne4/5oMKIYb1aca9zHTidhrNAA0YJQu9M3lhNEO
0eh4Hzt+PSfBt0VgrHJl7p3MHnCgZj6vjy7fkSYhshJ+iNCLtDdDXRo6o7hJL2QfJkVV/AjKE6LJ
BF1HQSnX0tuSdmJF519/tFFhU0mPGvgEQ6FMRUZZWsFHhusR+I1MJAlQPgsCP1VYj2lG2juMeVad
UBdSLf+mzq6Kdw70109w1g6srWISTnQJazymRojSZJs7OTvcy4p0oRUji3Bp4E38fGryaqqO+CUv
8M6v5uYpMPbtfwKBUMa0m/c1GiiHNqxuHp9bpYemhJhfXRImwQIQIW1ZCu16k4joUgwyJoF00Y8P
ZCEoQ76t9NBfsHVQn/GH9Oh93pUzGUpmcbmxiWNWPoLmGIHn+dSZYpID8CjzVCT34OaqgLGpkW2n
mbsB5I2uWQvw5sMBwW1XMJHtg/nEx3Zwu9bg5lPXRL0PyF7BOOZbOoX8W2mROE1vb1BsYj/OZZSg
qlv8fF0wNazD5zKDuHAn5KPx0G5psXCjWCj2zwFH6d4tvUvb5A63aE98rT6r6fN9flKQzk62Ovjl
MB0Y/6sKX4+ZF7YRjaB5DmWtyGwhHrRuCUK/ke7ZwV2o8K0Bn3Zb+fHbCOTplDfl59kwxMarrSDv
IQTvF8tbRVN4ZctRqMEzdpdLsi4N971h1RasmebL/ZsniQ020+Hy7FqtI6/1B6Ui1KnrUoP0dtHT
msosHjnLH4tll5xJkogwL5s7wbKBPH2rM5Mso33m+Cu8FienXWkBpl33p48uDhDyrw8bkZTlvObo
ydL8EpHTLJREqUb8qEyChmqrWRK1CdNFE1VGNTVwMCmAZ6f6kASTYlE1SxkvSHaxCM2ZQ0TXHcpU
cSgacI7GM80630hPIUlwuoScqpcjeNmr7IHUXPVHZcvc/jsWCFhFSQ5lll88MHAUFScIuIbpvjrW
DMTlW1LqUpKsf2Tbe3/v3kk09JQLa4uQ15SGTcXAsAyzP0oxJBd9qgHelHbqPbxkTTioOUKvFhDy
9e0mjEPXt9C8jaNsSA4zaZyRxn87NhPqzEz6N1GhJGPaeN9D6iW0wuoUGLz2Q0To44VdKflhuIiA
849MreXPx5YEVWYOIrPYAwTQiW01OUlBc86bU8V+IvAQmI4UJJMRRDFgMYjHgDBo7rA40qLCZc2S
7oHsLGOKpo8tVzitqBwaiXHxS+lfvd4VX7JsfQLm0jqlS2OC6UH+T3aioq/ZpSGDAMpyMR+3Q35B
vgYCXwRVNKmN2J5Hm8nBjNN6DQj5FXKwHFjUWjCezx42dXLWaytm5svXw5qEpAcGrEnHQSxpvoUl
9RG0lwOlTbC/sFBBzLZ6VZgBWR8sO/cksaZw/p1g2/Kg2nf8vSmdYR4J2MzkelssjYDW8+WZg6wK
oIWix5OoicT65fmAIHLEBK6fsgxQ8+A6Y8eK5BAIe/9mDnUjCe+tlzfh1XllgEl/r8d+3FFmJZrW
1TyULH60DzyQV1owWwYVA2JfOnCJ5na6XlBUDdW+qa+xJXLoYdleq9LBC7m4ANaehRgrkERUij0h
w7ghKPQXzNGQ/jyuoPH7ToS2AivmHFHcVqEnz9r6nBYKYxMn8bXO8z/JS8ezKl5/pFlTfQs8xuWF
GUGjLFuJlp9TfhLzomnOOODCUu8QjgrbUY04wyz7i/0yN7plB/CbDg/PjHqtLIMYaQvUNVraSh2C
9+7RNa76u1pO2kHZLymboDXWegsB9510tcZM3IzjFWMn1FhaTrqQRRwcuDDRjieovN1H9May7TVG
KFbLT3UnQloFeGp7KZolGJRj0d9PgG6tsSivQ8AMNUF0vfge7/eTtbMtAIsMvNw5nnURpKY/r0aD
vRZLm18rpOUJTyXPzdPBzkX54Lz1/2i60BttQ3wAl+Txhgw/iMU911Xmy5oxIu0Et8enDyPAx6ul
mQLKkTLpVWyqWYhzhwCDrOflOaC/l1JP+Flv37JeD1DFFk7dY8Seo6JPgLEAb0PutXwgH7VHfxbd
AD0H2umu8Uzd0IMkNJXyYjNxBSPQvgEx5bRMqWZjaM0SM4aYw5rzD9WiOoua+GXav4wN/1aK1/ot
4No2bI8Vm2yGMchnOAFhOkWZEBaS8f/Jazot3X9BddFlgjHim+rFh8zmyEQRayJA+F8kxeKLrS42
cW2aTYl8ExISgWLrPZps+plFN7aWcox7DMXaIrUc2SeMABjBUMOJ0lSE75IOzF6prc1hGOoHmtx2
bCP/rGfafyht5dvrNX1RGWTKbVqvcwBL5iJnImnFgaPO0gLEFm6/hGTTpTHZKEGEkcgJO1E9wNNg
+G+jFRby9GLD63Gnc/GMI9TmyQ4rsN4gzhuc4k/LXr5ln01akoOP/g3jplPp0t6vbLc7AXNk6rf+
OFnwCMB8PsZrRGk2tPKXlpmmCi6sAKJ4nbJ9JGeaDsQxB78fhhKkNVCcLReWh4PFEkm0qPa0qjIH
qBQROC7QHrJBPnJYDu2jKrIyckuC1GonZGWVNGz9GbLP6XUg2368wmXtWmKWJvkM1nT9VGVwrPP1
D2bFmLm3UqlrrITaGpNj1AEkGKa1MxaRAoHAj8T0/EdXjNP30Ul/K3dI3H10c4ZJA5IThTRfyUDM
ZcwWxu8zsNSkVOLvqaEYw9BqvwT9H319B1bfx3ncseKX4Q2kQRMblXF7pghceCPK4X7jjJnd2Q/k
V/pA4m7oZfXcC0TvLolp01QrEozZ3vG+XhMwZw9CqU157AOEA3IoEaO8/6v4gy0+gciLM5k4ZzNP
jkHqe2alyeqNYNjdovDca+fe1b+EXUP/uNaTX8TBGEvmsD4NBmUducFYKAXIQvuvG+Lm98aJbQPv
uwtbP1mjiG8d5/7O9MjDUHZEPUPqhGOX24jONBfpTHQX8wMcmUrJHX9Z5uDfjQsBZdM9x9u3QxL6
st6zBhsJLUvIBiqm+YLw0bCnSU4xV8/CVijRSpUGNXL+OpOz9J3fSDXAqXzqINFnICJsUG0wuDmh
nfM6kc8d0kTKKsvwZPItckvh+rNJRawCxDgdSRRMkl0t8ZoA0f+adXGEEYPTT9i2rfwa9efXhQuc
OTPOpqyuDkC0tRwOCFnq3bbsbRhjKT5qRVuc6xgzAlhA+UBbtVo/cZOIPHL0cNprzL9CzqXPiNrG
uM6MzG9qbZ2skaT0dp7ulnMAKy2ymz9mecAHTAw9DTbE8tkSBdQWpMakhOJVrc0NBZj6C2e/Clk9
mMmjU2q35PeYTZbYjsaikBFBRqmC57e5xt2CaYjPqQuOAjyTAlaxgDUyeUfp5LowIyQPigXpOG6R
qa8hsLD+wa0BwWyGhFAwqcLo0YTwjpLk1uSxPDlznyfVSrYaPMZeZ3ArnczQJWzr7gQZxQq0lIEs
GNUq9TiZW/+5GxIFGw152dA9LIMi20DH2Kb86fwB/dbfgMpyWN2aIp7uAyQ8LibuT//p6eVXP1wy
ARlI+so1uvhj2IGBTcbooABqpP5KhUdjP+1BraUaFvqbrgU/RMwJyqhS+rY4I2C21VNJ3h/9iqT6
2AXZEXxA1U4lx3MRslnztUMExpWBCuk4NkAUsVIv52LohfiTtHSiwgmDSbk9ZmGXgidMXrKVwstN
W+Do32h5P4E2IJtC6CA1RJlNj2fgXFp/83b6ZcwzIX5wnVLOHLSamH7LhcNJlBmtECGYs0t6meHi
mMuPzWaZ0sUizsQ+9e73aTwRKamZ3bQwaLynLwPzMjegZwGitM81tIHHQYZT9KKhZ3vW10WB3xqW
KE3nXOVnegtEpqng3xxe2/meTh2KhzYKoafJPWqFObgo/JlYy5z/dex+7Qwcd7t35wWKXkVoqZAf
K6AJHrlfDUgLqvM/Bza0ye6cW6TCO/e5fRJR90BZi49YRNK1XxMNUHcZT8Gr1Wdrdh4b2QvP2k5q
zG/LAzG6iuQN6N2tD+AS0YCvOSj1NyBFcQi60m2bp5UrDWheXlEPAdbfDB5BvR8VZkmlPW97w2yG
9Cd9UsSeCCEj4Vpk9lcDOMfvoOvtQmQJTpio7A6QDM7nKuIpJBqUXJwcbXbHfDCleoAEfeGCFN1x
rbn68YagSmjIPDeVNztpjDnJrarY7opcYL5wwauUlfK3o0nbwSWri+S2nQPtHs5Cgj3QlcBYDgB7
I/syPU6bArgcsydNDeidkzqi58QurnXZUbyYYXBmSe7bzREmnLBidS+VQruWDccjUz/aF88VOC/+
EP2CfgFUAPEfpF0JfhhZxG1NvHeq3rtjvMKWgcKaa95ERXa5AJM87FzO6E+I8/D9Ic1G9BcbwTaz
xDLY0h+XkKlwtHFndDpxxvx0327Y6DGaYEno+iAsQ9pEOqv8cTkyFdEqs+yHeONEYF6W6fYDxgsp
9h90BxVqnnftQzyOnKBJvMwe8fZIdlfC9dgoYTsNBKKEfxQceQWZBNLHNbkOIKH4IJvKKEcGIHXp
Xyife8CbYGMvDlHMWz+XyZaJ+hVVA52Zr+BsVl7+5GS1dCXW4mnHlS00+pSC6hQa9PZNm6yIx8ZL
wbZ6RBszKownpGGawGB+uBzTHhpET/B//l2/rkyDMivXBjJ8ClwNSCNsjCmnN66umTRspDfIpa70
1JfBku1krYJFNjBdauZGW2HSHgAOezCbovKhQxhwX1cV4NNwGSzQ0vslGZP7X4/SwUlX/04+tpEc
1AXs8+aONVcvyPGtThDIwVoCvei0DACfh+JK7TYhUNAp4mHCkrmkCPLbEuSo+WAfO6dc9x1ObpQZ
IfDyXJL5kgvcGTqpiYETLE8+KtNQgaG37m9Dacc5FWK2WupuhH3hpLUjVl3oZPssC2W/AfsFQSbK
gf8NvyekScStHj8WRE372ndahSCIBnKtPuCSM2ouEf8m5ybTyOJoB03ZtGYo80KQj1OhowIcsod1
cT6Q/iDv8xm9qfP8kp6k4yHUZ+ZanPjbdjH6CnHFvmoHP561L0q2RpIe25dpZG1Dk+RbWEmpngIR
omIlEp2OjoAZQSxsqbHifNgdn6ZOZYb16WIQGdXBtT+ZuUJb7cWpVfT31AUOzVgVRS7BqeD1a1g5
IMdR/b2xUF+XVqUXqwIKjQw+A4TXwZsPyyp36E5B4nn/0hhPpvlpXbnJEIeC2K+khhyAdrwIpKXp
yHO3qpxVtlLy08Bq57tCKKPPJ2CwSNvT6gJPqbcikec6n98GOK1TEHn/DnOkv06hos79kWt1tW5y
VJUGc05eN3RNGRKa3VpMH4WBH/+C3qIa4nu1EngXiGojQRoDeNkkFGJVuU47Q+0AoBEP590dsFdC
eKV1APvJkGGh2cMtVYS4KVTYw7+5xuCWZa2CrSnYLUaiqJrrQjxoAdjs9xt/2hTq8bpvhIhYu8/B
jrnlpLRFLXW2nrnuslIIv1L7e+KXIOhPtYeumfx0ezN6d+T/Y6+uWrg6s34jz7oMCj8I128lTaB7
82EkKh7tk/n8mi9ID78F/rIIo+/ZrleInoWB8w3TYWX5vIzXbv6hnfnI9BqR9FEDWUX9xPFUSXiY
qHHC9AYtX+3AywtONxRtg2fE+JaJXml1qDo/3K6Tb4pJnd4NmcFFo9zL+UyFcAkqMPPz2zI2jijM
evPJV3hN14i3gLNOFjdzdJIA5AwCa45xMGBk2j9Cgfbr/9/flkTIcGl/1ww8Bf13WWMbYaJP42tT
QPgl0KCbiDMrGCblN/1Rjzj0Tcmk5ReUqvkVjrjZsocJmvgAve6AJUVmkipzh4HBDezljSPF8YLe
G1kVMlvhbb31+7z5q8jj3dznnbo2F2DoxIN/9P/1vEyEFTSiJ+qhjyWcLE2NsGUICQYyHILi4S5j
lczVOTfgGh+rovrE9aepNc9f6Eb3RTkGcyMSEGwxXTME5j7UuVPpa3TQ9wjaXroZudBuVVedQvhv
UM+DNvRgh+YXOIqf/rnNa/ApbpY0SzkDny6BNGTF1JYuDN7APb3m69tteSEM2LyyqaWgWxKpblmj
ZT3YUgoQ08alVXM1UbdiKsURbHdpsoYS2fw1Ci6GlRGAmynCQZpo/sb2LjGibnlOBQRfA7Co5G5t
PhBtpplfnRvsfV/TLHnZGNSc8yXtoHksNo3cUEhd5It/WRobJkp0KeOc55H5Lsy5gbMAzxbxH1Yp
uI+yout5hLwvzQvlrrYumagEO5lpnO77BkNt2CP18Rb4dr8YM/1bkPIRYUbXeXVF7HxkH9VkVDZx
e9lvsNHjBILjq0h1fGAqwPGedc3o0h4/HpSD7vlHzCTQm6K1wkiiuEvDrJzh6fz0XFuVefomNST3
twlFT+7ihTLcZYQDefxd9OPhn3s9UHV1IQd+/QtZOK3BvTnGNepk11fLJJ+YAFFFT2hptEsIvNMj
zqa5tkDTktQoDUDSk6OxXnE7z7pYZUW/CZljpTL3WFSSVqNb5UusdvZ7mXYXilj3D30Y7zQiHn4l
Fc7cKXJtMTVf37UDJTwmEr2Uut2Ri+gEQytfqB3sy5/vrWsoCa3J9+KUL1KNAEbfBmArhFLDZyDL
cZr6LOykwB0LW3D0a8hY5/OzIwvRnwiZJk77SxhTURZ9qAqxHNVSOnqAORtEmVT6Op/bOxeD0fGj
n1YXlcRhR8/aPOgfncWPhJvZsmyrm7sdvWBKu+OuOzZ9ocCIZuIZ7DnIMOcTD5ve3M4GAZXg/0R2
f4+KSD79f8qhxx7H0CjxTqw3GLuTQaE7N/gJ9mvAS6jdjMvSLKywqRFZNQYt9BSl+lFrIT2OfaDb
7aZOHjqeVtAn0MCbwJN0JMtb1EAPOjEEHgqRtHjHav8S9uQqeqDa8aGRki4MEIea7TdRbdPYiWBM
pNDUcB13Kc+zBCyEP4MmtYSZdcwj/ySnJ7JeFE0ZGUGCBXVEg34Oa4SGDBzH1oRr1/RXv2OEi/vi
kRTy7cUei3VSX6m+Fbus52AbamktkA/iiRWDgVEvO+oe6Adzz5Fz7Lppeqckun42883aQmIg5sna
xy+Vh85X1qjjMpGjLfm+OAtWCSXhTjL7Cz1qAgCbA/3XO6AQFnaVsZLw1gzMoP3DIofT+Ii3ggiX
EHldrRTv07d93B5R6MS0q/dJTmir0Ii1QQqp5h+T6eDHV3M4jlQHjw524W9yqdJPAHSKDI+Mc5Pv
BlArzhFdcRtnQtUKBppmL4cGP+83PhmNDBmX+Fpr2879w71il2DIFZlk4iO8XmBLbng0zm3XtkIG
EniY2HPZNhUHFHtNDSeqwvxvP3PDLCaNM7HWHrVHQC8NNC9hoA/n5MxiwDHlFLNZkU54fbLTN9A4
+HLvJBSYTSRg5jHFKQSSHTUwtmEjSRqXrhX5iUbxSYIosrx9FcgDfmr8KzXH9s5qKVIQnLLNXJkN
9qUCKUomZ7+GWEkVEQRy5f4jNApGlDtIdOZIkpno9H01SZ+bHT+5qdgobO26ZYHrH8c8jaCOfqL4
W45Eo5cQbtBy5JVHIzbLlFsaaWZcAM//EqKOLdtUIMJhbc3N7e44mimlqmNZJZ5OcJp4Qf23ucv1
KrO5ofAkTjKv9HELz2cE2cC1nAXgwY3HkKiHZNZZytdLxkPgv1IYrrWIgSD16llE15m1nC6hP7oR
1cF1yG6q9f9D/B/SxmI6Noez/AUqqs2MPLesnxSKfwx7tCPHwCuuR/lvAEbbzuPafNLy8E7UnlbJ
/3IXgMrRdN2P8brTxcNJOk3QWXmYfrqD2uOUHoh2gxLaKCLIwGUX14aBjmr5EBDIkNiG0tackWd0
X1lzsnJ7SWmZ+3JdsgqbU8VcCWBIMBN8Li8l01Ffd0WACnIsn+7jWzgrmrUuV/eD5WeAg2Y1mrm9
cwJolmgvDegGGkRbt67AJaUNTwfYrgbOh5aIiY88LV0F01XsGumV0c/i4FfMrcP08C8M7euxBwgS
sM4rRQ1llj6hsFrGfJD+moNppF5Q8Xk/X/ZSdHEOsYqK7vNRDk6QSD1yDL40PtGDMdJe6b03B+je
M7vFGvKiolSEE+S25c37QDEyib6Gp+/3ytf5szdhKppjKvDIiwUma+Ijf1DVAVZ8vjSyUnL9DsKr
dxBjsBEyd4TniRFD2ELRY+b9zBkwQD39ZcTyXoYqHC3IyVTPRomO9GbRs9X2e3nHu8SIn9cJpkfi
HxAwPUUSYXA4liUec7JQjjs7qYNzp8QMCkTrizh/Vc4wGgR058jQDUqPdYFVU5epp4POATUVE3xb
Xibnh+gOQm/Fw+5C6FTZe4/BkZNShwpTF1az790+MrkPBt4a0Ew6gU0hwixMLyxwbWIzAdAbjKM3
RbaUcj/SGV/q457h+38HIK9vowYWxgybQZ09RN4L9L1InWZPi9lL4bkQFkouiFaAPVlUEfwVhv02
3Kz4xq5aHK8wNHwDbUp9XWXBlffZSY6MinyOrg/gSZZqSsbEcZR29LPRTtai7MFh8W5i5kHuKWWi
O94wrpusN5e09H7sDizbow0AocTThQA0frhoP4S8JhVYcFpvDVwvgWyFxYx8JMfY7ZscwrJ22iPh
v5poW2UoQNyw5+S3E6k2a0Ynzypw9CyvB2bmN7PxUn3DIEI4a44hWWBg9zW0seNqKUYkSxpgVorp
Mntmr8mY3p9Jcic7NL7w/bWTH5oDoIJpACz+/UAW6vBDdl3AjKRxdnYEAGVNdZLOW8ugjJLOutFB
FKlgs29NDhe8VMDVYCLsNR54OK3J0qH2pnGwX8egV3WteE8GBOM9/llS1vVV1qHJpHDtx9DWjGWY
u7qEjpFJC1lY42so0kZ9yG2VxTtZyOEPfuVIItd2A9gIsFzDiNCCJ5UcEJ8Lnm0DxdoAAHygzx0l
kVJdFP2zCb5mFj1zUUrt1NSNSumWJX4VbVlaJXlo2GMIVXoplhtqqUpXbOnVqHfQrPhQmjpO+lPW
T9o4QA3nGBcke8J0E0229wCAc1N4EWMEhSPWMZbQW7bPwKQZ1X/kNMjpetiTiC90ezAwDF+ppznm
vRWYgGFjQ9Aed2rSY0qyzgzSPvSiY98yAh2OHi6QdYa3xMD7ltzI8IYJMUsmiFhr9hj29xGkOZGQ
4mo7PMJZTx7P5lGA48W5hbsvvOTUwjkC/Biil51IPv1mJRTi2cdRAzXhZqALLBIVnxLQbLt2GiW9
fL4hMQ8QtqKNpWhiOOKguKOncAa46fpWHPQQkoSuHMjx1oWHOEwvUpllg/SVkqOSMfIB+q+/RX9p
IVTJf1EOHRYCOdgiVFSYOkxIkYm0yFnpyKl1X3ZzKzF34X3Hlm1upDx5dFnBbgY+nqLYTedwOCqx
fCQG0kvgiAZlMuTQIK+oz696iHUDStw6ylJ8Jvnw0bNtm0eCRt2xRsLalK+t8MvnsY7i8fLTMjRr
LIIOeKmH1PFr58XUF7Sz2nWGHDmDCsKHCdFLK+5Yait09Ix4dVOgbCastRPzWj6EGTlJQAwIjZ08
7XW/Tnj9CeXxF9itmVCu4U6EOQH6ryMeAegsIkOKAPqtGhF3qM32o+UTcHpKluV5azhUCwoAlCe0
q6mYOurArP6nwNo83KCbn40/wIOgakaGND7WbBZ8aY4UoVBvZrP8RlU/garAlMbOKjbORnS20Ukr
552ZM/TSzYl07Vnu8OYAJAn8PJ0t2aoaPo/ruNC2GDHaEhEDzfIG8K8GdYfPrJ6hAQaKUShgCXL6
LRvG4IO8ED6xtCqfmSPIQjJh62potq5je+cRYrG94aVWso4F80mf4METqZ9rxdHqEfAggfgbUcyr
sZlloPvZf34ONYIJXGj4PCYvDNmprDw5LpeboHRvA6Cd0FFSMxpEckzgQvOFqNwnK71ZoiXE1RJT
MR7sr4UK+6fcDf9rX7Uin3PfcgAzfPLRMljyrKg+WayzhWlXO6b+kFjYj/Q+JSUdS52HVJsvGzLR
VZfOsZZM2yrBX8qvErrSdJdpJ5rC8ZM+LADe61p6obEjPaN8vAkRj1QMh0uHmrcmYZt2roh4X9Lc
C5PSd82g5FAIpFuHdyiyqg1Bs5wGhdYsXM7YA5NMgjBqwrWQFyPjaXE4GNownk13SykDD0yzQrNb
+Kz5lYs5TiX+JdMQ7HE83KR8kIeKHJIK/YArrYzY0mFwA+uPN+a7aFlHdx8soc29CFkuHIuQGd2o
YjUizQE15WVZKoO5ISUVOuY4sslIcA5KLjtdrHgah+DkvstjeQPwb0Ef0YHPcSzdxI1XVyU+wZ6p
RfI2dxy4IXA3/W74iFY2SYGKAxml972BsYBzKtVKJ+B/zjpj0cIJ8OlSHhR8bOT9uLnD+ePmLnzk
E/eYT0m1ZYxSsMK+FIOyUMRiwzaCztpKa76uilB5PiZH2BrnhhSLRGpPvOVuC1LRFVOEZziQIzn3
UiXAXNTCHTTWidufyVKnTjlsGkSXfziB+hov8mmQo2WkaG/exIGIobtJTFXI4ZG+hX9rOYhCpTzB
DF0PYaR+XgdwFO+adkNT6O1asu7PYUCcXHYuCJqWsTt80F3gt46dMAv4rwiUckaKUzTDEYnaRbLl
MxExpNGBkB/nclIr26/mE+wxiOYRj72BX2IELH2MdvJ3BEhLs2KfJIHm+Ws+9Quu6U7qX4dHcFSn
iRsd8Q+2OC1Y9Oid1VkU+Ao7ijEbvFO5EzShU6/tiPbWOnwZiyF4RkCzptuCStMm56qRRJtJdUqY
pP/zL0940Ys2IE/9akLwI7siNqkH2mnx3DJq1B13a/Op1hHwFTEKUn+d+3qnR7cG6GboqVhlnVPu
ejq4BmRSX2siRFmRBEq8vijvusnc3xj8lFlaIHT0iU55dAY/I7dap8t90LBk65/gUVPe3qUbP5Jx
k5/GXYO/sgIl8w22IjZCorcv4+EB5UGyj9xlLw0CT7266/AFLMvMmv5fkUDkJkHbFg4J/ny/WrrU
5y2zQqRvuqpUT36qWWFx36RPICFugwj9YtnkfNZTKLWrptRjmf4KS5FP6Lyl/U1UwFeKm74F0h3h
7N7K3ieJbCb2CQgA2v85vpbzLBTJSHdBuu51NgxGx30ktCENiU8qfSdgVKyJdFZ5XxZmiwIk7DUz
gkUrxM+b9DqHQAMGKqegDTUFOxtDwH5SlsIqycZ0/bf8QVv4FY8X7bJH1iF+VPjOSSn3vdrAxxQj
9bU87qD/WyShovg7YT5PfyjHvtQsMCiRbPiKEeZJF0FYVqtb0uHfuUl3rSwZbZoj9jfceSpJbpUs
4JtwFsbh6wEdHjZrZFbAaNqBp3Fc9zoqJWowcXaN+BaywC8DkxM2SWNfYSiUNpyxH0urVa+6ogOd
+SATQ94q/zILOWEQKn8cQU8NC6ecA2Kf9y77jOW57As9z8BJ0PftWqeY61rKist1cJbHyK1zFcYv
C09kEXbu7YYl9C97zgRRySznJSWK7aIMxvjQ+s5nztpeuzHfp+By04l8DdWdnFE5lhCnEHkb2q8r
1PzAgjhE7XddMS5W8Tj7lU4B3iJxMdSICww7IRHFN9edPJJS6vymS9AWl7L72KKmYppdlWoZbhV3
2fsBtHvtfWYDTVV8gVxoMLVLnXagsXNOjGXIzrIJbMICXyaNbPTjoSppGKkfbqYw7fdYizvmBal4
eYrUbnVoW5aaMUihR/5aFN19wlSm2udR4y2lh87NAjjKcpTe9AGpVYmL5HPkSOur+XnSDEnYn5gA
h9hjR3WUiZD6CsULiQsZ8fO1DJWNz+denyNBOcnOE8WmQLXl7w5U6l3YEu5Jerv5+r0UWMKLypDn
a/ud/qhlog7HR9ZDSIpQT6t+ZqLktwHfYueRvnZdKLI2odvj3Trwj0NNfHwyDzqQDV9hmr6FUw2M
XmfiyeCQEWBgDUT6kt0CKu9GDUxeGBikNsfREqu2IjxGp2F4E6YhyF6TsB/IfrhjBvcghL7QLVEa
48L9WfPkLx1wL5+/UXQcFVfkjddKmajatcWgLNPfZywF//m08iMijV/qZUVgy4P09TQ3ACwRk+8h
M3tfSZ4MTHtTE4q4K7Zi6wnQ6/qtWSnYPfx0HzY/OlvSPuDHZG4ZYK5bpxQIfqq2FJIuQq6CE1ew
cczjKNEA6mRynOM87gd5DOuE2qztABE4RsfsHiLln0P+M4pirwbpnniAWnNXwL2JlxJ10DQtcbjI
oHYB4hl4GgYctJEpJYOADJv/5II+vatVWcu9/Cc7/lMbJAScnYY6vR3j9dDYYcfG4O8s9arQz1mk
TUggQy0lgjTfiB723fyBoeyPU2CxDvxVGVht6PDHcXFiNspBmSvFuPpAHOOc2T5+C3pZF0gJ07bM
NksXPAv6gbsKn67ToOs+gQiwnPSLDUaEODl8WbGLNTHsSd1k8N2CJT7WQ5DZuaBqOxS5GhiRyROV
/94OZSmpqTUbDdlVdteZRi961CnTjo8i8Kn6UHxzNnmkcFaCqAaquxNVODLfU2pbT+ieQ4PKr+//
T2ENYTuC4cz0UNoAcJ0X2wI8V0kNcgJGwGWBdar54lx/QvbO3l7DY3lkxP2dXCdrB7K53/Tdn6cc
pNU9Tv1DysmhcFYZP6zhTvk51tcMEOME5mhFMmSqqiPRC6zkArD4cQKq30YWRd6a6BR+lJu267o9
tGAvhDdNve5nR68cZBpNNmpE3t/I+b9/oxFBbbbekk4h7hbvPDkFB5d1AvoVEY38nfw7nQpr+Qr7
cu2TR9mvDkW6m3/4c+aDY/7V1RGgWasl5nqIns39F44dccuxEmzq7mqTA2TQvlZ9gJefGMOqJo1c
NpNuvqEwZew24Lb95W0gKKGNVh6QSxT4EJWw3vMCaBMxjaSfcBHsLNctUuZw6sMFoHLH9FO1bspW
rtv1ZBXRN8h8/FSSc8RTLJl6kWgUfENZ2GGo46b3mr8OtGFBKg35nrnPNPBA78EVBh8i2kqWKtiT
89Mpesh8Z2sXNMnfmhAvdZsUEGTX6I0XlrPYH9Yhi/6+QdEaqbqY9flVebXWN66zVYJ63PaTW8Ya
M1jT7zBAJnpp/B46NaZaTZZDX82pC4o5u7ahYLQ/6N0mE0XCi0GGrAdcBmwL7mRtLgdu0kGv6OxC
KJ+sz23KJPmkaLpSEaum+OP8Q2n8rx9cATb4ld7zYtoT060zYrZme0U8RBA7M+BgSeMtz/g/K9bp
OMvl92vZCRVezlA6bH/hhuqEuwPg3TOVpEcPnr42jEE4fE2fSlvufI+jdg7+A1KyUNqxn7NaAJAf
umkRlAlztkPp+UUN/2pQmoUu6hVa76dYZTw0pIzU0xSrqNf/9vIGsgZBfg2no+3kzWUWA1a/gmSg
Po+7UGK+d8IgCqJlkk5PMDE2s6UAh1/dcAqxq7XR8vvPd8RYChhOWgbcJmn24qF2eovsh4R4SfcD
naUZAlFlzoaEXyjmUnaieGBNfnn0WXIuhGkHqsvDBH/BM6WOdto4QUp8ibTqTWQjIx6MEN3M3eU5
cw1ZSHO2zP4j9vuu8aG38VeWrUet7EHqGPGlD5GjKrXIFBYcCueQD2rxT8DsSs6/1vFxnzYTFPtK
DTidDU8fESHcxvyZ/40Ap7o7GFilfwn688/vVYiTGcjbUj2NW6/ufsfFqeIE3zLjMjex6Fd4Ljer
yWXGufWKdpZdzpdE4QGiFnot3vSSVnQnUEgaO8am8E+k7CqCrFfgVI0BqHhNhBjFO3LS8XugZt8b
4xS6nxdajXaj1B8yjsBFzyRkPmOlnt1PgybK1D0SFqmjDRmBQuLrWTDHBjRWtJMOp2n7gCphoe7d
sqmrcPMYh/Eph6Lac48qbS2JC+yyr+FO2sw+W6sD6/iViiKRc+CmvH/HnS5x25a1xhNH033PHEHQ
kB0bOY5T1wi6v0OUexjGyxJehKfYk/1LW4fMxd3cixox6GfA1O5iqnWOLeSt6gcyXX/+BokOquLw
2X2V3A9WqMi0/ECwRZPEPxcECZi2Z3mMDYfv3+hFmSjaPKi9kAhcdIEZ//p4La4y2h2HiUPt/iSZ
NwJTUks3VaO8OKwRjKkqC6H7iUVQ5i0nBE9wWiZNN9ZjUPcGJC9OyMmRkNpnV5tXyqhIyhO1rPbA
ArRlDu7Cm6BvUAJih8k+0ZdTa8beOhkTg9v/mVPDIvL1qO5Pm9pC3ArAjitfAXea9bUwm+WFoxLL
6KF9Osgo121Ircgl8pffODwy0srQZSCDyMRabMnXZgSYE0XJfyyDqGy9SQNDP4Lzmm0u5SUgT63C
ZX5s37sw4WcjHfhAi5SIX3xxaTyobIZ5RjfUTIb3UXmZp+1kXSkAXKnMuFp0oISLP7algnEZEAuQ
um9b7LVmJkWYv9X9xGjPU4toBGx1eMpyjaZo1yybd28OUmAPdo2a6Y4KaPWPRShFvG9zuMwcwM0Y
nLfdrg9evmA4369fkqr6w0Y58MCOSA1QghEgY103/9NDIZErqDS6cYckGqQAKazqPTkPPMibOQCi
MlauqE8bPmSKC9hw/9FJB18dpOJq9lEoZux1+pgc+SDH3z/AOQ0PaLYTpzazCqpJJDYlV4JnYbFl
uG4WfcQj75Hvp6grVTKXqLaS7lr0iAu7dj6i/QW4Mla/zFwx6+Fu0VsLQ+fYRYDCyOOPu2WUOb8Y
JMzBt5v/R0cfuVE1InqAsBp2PKwjMcugH0SF3nX+MhWixc++oOVc74n7t7OFVZH3yTr2l7GgqFZb
LNla03Dwpi5g1Ywst0WWsDM1Ic7ANIszRt7Q7IQDyFK5jBZHSod+Tk60ATbd5ME6rt5PR1ngjssz
sV7Ju5cLVinrNlD35FZBmmW7zz/LfL/FSYR5Wl9JU2W0Mb8HayDK1CeizOeJMP+elP2pKhy/7pk8
NxUfzImI6UUCYP6TCi1zSIcRoNGlW665nDve7jV1YjZhkbHcq2q0kiDE+jhTMuTBigy7xhTeypSI
fA55VUAIzSx0iVJ2R1AJXFr7BnFwaWsAO2fCEQBAgTXnp9Dd3LnZr/Euu61SV2GQJ89U0fUN2fzV
tCIp/PgFdRwoUkbJkojP7IX4Sg3cs/NDSxO5B1QSzBQsoBwbK0t0Z1UYP4CaOGVmIxarLw3V7tQj
5FefXr58NQvi6CPJPeSOUlJ8Ij4k8mbKI7u9qXePCKpAq1zbBkCa/Hg1QX2xKhgvVT5YF2++lE6d
YHmabx6obdhxDoXsWMQS/yobfgEzq/zQ3gcvCgA7aTSzjoxZgPd/TIKv3EYocYFnr4oeY4eRQqOu
FPkm0Nrsq5QAyGYGrC9+41fM6tglKZhryCNls0PmWjFEm4A7xoXAbezgm0cpYK5c3M05OzXg8Er1
JOaSpjhrxws/0AQmjX7QpohuLhW//u89EVRfKTy/rosi+MIbiqY9ZeS5qhNXnnqNJ2ooUHh/uM21
KGQ5FyKyFH4IFv7dbUh9Zz/JMoExC0scNFDKN6Cjbo9qSZdXWiqmmgyL2PpnlldlWBb+w2cryLbq
ePWsWI+Ch/Nh7To2wFJO1tJbLxX9K4FmZkIb93nsXh0wrwhcXAgduJ99MtYkrPyhrtZViln+8lYe
nWjvc3XxCZCUppUwBAnbPTTZK7auhz81URMYNB10XmAfmjePdtz8kRdYLJXiBeD853oiy12WSbIO
/XvZMWady8eprvzm60sPGaDecgDGT6iIxQmsTNCUB0w4q/aydbywP+Xod0DxfHTIK5p69ci2bRAu
2lXfQme3cQpU0RRXmlhwzgrMptJ3zhHj99JpJFSqo2t3Yl8b+tfzsR2PgCFit7aQU4wTGxHXBV2n
bypHaICpc86dH/Xhhx4xjGTX5APz3AmPrVZxMiw040IMTE7ThQutnO8j1guVB1XUuBO2bjLCKdtM
2qHmEq51pQZw0cPQ0VzBB2HAqzELG9LgMFD5ET+zzO8jX9W6yTE2EQT6FBlRsNe8WFUFUff8IPol
YEOZgjZ2GCByxuGYXdPsmsAonCsceNPagWgO2vtlAxUYa+ZuSJuCmG3Ky7PEDz1qOPTbQKN1dSng
YqThzvHJazwJzIpRCEPc0GDwrUKENA6i7NhI1Af1+77LEteG3QT7qStbBwT0Zh9EaVZARmbJRatg
wPlOrNvHh7xEBTsfK6XZdlxRHCKag5PI8QcbxPDhZVSPmcW0jQo2gSmonQEzgyoa2morRZeAOBhw
dSqGMiqyTWAGnIKH3KqF2wNu8Y+ZLhcz5VwQSxgG3KUhWxn8P/EpRm3npK1LPVkgbNa0+mn1Ul2J
OkJhK5tA4rNcCnljIyR6/I3eHsWy4FZWwlXjt7avB3lD3j4/UG3wOMEl/pLh6kbaJreJsYxppuPj
8hql52yVJOJmw4AwNh2++Edl0VrkniXynQ2IzjPaffG6H0ji7yKddi8Kmy+CWCKt1RkPC1MvUFEC
TpknavQsyZ7L3fK+od4YfG0bLqdn4S1O6oiJoDBsvcG3I4wl5ANPRMZVeTfKQM2hx/JBxnVMMTJR
40c66KS1AvwelRxardNYCmUw1iE4/JXWeFEUEmYq7rY1oqOkkxQODsdgBFcSY8DQ6XFc/UFERBJK
Fiz/WzYrQWBB6AJg9zzVLLRjVJLIHKuysrjdvkRv78j8tq7V6D80cTtGa7vugu1kREYCCvp+Tv9Z
cbDyg3uJzmlZoM9QZmD6XSqXqARVPzzhF0UnYWqzoTJCYgllXvxOGeFon48ocv4AO9mrqKUFfAAw
XdJMV1CyoL28OXHRma4J1YQBCEIV0rGcArC9vqBlwL+b3Ed+yGPZgz9VBBsIw8kBccAbK1iiPJqB
pRBVVLfQmMMcL1uQtNEZs847yWWTbbqDxkiL/3pl3XBBkXaCukVHuN9iruOPK/Vp0mObpHtLy8l7
OxNYUj2zmu9VU1kimq+IDsL7Uri6+5AWxprLiz7sLUk01BZOsW4qB1qut3MRhs7KCKEhF66CdSJk
+GUZ/z5EH00npq9vLI//wcAPsN35YlHCVx6VQa+Q+kWLpXqOuwCIJuM6aA79wcCbSZucXCawa0Il
VRZoKQvAqLWpkaZsfi/sg3KdjNP87Tabvf/qbX8soFmKUFVotNEaaXNwFHp19+atYo3jD+1d3mY6
jFN8N9NfsB/+9YuB8isMp50ewE6EORrES4nsKq4G1+F0QGs6ja95BQk5+ZccQVnhzGCIpHC+/uq2
aaE3qARiDjrchzCcvFFLqf58Z8lRCZ6bamgk9oc+EFa7dyQvsy2UHtmOp9cEZ2UmJ3veXpqzEi0b
75karXULTbk7VjZE125pyaXj0xculSXaIUUEaG5rEyCAO99DqUuWXznyHdq0uSwSOB9l9e0XAGZn
q6KhehhhT07O9HS8U0ioaea99/FV+kOLvY79GA//5jPRYwbduwcd+yGxwsl7FUuD1Td7VVVITncx
Z4rNU0LjyZzmf3FB95RRL8nf21/F1NdKPgXNeiEwywbYTHimRMIrTLeuCXgeCMJ5vVLB/y0X+LVt
ZnJDMVCjYuBEJjw7NhUHw4y0ieGo1wFcJWt0n0rIU/xb4+krQpDtEPp+eBBBZuy/KKhmjNuwQZN+
YTDUYiLAyOTxqj+5QiuxchWquOxaTVuDmNDYeT6Rlq7olaaIFNnbqSVBPXXfLOJ0W9V1GNkZdLs6
WeRf9Kv4KJY6BHoP6/Qpi3uO37XD6yiCectpZWb/kEWyTXZSYTQM03z165SZWuaGKhxBxBZ3NfR0
MescEsbCBMcfxmSJILoIAcb+p8ZKDxetL8PQwCubGfIlu94z6K++wBypzhm8JRJT9K+hLqLL7CMu
p1CMV0YX7DIwsG2uD7Q1ZjNEtg/tKKCcN5e9NXyOKNCY2KJkIeikxmSLr5YuNdBXYG1HFqQ4AruX
oarUzBDNG9ed02WUZCIVwZviYQDWbgiksJMNBSXFdi2j7X/jGELzgXdZVm75XuXq+DAag5wfrRp6
F7VpzFl5mFtjrtrwk6W/B8KSlTjc858IFysufsag/6dHx1ql+EtqoFLw02cfYD7wmsVSRWquC070
1kLPZnThOcQId2ZUsoF4IXANU2yzGtj9zGPujsz5Esrm6aeoQqihDOvPX/TyBBwWvTIsMkOWKTnX
UFsrDRwvI0r63cEITyJkiJk8B1Sg5UwDbGr+4ZTimQUX4zDCYfHGbIhbW0P3V/Uf/d8dXO3x341V
hTQJ5owQ/5CkfNnVQ4KOH5mtqDSdkUACL2Rcte3MNFuEMvFmvMe3NFBvprmMBfqDTqihQrOP8aEH
Se2CVZKtNY2wYIvOG63rHOIhzhGFZg1CZulcnD9R8/dFUNMry2IBT94az/IG2Pzeqq2DCzWZ36BX
I8zKwBm2OnmReLvQ35nMyvcxtuekYB7NBtRDf56iXYx9tEj/m/dWaUSqRPPGwCp1xpvwKX7x0x6t
vdXqRcfDcmyZDJx5BKfzrROr3Xo5HekrAbhohiVcCFD2BHYP3xIdO6DNjuYNPJJNJk/chT+NVFse
WzqVUR8kE9wfUUF+9D6f5y6bmBVHEqFhZumlefEnMnJCvFIJIuJ2UnRrPt0k39rDdISgSCqTdJVZ
3+wfcfKzIVREs9V6hIgVRQroFNvz/rxPLyxXz44MEQPLWcxr0egbMVeiCg8jguG1mOq2kO29wss5
JTBVX5AB7FuhXCqSzYIo1kcHYkgtLY07VgtL/be9JCce9gCUzMVX6qGiLrkZACIBldrfkWD8HGhH
1pjOKolTapZ2/31kSEqhBnmitxgcWq2h0x/BeXgn6RlLbsuLfAeSsY7xX9D6xJ5CNK9gf/cmgh6E
LNVJ2cYOwQ2z3UJFF3w4tnX5eDN5xpPD0pLbwn9tZjnup9axDKIf9UyOb4CdYpIwNNCNPcUaha+p
fzC7FpL5RFC6T86/bSG2TfSRS1CWOXXnvu+uCEAkAz8FKIKM3ziqobTDx6Ho/7Ot3r8tlcSymhHi
ryZFQ/JaEZveVUopCKZaHwrqlXSROeoCgOVY83kC97Pu7mFacXpONJ3LFYgYqUB3Fb9/ShG14bVT
ykhaSw3oVkjEBVpnj5caAaeGsZu1FzI84nfQ+Qjni1sP73ywEYim22mWgfLkvhSrzgJv8Rtk/8gX
0ji4DI7SjsYWW7DDFKfByXOudaSSL/E+Fr2DkkV4esP6hpwnR/Kl9WDsDCApNwwYiYLNIvWXQsyH
ZpEiiGaZ38ufC0Zog6D8SSUCn1+2JE5oqdh/3ys7vNbmhcBhXMzhES+YofdC3/U50iAMRDQznVn2
rHImjlzRDz9+FTAUWvMdZds75v4KXAZbcB3hoxqijBghR2hou/4eOUgwf0mXFlAMqOYjYTN879b+
L19WR0I+3HB3Cz2FpIGyLD/USGl+7zTiFQbTJ7mZOwnC4XQsmdK5v3Pr2zh67cGKDB6W/YVsAHIF
TjPsCUzf60DepVwens+2kAeJlnZWGEvr+sbaZ7N84xy/DcXEVzOVc9Y2MccGa9wrnEPyuIwrUMEo
NC1o1VWenACP5UTiaviIub3h9SmWqzdx8HwtJS/oVFPnu0dZX6l3sPwnDX29kMskiYGXUypmG/vT
V1ykvo3zZ9MDWL5eCB1hYk611yZYz3WUqzPg/BBCtFTSYXjPE7TVR3Pd1YB64VkmKy1UD9zPdgun
Ww79g7zQW2x+zHTlTBQ6UUryM3IuONluD+cMI9g9ePoQOlbZKB8pNwsTdt7es9nMXFMqMtf57rnB
XbgufIW0cE6APtg2xyF5e7jofJGTg+/SILXY+exbz1Xvk8HhoyJoR5hzjdCRrOQzpttnvJ5/wJ0Z
uSrcNqUZ8V2Vgtqhwu91AbcDBI6C6PcA2TDvS5ddANhLntwpAzxKeSAoff/Jx3QRDJ7oOiuCCiD9
HnDVReNpX1rBHFPo0rHA2kyM4vg93ftaHyXranRMcEPRpOi4apCq+6JEHNOqTzRFtEQH5JVVjJ/d
8KzIpxsb6K0kMGtpcxIMLDsD1UfodRVZorcHzcrMAhH5kvM3kJ+9jEy36AzClVhswqDz5Mz/MeDs
iMzNGVKs2H4/SI8y7nfW6pnde6saKW0HX0EB0/8CP6raB2mo7IUuID3KwXNtaBtRhhc5o0/z6aGW
SwteNpSKPem/2iHM1ZWPkwrawUzLIkW2q6V2uS9LndU4ARDWMRmZ27k9IwsgFFy08h3uu0X57UEy
XvVTrlHJzTmZ0MqLs27FxE5sfW7nSne5GVzZspdzKQzEP7DI54TVkCzdhQcF+j0+KGTwu2iDhb/V
iVy0maRyJwlYmcAnnJvHUrfyW18CIF1EVPWA3Yb+SuoovYQ4OK+6/U1bIB9827RrYHAdaiCQVU69
8iJiu+YSiqnxh8C/RBW9hmFldMh0IzUjhZGZ6cSOuuYfE4Gp86tS8XpvlMECqqwJvMCKtKTPOfWJ
rczuCIRoPZfVhRdHAk/SRpFoW09A/TNoaAPk0e4JjdVu6zJnCzD94w4+4SdoxMI9mU4BYOYt4X33
A2iAeacYpO/STuwOlgF0daPB2XwCzsrs0dTWj1DFiZFP/7Fe/hYHY81+vVbke8QWxCfZEAgvEs1L
R++YFedVbfShnjqWpl5eq0tQngAKqsaXaQnxCJmVMsafw3O5sO1Jy2HPRimh5599qdCSaXAy7+uR
6jeHqez0PTevllRH/et9tS3kg+ewOSt1Pb7VdeFbSFoQZE1ffsYQcQoYzPFkhWwia84TWwown2x/
Kof39fQOXglLPHLFGvcUTWgml5fYAuJmI1yBw0JhAjaNjpXjyCqX01xtk5eisiOvph9yBhdNUhp3
TBcCGTBSnIFVqCadgSLo7GDfSu+MhYClRmMVmh6lAEC6B3kRHKu8C8U/J02seOLTpAqvmEZF3mvl
IESAXR4MAxQD8TD3aYkY96YJfezOzenn1gMDC23XCQLgZHjZn69BBGVLD5OTrJaA8EDzxqxB46R1
3ZB+3jx4K2hnuyamADpbucDqOqKjJm3xQcaAiIxfpMfho6gh84TmaqUr7+BTo/DoFRUoivF011jv
qmM9ksP0N33hP7NBmgQQZGgHlMFTIMqmyqSJNjaf3Y3z2A29prTdlzNaJEMFltwAbz4jPCvY/abr
XQn0bNdPrUlHlIWRpjb1dAkztETRqJo1HoTVIUugPZcvsOtdI0bGZL5mk6Dn97MF9CEJJ3UfXj1Z
mwwsKG3+LMqgu7EeIG0HMnTJnrkvgPeYC1Yt+A3A22XPx39Fyh1qD6zgTtZZyy1PCZ/TNhuNgr4u
6is0/BtzFOHXfd4fXmo4zWTKYkkZuiMc0wu0i1Y3jvNvjD7D1hgXpcVbwvv/PoLkOXzSqQYehgpZ
Hxr4pBDsfkxqMI0iZ36ecj/6tKt3lI9bspnugMZ5tkwWeT+Yr6fbTA+mnMIN2Fg2hZf83EkUQzK2
3hmzwJelQbn1QsmvyHBdEOLa80Zsl7tc8zEyJmp1q/JQd1zHEbKyr0isQ9HIXBlQfJgeOpycS4aN
9QNVNxV64c6TONh/oMvRPvAWpWPpzZeQIBsywWc4P5SpzdR92XTAzx9UvkRgwsDLMGqjVY8qCtA7
hInV9G3Qkuy2NXzgG0j0Wz7AQusvxntu96Mq0hqzGIdabSNFVgGuWSR6eHelf+aYTnGxFHQCKY+6
ICwz8Eo+vbUqY9dNsxVEPIb1kpFW7AnrBdz5Tqim0OgbKuj+gGfvwzhLPwgS4C7KI3begDyU7uIq
0h6vQ/JnOukH2HTU1wzazH07+nlBzqhXq4M2hCBuLotiwy4zbvrpNvREi2sYGD7tJzEEVv2E60gP
a2vBry30h22osiFdvubdsvcDuPwaM2og/M7s7wza4bhEW/1/uGVK5mkYzTVvbPzSHyXLsgHYqnxx
DGfSMAG5905bXzeYg3UgGc0PlPjvXWHeUHEib7Ghk8UFVBakFzJaIp3IwZJr+yBweHW9sTZYNlJS
a01vGaIPKLRjur8+AFZXotiEyJoypwpuAgHccNWwacqmCGmhGk71FrYTJOB8evVfTyz+PV/RcD5x
QEao73/lrcQAPLazuHpw74NYtT0tW1p+u43VTR9h4GkmDPRn6WYY2D2/2FqeoIog991JiMm1QIRG
4/LiDA8N8my1qsqiIMHEGLFP/JgXNispD6ds02Q9bVOPl+iYqK3yrn6P9Q1BGjjexINcHdHUrtm2
1Jzo7vlT/Ej4mJfrJuMPDO9O57AfsyBUSAlo/svg9zLzn3jPbLvO2BcuYfeF9TKWDSumv+3ySJ54
0rptaUofA6rv2e2LUUZlUgVID/dexyXNN+85NBq2Oi8GI3oynMlBAy7YuGdKMT2j+5SXmh9qJ56I
AK1Sosm0p7v0rENqpPZIP8ZtAEF2xwey3Lto20EtTXk6ahDbzdburRLRBye+E/Qo7n9t+0IMnwUM
tGi63lSNPXRRC3JgoVLHoMZ7eWOV5m77/vRoKqfxF/FESEL+1tDYJMyRgpIOdSvrZYrkWnY41CN4
RWoYHkOorKZbabBaEnP5KvDNDJEBGIQT4wmULPTHmGoC2Dw2/OJwChA92gX9HN0hPRYVNnvXOPyp
sC/lsSO5OtDrileTYfVmfK3ui06hZCTTwstZHbA8knAKhyHK2muTUO3jIi4W7FAjk9AQtL0obERl
da3cf5QlBoLezRAdPpWvgjSRkQ9+2QT3fSHBcUKOuggKD/31SGkGrfI8ETCU/gIgHM++4JRciZFA
V3UEJhXrTCddvgAQ7UcborLeS7GfVstY4xgs12WIIJHCsGME1xwfrLCA12JqEmFm9ERmr6psBsSg
nM8w3itNQlT2dyeULmfmo5MnfgeIWphGEGR7MvjgB7HYqTM4RDBudV8E1FqYpU7G3jiVYILsRwyE
T11R0FXZn8rbQeV7h/GK03Oclo1mTyC9hjg2P1L7uuNNBgtp8JdAtbvrTlxW5C9cWYU1NC4RanTP
WNnazuh2pmdxe4Xj3BllE4wbCsmJFH7RxVJDSrVoQ9pTS1zKkQDXCiFgRYZ5/dv0qKTuoYc/ZGGA
hToJrHDAwWuFieqrwJev/suinFpRTTlMNqz2rLepCFbVeQiKXJtoNtEoh5kI2MNhzFdkdrXZ4ZG+
u2SiChqP/hJRrlJoPrjYoFB9ftqdj3rd76A78bDRSjHDdLLoaAjAVhH9iF6MgwgXw/Mg/1c14zLm
9yc24xsLq4WsRcoaj86+gH5lEbDTEj1+kWSc/uUxNahor4cZCpkxvMFWoG8w5q2Sx86sC+m2iXAk
/EaWQ5rKedvHNLoJBOBtIKEyCeTz9oid5hagE76un01G36R4lppcZq2qzleG/A8PF/zmogwljSpu
gCwy7TXlR5iBa1qR0ABPqjOt3pkOREu9a1MA5Sc2gk0VsKYIBh0B9ZjXFubL3oZqfrwpxuT17tzv
Xn3GhEOS/nyT+70vZwwenNwYWOymBmii+wr5R6LnBSAU8exE0G/gjYxnz0KmFlOPpDgfYAt/p+Fo
1s8ne3Z7HRazoZ5gUASPdwh6epTW6Aa9CkGFFHiqaYX1D3MB3kcnas/ZShsKHgmNNtOGqUJNT77Q
hMr1ggSjZDvf1ngswrSADvqP1IST53yBrlmIqjea2lNTo9tTotoGo2OAKrqh89PBGoFbxfInOLsS
NI9z0ISGHstLEhk6rC4xZWhg6SbnT1pApOgzo4lmPdNwPsLG/XiZmYjKFs1HbfHoH7vWC/gnfWKJ
daUmPVYj5CKiLU5CgVtsOoD7UvQA9kErHCB/idPl5P5gJcHmv8hFuAsM+skMh6lNN5l++kuJPKyf
XOyMuPaDxhLn3SRHeZO3R3S3FMarHU9rOSsi6WLrosPSEE6uzRia8lhb38DVm1BQgYuN1kcr8Nla
yL/PnBm5R1HXKE0YcFsOTskKAXEnb56h+3nvRo78SCaN74lzIlDQk6HHFIIb6j9H9UVLccJiLYFj
IcymNiuYyIK+yUHlMOBRHpwipBlZoi00gi9jgQWm81/J1iOGbG/lrmfrsNCFadznodjM2tm++n63
0YvEsQL4Ab/39hpNOX9G3Cz4CnsrYgoQsDctm0rmQQqKpdP2JR9wlldmj0Am3P4XjHjBwiMxWVIS
zJ2xR0BBEwuKKdvPDpNZuBaAgGclniw4KM1zg2oq6j0LYDpzWLnTpC8h6bWYzIjEXusRn6QaWFr0
bKf5Xx3HETiYVKwdA2qUNXmRUrTeYzME1wDrL2QitSeIZwNuRzXFcDT1WhzNzU+ZC+tY/nXkILKH
yxosm+Rf/Wv/xbuCdgtvn+pMOv02/rQZ5qbMwaXdUpru5XlcCBz2TwlPZ842/FwCofLt7wIMDH8O
H56yCLVvwAJM/Qyo+cy0klWLS+2/McVYe8dE9b1tdl1JBLDKSHT42RRCPmqNdj69ZSPOMCIyXvmS
x6lXzMrB4iqSDaSDCXEBGGeqDNFZCPqCOP6aynq0GHEwAFD9Jou/K49ZeLc/JP3H1AM1rMhjRxw6
EGDUDtO5x/lMq01vP+YD7MKhL4h0uBTKln3I2NhrifEib0p8hEH1oOSGv9C679CxE5lPTm6wnQwL
hFdmNOYB52SqoQA3v/L7ISVicCWVWgjHfNRTYY9A0lQKZRPpA1HZeGHuXQ4GXE6m6XnOwREFps/N
te9Ddzsi19usrlHYtdLZILdSLEUWBIxHkO4pJqn1nBcaaV7sIdWFBKLTw9d3GhWedKN7NPA9Fo6Z
Rf1b/d2wHWIjxevwLYqW6mTpWALJphxQMce1gm8MF9c3cPi4Xz6W0Ve0p6IhLPakYqVG4xT/mZo7
Ags1ffcQVgaOfGhWNLjTicV01bSEFDi/O2sLauqnfxwHZK5HVj056CLsQFtvhRinusDUlKoM+2jF
T4UVa7N0kil6lo32CAq0rk+xzCeHDtQZmHm059F2oQOg1WnZHFXYGoQv3hqV7XTphZ1z39pCJhOe
g+EiQqkEhyKVQOf3nn4DQxtnhVGf0B1DaewMkzFWbRPJE8joZhQg0MmhnXxS8obFn7tuK7QPF4s2
Hpof0eNTPWw3ikeQWz6P+ITi4KQBlJ3Nmo4mIZsbmQwKvuLDkW+vm4DuLHFDoOPKFRS6tRtcUrIb
mPFgnaDJEZw08ZLxv7zjjQj6ML6NejdkFpd0PEZg0O3NkPkq7eqOcNrOE7y2jtjtUF+qzH+cQ8DV
405P0hx1c2JgubaLqugKR2e3kkg8el15z6hCOWFMqvT7vFdWZaCjDaNUZb2io8SH8xmu2vmbiVFx
c7Y3KXy/TzwpT/7sG4qazKDKMyPX6AaKfShohkBux0N5HZ7lnfBHfbMbD4roBiIR43aV19X0a1+f
OtILr9nKrugMgUtaatCAySeDDL2f0+b1n/fELAk9OYGlr/x1AOIHBuVvNvyQZzShdE7wGQKt8WJt
OrC5lJDRJC1h4Xa8aow+igUARhKBVoMZCAT1LRy92PcTuVcs6r6Zy1fv7uRiJ13SFlMaVduKTWPF
BukbeOAzt5iU4hDHGg65pH/WSaMkaMksAjWI24gws4qGajDNCLQL9p/MWq6WDjQxK4InF3DdtR+l
7f/vAYoqCc4TAjf6qyiRLRKyLghD3FaMG7u7N5IThr0uCmtJuPdZgtp8rw6OZfiDdd2E88tVAjSz
yADPmZ1sO2h50/inbRxE5zWPBYwOj/3HA1mZjoNDz13+IIzr7SLPDg4bEULi4UsuHdkT24otlYcm
8NOsFdlJ1rd2UmCXpPhTOb8S7+joTBOXSj+rTdwEfbX6D2F/afD1OennIC63L3kZidLi5i9EbrFL
MkLImY0/oS3quWOR/FDXH4+GrSfAj/L+DrIj5gWOVOc3jp2TVJU+WihYdkaXtPRpbdQgbXzIbzWp
w32aLG6L9kMYYyOQ/0XN3wTic+shenTs/dFUKqfgbB09WOubxUkPFLD3LGCSlJ2ogJz1BaTzWONj
DD8Xc7pX9Iy0itTXZXCp//zb25uLp0Xn9mlopobFujIOjAxQK8oQQx620z0T5aOmqWJ7EKLYNdK+
wRdgZk/s2/Q/LYID+0spoqHdReEOiUPCp5h2aS0SPSm4NgQmSGYSMPCVnybUJ4gAWrIMsgARmP00
3RlSMhEzjLseSF4iJ5E3Dgt/bCdV1SStDXUwfjv7r50jLGXfCt+FFFB8I+E0lnXpJu5L4v9DIsO/
OeYVzcLkAtaWutFaOy5ewXPo30i+sapnaP+pNk7dnMn/tTRrDpcNWct0kK2KmE1UtdTG+u0QxT2B
EC7ZeaudmSnZxXehqfwlGfut+tCPTSpsfbDVRaVkEoXTmVUFQe5vtBAhMH/3d9gTeGfnE3NjGupl
KUCAlfEfE9yLB91SgQ9p4hfWMbFb7syx+z7gksBUHXALX5OEwZTwhx9RwQ3iM1cYVHraWlE/253F
bQEYQiGGh75eQD8qEt/kqF8tw3fdRjxiOTVwCm80OK564/Bdp+BvrlKF+Cho6Yf6xRvh+6NWylMU
S0lfX7EGOkSuX4EBfGPhQw2MlTEsC0vvYdJCusdQNEdiCF6XE5ojejAFmFDVZY3a/FokChFlKn9N
ONFoxb5vSzWXU6lwZzIZTKLoZVLLcYvqIlkW7FRK5H50IkLhfTglBJgIO9I2TRg7oWSjebWBodnf
beDCbywOSN+Mi8c7UguRqJNOdHduw22+rDqUYj7SeJrlwGZhAuWJRyV0GZUnmonOBI3mCdD1qfzv
+hfcmfUCyaLP3V7wp3wwlK08HOUjEAOG0N+lc94tDcYU49Hn7sSJAQdPeYLqcWvUwxr6zngOJ0IK
/FybVULxGxVizFIY+YOvCeep+j6jrFz6Rxj/BmwuDsfKW2SOoCCG6K6VJRcSMvg59bpycYaSNX6x
BVMoCuUxhhIdjfBt/QMC5plg91DfDIYa80dwzeSkvl+OO5F6hnmOinh8cvVW1HM2x+QsxWT6YaXI
JYJX4FXrXWS5Z9nKQtFvQouFKv7Dh5/hN9weJMRP/iRaZl79YGlvCQnhO2MM2eF41+XGA7/ljfMR
AHH2YuULTccgLGsUaKuRbsm++kfW4XHC7QkoFHQm3JtEkNLk3W58rcnYQAKfCiQe0QYwAIT8PKFa
TaGliKDCOg4qAdtgqo651+pJmxgW3xSeyFX+nLXppyHE2q07zkJjMxIu14QngyavFvwkf9q2P2+u
Hb8m/YDhdoRWRc+V6TYMDTDwHJfdEUkQhEPUVqUAb/Vbz9aNqjt/gUwI3sd96fJYIEF+L42HM7g+
ZmEPdgAcFU+gz2OmWuC/eZ8M0Njd7XRaW7S5MDUg4YsMeg4CQSNHvTzqo0TD0Z0MYKe/+Esahg61
p6lcO49urymwkLUnP2H/OWtuf3xS7eH085g69wqlQVEGOcelYRVUfOmOFWZ6ywRrErjyygtPS0xh
3W/bc6ZmksWnUApd22jgUzJfmqoeIFAB1YXc9aaP+E4dYMaFUZ57sITSGnjzeHTkqCRrNy6x7ZX6
0jtiN9Kbwac/K7bjCKXTqhords/Jg/80zyaKWWWyQfl138pTSRZpofszEOaHvDJ2iP86VjBKNPdS
Te9vQajD53gfYH+uLPFmkbDoN1jqm5bH+QniB8zIlmVdibtj5cwWIO3MD1auWmR3Vp3DMcon35lZ
fgwg0HMIhjxZ9GKv7y6b844beCAOr8IqZRH+NPX2nkBRAx+m50CNwqcW/K4hGiyaywAx6mK7FQSn
Qe+o0zML0Izd3cT0y2US3Ul9qDQfnQoGhyWX0NRX6lrGMVLhRbKMy6XQ0c8SBlIIdBJKcj/gXIif
zsGMAMFMsMMZY/nIiaXdmeFu3/Vw/kRLyHvCStESnlDEK7AA4jzInJuQlwhCDNOndHWVyHDmE7Gz
tKsA5/1IHN1tGoyVO087rFF50PMPMWNPqPzM1Cn1EGxbxIGax7N14XpQQicSnukSkxPw82+gOzbg
r+h07YMW+IlhXgDK7qfaJDeQXzxViMcPMaM5dgYnlP3sFWbC8f/vd9xOK8tQhp48ndb2lkeDbMgU
r7l5MCdJsTZKpqsJmN9HQ4+JJYBAwd5GxP3zeNSuVkGjfPidDaT+7pk8467vSUILrJqIXgnwKWfe
H3gyYIJdyS3RzVUXVIyVmmuJZgaDCo8kPXVtMmMASiJe9cImX8UmHixVuw0vEyofeBnJ3ByJB7jh
J/I3D4ufha+9UPgbgu6g7/7kQPjpqm46HxVTBfsgzBfQGAJrcF4UQPnLpvcsGLpnT/4I25+Cg6xs
uYKUkgooxNDdhWPRTOiowQu8t44PPs/fGCrw1ezG1bNuyQpX65fUzgAabibEwa/3eKsuBtERTkWX
WaTfJyInfV8CYD+5wkrIbs1dIHDLoDdmmq9HUPqx1n67c23qgpAL+e8S9lqueI8kP24wnebX2MPv
8pvsIdqiniQ5NLPvAs4If/wLt7OaLdv3GdiTJzwMBT2SM3qZcKJQ8bngsn0HxmQSwdgMuNm4rlHZ
X/y9U5VP3XhGrglqaEH9JAylF3p156MK8+EtkAr0DBvUMiYwhKMvlRX0mGTnRBvqf4dUh0TxOB8l
gViBKME9UYS5YuBTjjUAxCRMu7cEwJpNNvLhtgs3Wzk6fSIRCv/tDzTUVRJ92FvTkE+9G5YS16Yg
apK07NV42h6EroZJX1Gtn8zKY7X7KbtOdRWnmWPDOd2DrTPoMVjS0Kn9JHHDpaWeCl1xC9QGYr0M
/ckB9NZlt7a2DbYK5kmrim6VVqN+7b1sSfjc74/gX7pUbJNusdsf9RnZv0ucorUMV18drb8pZn7/
lmAfZIsndQh78aZJtnkC4GaEGNTyLDSZV4dOGk4Vca9h1jS3V5PHgCT8B+qIZG/Z7YAWBXxXW2kl
6bJfKkL/CGbUTGLAd2MdAal9WAS6YMal//2PxWdmN1KHpGZ4GpYHX+CAn2vt8NJNWIbl7MQ4NwQ8
puRVDkLUL4fnhSiQRR8a3TsL+ROmm7xyV80L9eJjskHpNi8kk7B1DnCZRWKx/td4S2qTvaDQ1E8C
r0Vo4Shy4BKjmhyBATBYALtpNo74s22G+TBD7u8VqqwDsOvC80zzzA1p6allB92oROZFDuks462G
yq0bcgloBv52PFNx2/he3AnDCDAA7zF4K8hEZoBQubSvhgnZrkvPpKbH7KfO0owOjd6fZqCxULY3
Pwxa6M13xYHwIv2TVaPldO3oACC+oUaEu2LzTxRII6OQAi9WgRYxABO7C6mGqg09uwR4I++IMbPT
sxyQE+QdHIHyhMJ6DGzIDWzEBLYbg9OD5d4jbDsNmQFVRH4PbwtA3iXmr+PBd0uybwiKLgTvoge5
7Hkn0jlLnSDepXBCmLjd4CgYM0xWPZMe9FysjhjGhVEOHBOqpv0sdB52fhRMeasm0SBL6ahs0Jsk
r7NlOeNOLHpeCjnDrbKvoCdUloIi3N4WkaqPHuDU2wRbYIoL8v7aPPLgfcUQQpBGW1j5p0ozCoQE
wmFFhucJWXH7ZCfmx/R7vtR2Kb3i7t/mPtGDDbvCr9VifHkImgGn+ZLQ6wIwFvBs5NGs8jyyH1mj
1xNQ/PME+TzGxe4kshjjgNcYeUrlbpdGxwCZOUBR+owHHG1LuqmSC3hhEaTGETMEVy1uPOX3JZdp
rEaGp1J21SQRnyPYtJudtgaA7UjGNWtKKa8ZCj9IbCX97bFiIZXpUkiaG/4z+GL1d3xZH6xhVCBu
enNO7gxIbXKs0+EtqK4v0rDGYrTTMh6yRxRBNaASzN2p124VQxRG6iJWxJYXSJ5StWS4noOzEIDJ
llHsSyTM+xC8QrNYtxIEUNHMpMx4zBp/XeIi+DEnHNZck3Qd20tpcXXoge1N9cyx6+a2+KUGNouF
F0+hwX6Z0H4AfvpZYWSBrmdvI1JL08j+ERtreVM0WtRD5o6HRHd5iP6sDGkc8TSqKJF7+s7ZgrJo
vEOCbmkRU55BrD54LJBHNiu3DB+TB0IYCbw8ZRGdcPkPwZcKNhXrWo7qjYAjrQdF1J/Q6MYySLW4
T9puan91uc4IMd/zpyCjMnPd7Hzsu1TYv9B0H8JXuWO2Bvb5aTNh0OH1mfftwP0YoYGIzjvSNmJf
LYXp0kqSh2vIQbysdtmheaRMPsL8dW5vXt4pGVnyDNYQgxAYLe7i030EfsqaBM1iW33CGwHzUc/A
3Q9xMW65HrxMB2gQ+3upcImyjnfN2GmYDZUhXCNM3CrouYU/PPfWJGq/No6DpdQBuWeFya0jN1tO
+OtKhUQBEkFBoArs5+NFNpIXUnOELwLXpJctwpLBGS/P8SuyEbSplnN7rfCT56TDEGvAnZ7RR0uN
CmQ2EARH3judHqJAkYGaJuJcQ/0xYP4QziQpFtzm53F27M20/R+FS+vxuTD+jIemAznBF14IlqGm
eV7iMMRle3CYvzWRrFDH6Rl3A0Gd53qamJyu4yACGyL5IhxKWFoCntACvlaC0RKIVGSiXoz7YLVQ
tSBjstZJIDnKPIM+Zw0dQ/8G6eTb0M979KMxEfJ4n2KhcOaRb5Gpjmk1sCZ1UHCljHcjrYi3xdNd
5c9m06Edv/U2WExvLGaZ/PltZLpBKDFX85hTAJP0Ve5uG1P3RnL0Vmr4I7cIMHP9owufEaMrRlLz
qaEfGs7tGSKYI1DzMPKRuXreeEhdXnx9L7q9bFCB9XaWXlDQ+aWDN9GoyRFM/rBL692iFMr70WCB
EYWfOEOM4gPWUgvA86Unn/i0WVHhK2cDwALzTWGc+9Bi8BAEF5wUYvDQ0UocLnIpByz3v+sgnV6b
zatKxs7siptCcZKbQ0K/Ijus2UVfl0HH35aKzJy1Kp0CiA/41wGKMQyl66KLyhEZKbkC9V6+ApNX
/Xm38BgLEc3slhIfTIDm73KwF5972htR++vvQZDehXLefuv0NGBmvDd56MRaDKc2S7TlKzuNrFEY
NMlspxymNnQhDkNaEBbpGMvE5tPlN8jQqRPn3SJPBGCQFRwWsjr92IGzxfhI0EW0X7A7dh/pLi0p
ssA1//17A4wXWZ0NOE3mIs5X/RiozFCBboP7bpbpkHE/GtPLFMHosQpZIH5DjIrSrTKVrKLMmixv
Z588+We0oj8omwOMFTEGS+a/n+Zg7cF7gqWlqPBTvVPcnZjbSvtfSfMN27eNWNJQ0smrJaIwQAF+
lfxci5uFxCYU6ty4tOplIs3Q3z1cZagncnQUQS0jtdmwrOsKzVKyTahzz7gt3gf+8wuubg6GR7g7
c9hy35UXCXEmMandBbSNbtcfxMFqaB8j7Ve9y1G7sQu+k+JdcnR+O2ybHbo74gIBKgMSTXsT+mo8
HBOgxLn8TvKDC7joQM9kvAwMwI1y7LbJ3omOQ1OxaaKSpXJmwiZAimjrdtRzLBA59gDk229jQ4AE
x+KNwOU2Km1Dx0lEdpJQ/iUtqcZxCz5KUC9vBQGPQJbdw9qIHKtdFnHKjns3ojxeTYLpHyxwTjk0
O5dGkShSYu7H8utlIO6nGXq5zQqhTZOZFTcnCgveI9G/osxkwKh3Kardy7EIW8/5kJvooK9+PV5i
2Kp7DggI5thABuVd7IYj56RkqTOkJWvapsMjZICioTTk7CF1jmDieHW+vJzQwvqU9eWv5j6x4W/S
vbofAKp7inmu986bwyj501AFOEV9OKO8N1IAUYtwQxk7ljXIMbEOy8pP+WWvSEDeCzP32U4qnUoV
aFGoMggr5NAOAT2ewfxPVuDQ5Zmwn9ZmpU4kU5y98IJmfrXt6HdiGW+0IMWiSCBiCoR64B3izVNu
ZmKdRtSbww2/Xs1tD6klQNJaLR8J3CyP9FpY1pp19nsypqEWqsqo2K2+cqUw/KwXKwmV47XpV6rq
9PZR2OZX7M6IQ6kxHVOpjqg9H1YiZilwBdAnX88PpRPSfiizm4YZOU72xuPRuWJcMgLi9W2wdo5V
0vK0G6wXK0tCZ5RYa72nFH0n1efwEaEZ0TDf8lDui/TepPlY5NmqID9obdzAjbwS8bLaCuHJf5Rt
yJOEV0B6QaxHlrK5/3QcKzR3OGAuFX8KNpYIUixC+0ZJj9pnUE3Bis/+t3fFvCu1p3/Qfkb0pfyl
xmOaS4jm+ScBNNxk4+NYFIpZIsa520WoTCesEYjRYqLu8/w+ZfKm4Zautd8TzqBqPrkFOghyh8fm
dIO27TToUnPF506cBf7Eg/IcU7yhY3J0Br+0OBy9hf4Xxpo9z+VOk7IU6RjuOTdpAZSOxyUpiBko
8rMPHLdxInZ/0in6ZTypBSANSepl/Rum3Zk2S+PRWlih8T0T2n4PvWZLQXtIVvRNPlxAIyDAgFL/
NGlYMMtcBW1vK/NnVRmeaDKqyh8dmr5INNqEJVcRsvEb+qJn8tMQFSfcv3apqlscjHAFA7homEGR
pd2kvJCUnzmkq9at1A8A2RGr+VJGsu8VnFCL+mIJinhJ/O9zD+9x3QiF5wM8RGGkEW+NUNabz313
9eyXnfIbon5xH/cGeuuoi9I1lX2jQquNvZ0UjtJsdnjMEJ2qwhsXsl+K6Apqs4G64U4wJPGmTzij
QenuKieL4As7U3VdoU+AkTjJhIpQIlkdyY/ei37iq9ghYjiu6GVljceGxbSzpB5vHwbvwA0sNR3E
QCP4dqoNWNJbKL5ZcjzmjHKGVowi9ozPalvlNoRZMiN5tkbd6a7pTWScnDUz9VPfurs1KMQBNYgA
RgEwqrDDehW7EMt2jSv5jDqP+DUgkwtvU3jmUj0SWsv7zaODmUeloiHgHoltQIJWL9tTLnU7uthe
eQCa+btNGWiQoEgbK1v+VWpWc1BOwJCL6YvBNiFinv8ZO0Hkl9MYEimtB9YXBU2Std42kynlA5Ef
MFJlq0cYHOn4M3zqfnIK/1zYL5C20SBH5HNNkyD8VFKi6pbMLLodJm33U6B/xMBLi1ekZ8JdMupn
vXaheuk5/rvASz8cpIYC0pBollcOEaeoJl3/pVm8lXAj4xq/eRTCYBnDbPj+GK88fNTacSu8pX54
oo14USxzavRrQ0uN6JbPs+uUGyDgmDMHVp512eC4GYayi14chOOkbEwkzUJAlbguxXWQjDfRewtI
UyXQk3nUeLps/idUQkXfGe1CAzPiEIUdwUOnmTjvQTU17LnuZuWKietV89RTotL0H1IMZJrIxsZC
ccWHMUmfpj5dRKnVkWeW/PbP5XQEMhfDB47cYaLWUZ8Imx9ake1iGLSiQdHaPv/Ek2X/74+yzoTV
0LURwVjTEdq6fPRmSX1mpmHPs93nYsoFujnj7N3j1m4QkkOjOhZrpwYUxDLndtOTzSKk6fHfb4jd
0dpmmMqghZqufhvZJudDvzCa0AVj1jamq+Vs4P7kAthjmw5WCBlLyn4qGhIOE2P9WaC1YbFfQN9D
3i1VuVVquKPmhPamdD4DEXwK6oSdcJ6L7TuhWo+yM6zV+eueeXkwLbMiAwQMFfYtWua552aoCJNs
xasM5goNQdaIx2J6YGeUx+Y1fLf2MfhdarZhy3TTLqcFEIGE+GOpcaHXVzjkEidkNJKASujYu7wR
azHwnbHm3c/igIfrOKg6TM7cxEko3wfiqE7NnG554aFu+OVyTOQ45iOqcRUNbfegLb53/qbZWmV2
ve0mzmoSpK3CmzvYg0uafrTvglKW0lXtL/1STegg6IflnvEIjRq+UNPwCPpqGobq8ZRK1XKawGWZ
8/bdWXWimzpaVAV89hPbKDTPZSlNhgCgBN++wf8iOOCcuKO7C7GficDsqsCrF+iYkwXB3HiLcpPL
wSr+2sZV++QAMQ+TzgDGD9C4QtjpTWqC8bAgGT6K0q1B5wcCbxiyFVRmn6q0QlVH9OVPQeyaGpkp
WBeLF3pl61eQXV4KSedOKoyLTodOklwc+uviWev02LbOMkkNk6tR2sIxAcm8bEthqvPJoMo/VI4B
BQFd+DnOlVaYnkaS4ba48TIgXIZD225cD4q66zyMxI1lrhtP3O0X/+QMdqZPywCkoYrv4BAeJg7p
OY4Zu3/sLntxZrApi7WYZ8eEMcxx2MkCoXeBqgxuLnoaQKg8sct1I3l7FupcmutSHNONkoywa4Pd
SSU7/Mwvl8Sg2MhgCEn+TvJ41+Z8D3TMx7ApLLf0n891iP3WNajjtFQbMwzRW19o2bxEtdsZsDIB
bvVisHHHYyFL7oT8i1VcRzC+7FnavHrIi72dZCyqRs1uGcejo+bXmJEJzZV/5sEjpQRFRlrD14Rf
uWZyhWmAugM+v6ZP/yJZXjCsmKNZnUxxbfsYn5Pk1l+8/qs03npGdXQdVXuGkK1ZeBojunmWnYy+
TzfncHzZr5vEhKJPfrM1nW1npl0Gc0Tl2U6uk04D52TcmRj+E3Yw87+1HuWtfmPO1v4EZQU87GTE
USEk4inOHSQfgUsS4ouIcLGwcJIATnXyz9rUV56TIVPUvxLY5k+Kph3aj7LqBmNjWex3VJ6/aPv0
UKJz1UGPQ8qYfvLIXye5cOvmkzXN0vKTVmZFVONwN6unfA+3lic6oFilwaS2gEfBxerFH7Q9LMYD
yVZsxMM6C1EwLCjvELRhBFJBYikhCED/kmWkQNeXRPIiiBYaf3ePWXOEsrQ7L2eE3aEYN8dSGPSs
claolgP58TBFUubdmY22DY0kpPLntEaE0Mn5d2SpgrP/Qs8AZH2JubccUa9IfYta6HuyAdMm6ypg
ByUe6kEA+DxvxF1zEQucdwbc8W+cyAgfCIhaSZfNAO6R4PPlrh9Q5UdYHOEnVG3vWodXkqLzLHWy
Ku0ZAmtJKBWAtzxdPdbNujBOzpYG7o4J0LIXTzG+vI3QhqJj1+L902/GOvt4b647CeskD/3vB0Ok
JCyQTaUcQ5S+exrqMRw8z5Bdu+VVd+AZeL/t9cgP2rMR04fDn8CkJ9xuOi6RehesXlLBUYHKsYDB
Ag2V4G3r4dD/LXZN7zSx75+MBzQTFQFJOXxcpl3P/S92AF/KGAh3hiRqN9syqPnXzsbcE22b3Bpc
nf8H2A4w1PZOaecNn4oFH9enzK4ESSBYgNxS+V2ZiHw13b0CunT10lXzeBEJTHTihsNHdw+64W9n
2ufnoKC47PdoSpb7tkN3wPadG+Qme1rt6Xy8Kbcg8CQYjmGp5II7TP9Zs61OZV1nhzZbjoqoFUiC
qDM2cSHKxigxg2h49N/Yl8iXHCB/hV+ZWGG/RjRbk3mAeDgAWUp1op3H99S595xzK53huvIZ8hFu
JdOFmEY7d8mESLoIsExFiTtduU6A/8pom09jtVao+HYNKLZCs6OXFygIELinOgx6syoXJzOn/3co
5oAHJE0qOVjFtpz9cWlH49UlsBqcQx8+pXWdTOK5e6ToFfntE+Qpt8SVqom/2CGuDCAEMDnaxCWA
nzady5hvd9rmPdIRqA4RWojfTbe6A2x+XbRlVvR5UH+ojVS4eXYd16TS5qZi09h0Urn2Spje/Cnd
F6Rk9ksx8TmxLC6qLervmT+jBoKZ+UqMsXvpaRADbfrT9vLARxOIa1vtiGdt7E4WGpjf9C7T+F7F
1npZPNaVKm1QzqdCfFhRBJjS1pgyNJ8kZFpkbb2fGBdVDODRNhkH3cqt+mWPkCvv+w8XKjc5NMJw
EOYYgw8ojnyXtJAO/uO9sT2T0yI50ScAK73scNEvBgt4pwc4HOIb7lvKQaGUkH4n1CgjCQa2bZXf
v48OahtEO3pdQVQ2j3LMKPj92lvCRppziCLMZh8em+U0j015NSSla648GgYVT+PFFukmkY/N7Lpq
yA2V900nyl6nv6Cw7uGsdvs2T22hrYQAs6CZuesMLLTDAox0dVk+n+7qmh+CpdD8xW2HlC6Pb6Uy
rpVs5JyNYHhOSa5Bf7agkY2bYnmIqE2iFd6S4ZzneCa6Sy7hLQ4pDlS4V4oaP5ip/uMgcnEQ9deb
Ii2+8kz0qKKCfOikRUGVplp/HVX2H5BCydE3Ja/bLIwh0HuWqNK9svKQ0WM41JedICZMumvNQ/E5
BEjd/800/ApzxQ1AbS+fPl3KiFzScE7QujcIh26uMDtJmTQoxcGH3RuXkd+qRVnPkEnxk6umwqkw
KJ902epLvixwk8tCKzFGFIFxOgIlzKiKxbWcTBFpZvVlDjBraeeSdvNkjMTfYi36XlhAcHTqd6ey
nTkT+3D5OGHa/m0+15HPpt+kGQIP3FFlpaw/eUowsjBQb/7Ovvp8TfTg+w3V5EgjjLgVWOboHwtJ
UkUgl9htxBS/BZKY2fp7LRp4lTENtutObR0J1pOBMkp/cHRolkyG7dHiD8iebrNPrxqCK5jIMgc6
y9i4lcUQBPTsd06/p2HpJua9cWH1BI2Nhe7g3ocmYQ2pvfle7zENmcqIcTjirmgkslNvWOnoGT4q
HPa1gJn9ZOFADiYd47ErLy2Lqatq5+gP/1uWwZSjIK4pZqWCi53SHCL0wvEY1DejWLJgGFpixAwL
/GPZLMCQJGiwiS7lmt6Pn5s3bE8yCcP60btLIZCCPVXdE/7n+3k3B1g0wOeLsjDag4TUh34KuMXc
TbooQ5A9TMSd/YyBRMBoey3ZzR8Hn57uSLXLDz9cUjZvNyeJ6A9iwVnTTEpV3K1lCxHiojBjD0HN
NcWw7jHIt+xjpsMVbRhA0pejzy1xKkakeh/bPLFRyBXULVAMTMToXxRs98DAh0ZvRN71J+X5YejE
Ij6plWCFIWRKKgQxvTwlsFGfLP+wc5tQmHTxxKNU1aNVNI+80XH/MrUuC2ByRwvA99+1h7POphFb
KR+4rCM6IxnZ6srXvml4X8PZDuRF8SaZY540GFUe948JUd0cns71dNCvXr5lSXhyLat9QshLsxUR
E0iDfLpKxO+axmNaLJzfrc0Vao05q7qUlILxb767VS3agJdrXGq3Edn8dwmsDLehZD/e7eoY/B0l
z5bNBzer9hDQ1JZXIayQkgYvaQGarmFnKkHN7Oy/YAfWASRfl2Ok1GBNsBtx9uUh0wu4Hg8IAd0r
4+QKMo8vMhXXiMtQL9nx5KnEXQO7TnuC3J8hzSpTZHwfBEJZpe/twp3YHVAksmI1bNXniH6u4DTP
vCEH+UH+XHxIPKJwHR/2Adqwpa7fYgbkqG2TIxom5LNGHgdO4vStJQX5PUcWUgF75TqlpL0iUYBi
knxl1S6CNULvbjTtG132JwROSFSSrrd9HlX3qsL9TH3t7+dujGXZtgVwk4LeOFCFz1Pw2wxp/eor
pSvq2Rtf30piofIgxN7txQ79hZEmH6xVz8uakiB+T9Zjzb/9dKtHZtwZ+ShjDVwUPBl4czJte98i
oM+dmmVqNp3fZHFYYxEYL78uvTJ/1No8m9w+wG6LTPEZawZMyNckZrZPSSifa65G0byD59yill3d
FpCweZm14i/fdINSIX+cI8lAK3oFTsaPGLyRGAaLPp7WS+eRSUVtSax7d34lwverCMnth18RQ1n8
fdEEhJx/KUbnRSndA4I7ACFnuxOzi9nQ5jM5DpSD3r+9yeYp2KC7euT0N3fwPUDXH8fjwm67dZAb
bB2wxFHdfHeWC1qX4OlsggxtXRyoijYSnGFwJgo3gbw0a/uQKAisW2+2a3kL03nlpp8jqocNG2n9
pNH0/2J2KlDY/Soq/UozNnPTRavcnr/ipQUY4lhWTIMGSARd3KLPRvVoMq8+wDk+xklKCduhJqlj
AIcm2JUBlbl8hfsFmactPzZMZiLZNIAt3WSRct50d3JUCFpN/JLlhMxYMQH2qBVQ8Gj8kvJ2bO5t
JpdGVzZDWOXEF9q4f8KTGYp9MJB2oIBc3bRzBQBTPtFWG/pjAmrshrP7lygk4zCkJtHhrGVMc6FP
tYHNCzn6a/mCdvi3kbnbBtCP9GhKZGVdU0jsmuqsWYmsHhJQiNFwT5C6idhwJkfTscfMQZ2Z3QAj
+1bDLHFzGUtLd9kfLn3t1v/ds8gBieakznCMUL9BY+K2od+UgdYz0i1/p0LWeTMctAYf5Q5Ie0yY
OVSHTylUX2zLuR2BRcBsGFST+LhBQFfmH+ljTT4i84ICFcsWhew3+AkkV1TRCjSU2iOHYWxNljNK
tB2g8WVph4HidVQ/FjTldwjYiOXd/n+EgI93jsLsRfUNDCjGXEPulwYRdiTMF+EKqHiHXqHdt2H4
zeZbpYTi3Wlp1K3h6iA5a8zVR6l5kEiQ1BXoJCZ4PhI2nyFk9UlnUpJ447KqqFYFGKSOQ90kRcJ3
AS4uAGBJNKYiSuU6sHcMUwMfoOUWzET0e3sdjEbGnNaZneikI6BTqtnIqF2LiQuNhun+aX+4+H+9
/5a3SsHdbL+BfBvecKRySdPCtz1oNzbiz0RZNuzh+3NsBMIrJ0wouE0A1pIReyFpzCCMBuAX9KaM
J4g498Fx1LseTaMe7pvc50dzDgNJ3Su6J95HKfP/aXwJcqVJm/1zLWP4dpoDEiB8goeKc6FnClgi
cT50epgw+I/dwiakDsJ2eolBYShz3P4PZopw4Xcw4m+Kk1G9H24Tcn78VWVQSPFXhoOhjRJUh4Fc
oSTMaij+mmKPXsxLT6t1hKOPPdF0Gnas1AuVq7hkazX89DjSI15xC+v4pwl7gR5SB9s8uiclHfLZ
UBVO9p3HpELzwMzP1dBlrh+cSlCkh3ueYt6uFbU0rkx1qEYH+0rgi4ZhMKElpZEiVbfthTo020QR
fZC2roJ3dqccX4bGe2TakOqlL9QP6zdQJ7Jm79vQhjHXVIS0p/Bp7r1t5hkrzUR3tfBMCi+3fT6s
oBTUU+yEQiabeI2vcaGBevj3vY9MhyH8G0vS5qQznX11exQzl0jCV6qVpi8TcGWGwiUMVlRdStKb
DfcZMwev77AUcVU7fA9vFgGtrW+grtPmBEPSYLBlNjNLzh8UVoPd8eR1Spv5XYFjT8PA0bCupCVw
D5hUQj371tNJrNtmuXQMcWaTeW7WzMdR4Zh+83ZUk3Uv8jH9doEedzoelUFNidddpn4ZNQPw46H6
m9GHIg0L8Vnm782FS/L7l8/2+3LCHmHjUJ5iGcKEKMMDhSogX0DWvUlnUKa6EV5CzzztrREaDR/n
VBE/eH5H18Crik/j2k2cQbftof+R1CDYJHi5VbTfLQmt79TLlsOssHTBKxXVwldoe0BI7PRw3b5d
wJUW1+X2lV850b8WjIboBO0ke+9vmMGhRJaJ6FfNtDkmOZnHIvhutPOae0IX1tfWX2Zu9/J9Ez+M
8AwvfjBAwWqBa3+g532q7Euzo8pP9Tqr8b6NvRdsQVJjmHgQrC+I4liLqcLN/cwX42Wo3anhAPLZ
3GMt/VqYPsXrnOS2BclHJLDXfIA7/h2PFieIfb/wbwfFKhYtfdaI9iSFS2Z9NDw6Znx+LK3rAzsK
SaAhspoM8srIwFzETGVOfnG1LkUc/xb2QG88g3QS4OMTyi61uOAnoYzq6D+G/xM2d6HfGshg97aA
bRAbRVlQgJAL1ugcmRHqLg4UkJKFnVbLCjpp8t3DuYjgReaF1Xy+DAXnxfgWXjuLha1MpkK5KDjK
zOK6ZsmMggOGZXA5m2x4WJJDmwiLdXheygFlpeeex5RaL9Z6rpO04th+Nj+MQAhzqp3HdPohTPh2
S2h28nNCdg/Lj6beWOmLgyNIaDmqrnNenGtgM+pIdBYaFjVzGtBATT02suMW7lGsKtUV4501Mq2M
5ctWlQ8lxOuW1BjsYRhdDclxxvardO4iz6tegEw6kfaVkYhZtjO5ilf4vE2JANHEQk8ZmiLASbh9
p1oaD39LQ4ph2OwjMvR4sY/FJe78v050KFwFDMwIxI6MakntczCfB+u0eRIUikx70VvXeaEhwnb/
wiA7zSUWxYNmU1m3E+SHO7HMmN97b807RDw/XXVBpMKwk1uS08L9x/s9wfUW50jmQeoA96wm7UD6
9qpJDStg2EWSDdnZ9Gxswf/1aXmw0kw5pBReslsVhR6H51sq7pstmd5GbnOM90uSw37IlnHntOof
IEx+Rzd7jKNZRW8UJn9dm0JYrQCxZQYGx5nH3tLKPa4Ho6kO6rMxAjG0q90OTBCoxKZ4Hbl2hZqx
VPoU5OzkzJpNY5wTlyJ2827kGK1g238QdjXU/+vniYCoYGH8DQcOcDbTI8Xsjy5eA4FOCZGvcSXA
9nZly9cUVTlw/4FHd0RXrJP08rTKH988Rd011DqDPAKSHTUw9BOFdhz8Nf05N5HnJL3GAoNfuAEk
WLKJjgjzudNHXi8WFHh1DAWB1gG2dCOPJj9dx3poWnHA2J6hFbRA2psUb4k8lVlgM4pAUX8GGkYL
j7C532Tmg7ovjY1R/mLjS20NhGH6/QF/58KCScoqhBjCJPofSwB0P8qw7QNOMszOVqPfDliwiH/4
lG5VQfaLDceimz7QrNgA3onRgTuK8a9cB4Gd8+ycNlkFuecegZ7NJPcO1/XENe6GNP1WNApoV25x
xGQty/b4mCEhs7AkNfH7JZW/y+WwhjGBtNEOIlBkxg4begFBNx/imaCXWUn/VeImq5DKjAsQHrPb
acmRkLe7biPZC/urUaYtfoSgvKJFelBEjZ9S5UTi+JaXyHKbfUdH2pdQIVxve9AjSEcIvvnBtMbT
NMM1KRrEZy12mD6AwGkLmIZkPrM45YWZO4RMhuZI9Bmr6BZUNt+vndnSSxwLT6TDUffI4o6bHd0m
8XfhWxL1m22QxXimERineirx6oP6Vu8XUBx2FKayKqIK1O012uX0xNTF57aEGLhRwVTsKxzIW4VA
jY6D5Th1sviJM3UdVh9yK0ttKEEP56J+OmTiO+bXHP9rZoj3WPbt9O4My8nCH4pMhfSdLKehtC72
0AtrmrpX0FLZBS2BWeCWAgxxzOLS0GnAZB81h6VEuWFpZ5Xsjz6MdnoUlFotwzu2XuB6KMBi5H7U
cwPwmY5AcdyPz/b6qMMCm8wtc818lL+lQ7DIlZ5W+E8xqHau+1til2TE1hCOYOp0lCUFmso+gwsC
e2K6bA46Em2VJbbb5lRfCrlvfft1d8EdhWUcU8xgfDAXIRx7HHbedMDsbYzbC6QHWgrMa3FoDAUN
ULYl3A5oVWAiXjSbNLCIWMZSe3HrvFC2FoDdjkYYwGtTVu0yfVnVbqjJyHI1aVIeQSu/J4vnEZ2m
cBVPiJW5vJIHDGygnF0VGTFzZKmy7OMB6KkLVg5U7OjRNxxraUQZB1ih0bG86a4yu117xQVIhMT6
snNebVNucIjF635nU6h3nSkB4pNvo9G3IbXvhO3c2cdWjpq6/UKfpV5sFnQ5UCCG7p/shH+ui/vJ
s5yzbPVRCOtZArcJgx5m21ESTCt0Wg+0KKrmkhb3LCqrtNTOnxbKsd+FR1n+3WKjW22Q262z6fYQ
0a/ZhFiB6r/lG8XqcclNsQIzvNqRG5bSxHE0iow63vAMeWxo8Rfpzy56N/j5gyX3vaWxOEqvski3
0jb1cSkxb4R6Uqo4/1XHuboF2M4MwFc4vf2477b4/L0sWWDzpGuxf94bwyho5JC84ySckUaik8h8
+rRe/p3j5R62oqnoOD5j1mFzuRQ81vRZ0WNYjMFy66SWhHHjRgFk9xvw6r9ELBT2cdYGibCzGsu/
BB6KFZ+PbM4tZva60PFNVifL3/lKhTJ+sP7Pg/0T5eKpbjHrV57oSboXTrzjimwxBgHBgLsF8ACj
Sls5w9k4iJI1TL+Cw0KpdoEc+Feu0t78B9dRxiHrrLt7zBS5ajK6bKH/UOvxtW/YtKoY4Bp888TC
nzXkQwb5wSvhU+R17tPNBoHKAHtQphyHQ9C4xHfmv2Z8kJCawZcmthPBc+FXpq8WYjNc74GbGTWA
hcmb+RUccwYfnc9qDNnV0sp7mMMhIkA3lJsGAtASGaA7CIvKrEN83UwJAwXSzINR1vOt9c0AAuNy
F8OCadhbwygXm5Vcy4kiyYITQWmbZv3pm1Wtg3yLdOzCgfba4276jU509Q8sWtFZQRhbbi2T2oio
/eHmpvFAfXeVIk9tIWFAFMigJTJ5C7t/ofYUyGldRooAH8MfQkurCqgjLAb1Z7BA4O3uMT+nYryo
b4oBLaGtbdvxilWkKD1muKw+2XeY/N4m9tGNCX0HEAOaAr/rJNHDCIoD7WL6DJXwRVLb253dFSi9
hUmwpERVAMBzZLYwbv0kpQ2IAg6veuE5RIgvN4yiw9Yn6xVx1ul0vYtBkYxynFgzfMlBwAOspKzP
LtiyWd/MTVHfou8/POeXa7KvOOeneSFJhiYiDfCw9zDdt55tdgluA6mV9+dXxt8S6Hu8534AaHBM
kt2TNYuvZsS7XlMawIqJ5nNL5d/0HlJjybaFFOquMArH8o4zhEP7htbuvaJMtqyMHPtV+2i0eCl5
QGlFy/WW9E+P/nHiR+TZ9iQF4rcUQKqBLILxv/zrAd6aF5JnVnd1WZpRsVPlz/XZSkjC+w/yEE/L
ro6ch76dyGkDIesMb4ziOyI6DpR9qb/OUXLz8Xp4isB5ePURFfz33G/d1l0AXivOaBvx/ltMrw4N
wupr2b92JKvUY5phmfgLw/HTrmUxtdgBPcaKAJFF/Sy9MjgN5qr1gPzC4NsYHewnAZ1eyj3jiGNZ
DfVx3TyNcMpQimr2/TfGoXmfQEU1FmyA+CuoaC2yKDb0hdN8OFqDgzlFJNSc2yQKLAPxpP5qOhlN
vjPKKwYOKVRVPGnmDnly+LuIOH9fy5RycOjSKcxIVhJSLcKBH6chtmquN7XN1WUmwowGKboMGm96
qxxCVrH7iB95cUXYq1C6BRuCoeTZEq7rRtH48PEdnlU4P1u+sS2SY6Wfkv8/aeJy80eIjrZA2x2E
NFdwR7bM0RLK8n0y0FvZK4xZQ1siYHHpQ3l21lcmNbodRh0N66qeqUrNaAUgrh2o1ZlYPT0VYA7k
HNBcZva/vYOF+EYny3kt+HMfWTQI8cbomfN3hVmB4PfuN0hVPFlZuSdsZPxGrGCzGmGJaD4wU30F
AJPJeNDaI5aW34uRZvkHQbi/JIJS6pEv+tEX1z9CUGeo0VmLhFa0HxoR/uUFg8p1JaUrXw98ybqH
qkFcIGz17xpZME34msw2mQRIxcX66EgrB6H4M7iXdqNbQLxMK97rx7vRtO6HekqauylyB7Uu8M8I
9bH5lJctAMyrgLFMFZvCiLwKN0rJsenEX4uQISP0GQt4O3UZ3Cki++RdP1AgxFdppoPpL/PN8YYp
azhYi2l0eLIDKRGc2dg11Z2THDJ3MRzHNguPdLCCEZaNtEiBzf44NNqnxOk3bBPGIfG3qtyX3w8H
dg2BKE2hkNgvSjGWoZW4lwKVo88h5GxvgQsNgD9+7QxgJZGNwFRqaBj/iBjztJvjPToqv/NfF3QC
KiwpmjT0ADBGLR+FH9FVepzU7HQFf+WfP3A3Q6icFMhrvL0Gp2OQmKWX9CLQKRXyTVQoJjyl4kz9
pBO+11mfWh3vgh9uFjaYSO0+YFQhNyh/mJLPRu9dUCxpGV52fo1U2VyDsPWFzca597PifvWilRWP
08e5ddXVTwIRRh3bfo4JL3TPZ52AXC3r6hBtL50Ks58FIiG4gKp0+41Sq/NajD/aaZSq650APkFA
O4GJ8Ydli81G6MkrkEaapbUEALyKt2lArYz53lNiT0TZ4GoQybv0nyIsOvTgcLSDiXkygLiXmmMS
JC1wWT5lmSUObdYY6yD4oPdX7EAtBIhbbzpzOi7qefBI0NzAF0VlKEjbW6lvjd4JG3AIhALFUC8Q
/paiSA437DA7/JoV5gYlw4yFUp1L4rU31LwPXmqqmi2Fhoj8o/yx3dPxjeyKzRtkhggYK9qwM8kk
ZRKzwX8gDtuF5Vc/Z6WbOVv68XCjwHX91/nCLRDLZQZ/EGgDhHGFaPxOURL6y9BAoi+0q8AzTKQ6
WiAq134NkOV/Vn6lw7NHKXhrw8fs8zBu5oCoyUv2rkX/Nwtk3y41Cz6U2kPSz0w33BukTmZoy+fR
nl3fTSAJ3lkrd3xJBOJ1N99dZEIeyIAOrisLrXhi7ykYVERychoVLAazMqA4wy1eKZyz+MWVn4yw
VSB7PqBvTHlZ4m7GcQglflpMsdwQA9bvNJ53HCO4jPj9BnJ5v3i5frRY8z4mAyVhdWbTrqP8qiAq
ysbDoVLVGnrJwDmnTRjjUdt4eqYBc/pLzgfy6Cvt2cfiX3cAK1bh8Ow30x/bRDHSpRwZb4U0X9NG
fRs24L0gldrYQXsSMaTOPEbOtuEMnZ9+fc6zRY8b6MflwZyVZKGX5FmTA4GPQj8FDCvYuCl6L3Fq
pLoxfwYDTB1oX4h97+ZzsdA3syCmp6fjcK8viAYFqlxk3GyxNUcJuDP5QELMtNowKcxWga2NzkOZ
tCYwOwumsVT+vLJaGuYb2uIC31DQD1yvaVUBYzESElUbQlGAeV/Y5pwi/Cu5bQTKl3AZ2j443jj0
SuPQUw3Obruk7ERHGDNx/tL3nPZfCaTWQuA1pQRX8Kqy1GEyW/dKcCEQFCs3UPcH0vmO8T+SuVZl
1qacpsE8pMbbcbud4F50yu45YXlJp3xCNyi2zxMZpyeIV7ZTjD1AtEfq6bdRt6TKuHEWyuEhUZJA
6uQO6enW4HUPYMgYywTFwILvCehnUgN82G1zGIdDDe6fmiRaLImhlbHWzXwaRBZu0+EPxcgIvdSt
GFg+eghhpYRf2wVmAh6g7UafxSJ8IdirMZWQ/MWMVqQTRrHmrg4riubux8MwNqh0oA/p/mvT5ujF
3c0eUY4vb9PodQ4qvKp+My49m1lr7ZE2as8Rb9ywkFqowk3TRV+8G9jY4MtVI145NdbO+ZpniUdO
/2Rp6ya/BsQVAA4kcO1ECgkOMky++BUVApaaXTW4Oi9mBs1t8UWf3VYe05UsPy1S5tKGKfE9p76M
SbBvrRSC53VF1XeWqKNpiNPZS8DUtJRfLvAAihIfPm0KBMLSnSiMpuXrGSN/ZEZoalZX9aT4uM3V
WbVCniJc04ClNWPY4YIr+cVWm7OMknDsUUa2IIdpvq63AeIzKTHXDFzkVYXkVCE1Mfqed4jFuN5z
bRtdKASc34ih6YqX87oLTpebvvrGGzw00I6HCtDagub2lZ2dHUuNdIp/xVOKvG67Wn3G/hR9ilcR
eo5zE1qoeGol4ZHzaHqesyPdQeVGgnw5JPIsMRCfxhuwaZBSORa7kfRopSAvNZKl/+w76AV5OWfM
PPeTHBzgt1b1FWQXcB9T5TW73lx3qfl9IxWc8zTokstbDtR6Q/m8JHBPzr3S2p6AODPYClCoq8Cz
28yq9i/RT9Virr0YO8jvcPhq9ZOy757C9NEfbY/ufkr2QT6biLAqXnKXfE1JzUxAIcYRkEQfOTOh
HsGpjPjQUJqZtp62Ljr9zsOhC14DbydkaN8VS6uQ92mxiQbNgoVnhGeB6cwdt2DcLSetnJGxMMAd
B6KIyVG9sQiYroAJX3IbVdM+1BtGNYVIZEJRfrvB7S5JlMs5uFDdQTqIbLB+R+cHb+ybAHrA/gPx
wFtMPVtpcAPwmKBeLenUlA/bLl4tyJLJ2iD7Xg+3tjiEVgv6dTO+nxSyX3VtVoWUPfVVXd+EWaLz
1Yq5XiMHGls5t7EHtsEDdohq13VWnwqM5MMnV2i96vE3PWmpw4WSpGb1eSmBm5HSrwTOZBADJeXf
eU8fvp9TazLpf76myHpstZ4ToW5TnYLV08JGgTR/AbNdF+d+tZp4alkNCWFI94AxQJVrr74VOkob
LysaYse2JhAXsSyELb6mEeb+XvoE0r2+foegrZPnj4rwi64nfC9IEjfsG2tWbrd1G4cikCjEuTx1
mfwhHC11Cpkmvcg7enIDg+CMcWjjShM7VyauAPyR/Oio+gUUOQR30tXGhWC/ymhmKK5iJeRWIe2S
JercyXuqRNeMt780U/niQXI6K/s4cZauR+eFnYbOkgwZR41hXdbTNErwd75UMculfbjPX0WjwZRu
r/Z6UW15WIo/9VMZEoreObBzm+acSsPsESSf2h4b+nDa3l/qvhUIIva7JFyk1xSIiv6MRpegEigy
K7mB3xJFW06DmrS1YNEf0Yhozw+N6MOQqLdvM06I78tEncw9CJpXJ+hA5WtYEurtSl1OZpdRjxp4
xGThYgpMdUCoibEl6cTF3B1ROSbhaof9qtUYaYlsgsP2K7E4yJGTrNL+9UOC3cqbK53FCpOqyt05
qjksrcUT11ouO3Y//lOxHEPFbba6Mmcbk10JdLnhyIZtm+zWBU7DMGGT82kaPZgkaHUqjbrO5dVT
1j1haKPYiCx5h9e19R7Z2RvQI3qnIs9f+848sytFfITa1u6kqWCtQSgVzdN3LUgnEevpdcAxlBf9
/dtXAwwRjuJUJdjifL4Lp5aR3X/UIfJwd26Vp2spi7IPvaxqXxvNH6aEW7y6Bxf/OWYsvqhqOdnA
mMeaFqSODNl9UimPZ1IppkwB4Dwk73G01UWvebyK1h/gfbclITVl/s0+hy75pdran7ytAsJ2KQ3A
C35FxnAX0f3zk0wBnNrE/PDLtL7/owmeUqoNiSNsZ0NE6unXbpKppv/fH+zzKpYtH6vFZZ/Xa7cN
crcRKJ4hLJWUKMuDkosrWXeh3/WlfacUjzVN5lfbvfu10jYwabaXwr7fmgO4TcJfTeES5ENCu86P
ZmsRdbd4LtHeu25it3VOdmtiuochth0MrbfdbbAanGxJqJiRF76re6kMTw3u+fF8VOfPX5qSLs+p
7UhBnLIvzcz1KCYvT5BCMTsmhyku2GwvivtK6tN/fOxVUQfEZhQuhSF5WFDmmrYQsOMm7t4hJR6Y
K5bKxkAc5TtYKFs/RlOzfqbqBUmoCcEiC3e9yflIEeNhZVfY2+3+vFI7K/jBwalyCRvvYPACSY+l
dfJCevSKW/KCZo+tHM3Av15x7ArVOYriZ69BQ0EZYnypFjutHwLBUYi5ZB5khkaovZl+tCLCyLZa
PIhGLkRKj2mhlUVHGsccSd4gASHlfDTrAc6cgrr0rWz/8TgnqCJtz50eb6ZAYqoCoywyz8X82heG
kuYMj9KYcamgibojBYUNh1ENXWo6oreYlYcBBZbplnB25mX4EBDOu79UzeKpPLoW/wBwb6SIFfIB
INxnf34lKpTpEHp3KzXXXecM3fqYBWP9RRrbyPkZO1AhwBGJ22CzHsL+PNoqAuvNGehv+jAf8lyF
RUD4RfJU/LMBWMYXQRuHtWJ4TXfIxNu4YQ0gZalcfQVrB4oKtjVJ0GLmPtNAE1yo9jJuyi+KUyfr
/9zKNkw1IS+70asVS8EI9tqNGLPy1EYu45LGjQGDdQAfBU0ARdMR8NWsT5AbwzhgV4N6/YMS1fRR
aSIFxcH1o3/Ex1BD0S64xLVJyraWVyWe04RulJDUR/kJtpBjN4W090Hu5iVB8ZLO7u9TRLyxR9DM
zIURh/Bq6jV3bb8+xeP8oy1Zw3ZIWWBv41wEzIEcMaNZQuIX15kP9lZ6cgQRYTsGp4pbm8+TrrmN
q5SWGfeTxlWAIJwsW2f8fpxamqJLp9KRUXiTbwZwf1yxBhJMHBIWL0c4jiHlRur5ZTuaWouMM92Q
XqSxIE0MKbebzBg1ObzAPyEtNqSWGAQM69VUDnp1lrf4oKDtoGr1JzarCfP++W4zMghCgP/v2ESu
laW2i5EFdPgYMNKONoU2hrMSYc01F0iRPrL0JKFShdRZrNj0XsMQ+M4Q+GVQkn6/dDCNpSrOUr9+
UrOgd8/zWaOSpF9VPY5+jj+g8XSqpgaRRB+QijuXofWE/5KjynwkJYcq/wz547mtroNNVtPSaonZ
QEHoepha9jsT+TPBfK6oqgEK6a6K5b1dsOUvsTENL2ECXBk6vhT/QVeaDjGkGZURXZI3djwg6LI5
68DHbpXgY7yNc+beW555VVolkwno5XNLTkv/+py/e/y0zdkokPsb574DmeDMiGymQEb0QqpkF4Qk
OvvQoC6hyS7goTQ4/m5pLLkZrJ7M8in61N40aBiJsH1OS5SsqKFF2v9c59nRdujh1w46X9H5ZGpH
ont1PtvqxHbtPtlCPLeJilb4fNfygPjTjCHaPgkw+bRecxYNztMN4HDQOjwNLg9bVNi1HSpqN6jF
rBQYQ/CLtqIAEZ5W05QEjhoEkPJ02gNYUWEUq25OXwsEgdctA+fwhbdS+LvzBzXfwAAwI29NEWOO
JeQfUaNUwyh3XORodY70SbfgulGF2uHM3TqwWl56enh+yhvRt9oDr4x1KND31qG2J9TWT0DZ8JEV
9J4QbmP+FJKt6bhwNdK+JsjyKE5uD7lwh3cSbGd5AhZq2r84wvpS1ylE0vI5bfqrk+mqXt8b1byd
VEdvO7s8b+a9istw+JM8s/86l+71wiSMCYLdHQ0+rZhrz9ZWxihF5vPhOE71vfY6hOkFmg1YLF2s
KqoZkFIuQU/E9yMSa00RdkP6hDr1RA2RXB567ex2kZQ0pp6s7uT00H9/3RKglpu+r2QtZRU9ZXxY
aqYvoAuKGSSRMANlN9bsjV4wW/LTDc+RWljPqAUeO7a1y/QwaKKxu/C5Y3PpTV5LGjfH4H/8eUyn
NgKIeq0i7VL7A2sGdR8+ZlnZYpM19gAFotaHu9Dkphxz87MYWRIiNkpjFXZ+XRzHwD8bFEGnhuXD
92slH3Ndct7hBNBufTA74CQk2jk8dbwx7uPcaPFEyi0UhUYGHG0N5YFu1AR2WCLXKXmi1XEG7COh
LfMYT6eEmUBhmvYz1Hn25Lmf5nxMu9lD2ZJ4JpIECtS/5CWqVjEc5j1zSw6s99SEL7g4RZDXOsXA
dh2FNi3EPzFR9PO94JZfH64sxMYJO7p34qUL6jkZev59uKQdHTNV6xD8hpmYyqw5IucPW8Bp1hvh
HuPj4g1GHxE7TE7abRiieJ5hXKCZhtSfCKs9zJHNJCjs1BbQMEX5Xs3nMRCDUTTY7uDBPSB5HMiw
UIuCzw1dQQ4NanwT+NiCPOtu0SpTqPwx7vVXCfO98pc3Ux1pPxCFUDqPwpRAanGChnEThCdpEcfl
5bA4HOfzF/A8PKtzL+XKFaeHy9uQLaGp3AXvRPvly8uqLzPyDD4gbLRKmIacMp4Rvtbtd3dAi3UK
zdlyxoRvywHjPaenjeyUmz+3hFxZLIslco5FsPqh1XzZ0ppVMkxJ6XlgSIMTiTyiK5DZiIuXiPms
/LdZYo6gqYG4kr8M7RP8Gvhoe9gsRu4wpvpami81vyi5y0RjRkiAmAiDbNYFhKwddgcFMwt9nZUH
e13ok3RsGKMNGNgJrGuS0n3+XO1K81e0QQxtzdlMJCng1OKh2j11zRsa5r7+nR2MCP1RmCMoqyjs
6NtxD0p66nz8WjwyVLlRZl8XjTglsMK9hd1NAFBsfRvgBv+aUJX546tcVOLr+RP43GZjRhL27NbR
DO1egpEoLzDvmVvDac09eZ/l9UCWSwDIk1Ms2bIxnWLXFX2Z0bnGaYx8hC1DDSgqegukOBRxkppX
OirymvynsYD7zeRv9ipH0SCBPswzisirOYfKVMCLyQGN3eFTo7kjnnr7ZN6wPQqBAgogF/2pm2Nw
H+gg3W7Jcm9gEfBheBKl/lL4XVxL1hPaErYOSENys++r7MZ+a7oZ7vjXPCmkx/71Sxy4Om3xuX7+
h1Z3lV5Jtm/HLNy92ciYFi3bPTbdZMzdDxRG75ma+LMCFDOe9NyFsV12qReFIm+y3J+oa3leGr20
8Jjiv0/DeNn1H2mFopbUFspYuA7SJFj4r0HidAnLZeP8ish7ZtHEDQQhZ3VyYk05swEhy94i/WgE
YRjzcXzwtX10B4wMcN/kLCbeAaFjvBXDp/Z/fildMl5F6RPOWD5kzVbaYnEYWDk/O5YWGhwubyql
xHCDpQnbJYnn+8FjI6WyR8aaz4lusyAQxa9sjOjHU1D4MF+ulR5BHMIZ2kunaWFjjpuT0o1nJMuB
6JcZaHzBccnANIstW8vkEAVJFUnMnw7OcqUhbGVxbxlBTygH+uIpXI17KJKpXfwMgTYbNX/8WnMj
poyBah9f3TKG+Eno72HGqTgDODvS80ckQZRum6SJoas8nH3nHNNuQRZGUPi1NLr1XpJdON3yH//4
rXAwdMB82d1vyjXRrv2HM7kuDPEdi4j6yHT5DV6LQQu3D1VC//8zpa0mGa6cvnmkHceY0eODMHoV
uIJCA0V7XCPNnBxlLQoFkJxVwLvys+cyby5F3bFZyYNBM+aMyWeKNTEdM5Fp6TeUhh8BqmLYULbo
UY1HXcpc6oIJUGxlR/Zs6EDgEpes3yhBsqfsjWaDW+K4CG4EI6v1awZEQMG9TbltCudtuCar0ole
EmVljlIqs1scTKzKH8+RehoaVDORSmebCm8nZqBjKJqFsIjnVXpVW3S3GUB6Ts+/TbNQ9SMsgBoE
6Zdg4R/VqgN2yGqo4qe+vNtUvCpJBX3kBnJn1hoTe3bmR7/7FDXpH5jnNjaY3de0nv30o4rhhk7r
GkAbNf4AJMTrpOf+/gjgcA4CKh6to92sq/ZkBz4u7q1lVsFCHfp8gSHkFEesjIE16dpXYahznCZP
C8LxJahExg7AwvDt1Ob8MiHjBZTCaxF6C2pD2/WVHtIkekyx4bG7bUzLrtH1Q8aWzxovVjSqcE8p
n0zicoLsaZNt8kPklx8Yk2Ay6kFOLTt9sIhEzyojoR4y5HVeCZ5y2i2Oni7GiagoCKG9Gxy2n5sh
Hp6c+l/uj17eYQWCfezmojiwwdk4tGdr8IqWTXUUGfy25/E/5v9871YQBjzQ4qt0OM31jEO+AWML
neBPlPWe1qmCF6pJX4iMUXYFVXera1vwScXP48wpNcWa2QZa+uC/bIIbATsU7YaZMYV3BmQYXuwT
XqdBoLDp+hqwpLPc1xFcftFRKiwRZ16M7BwsLlX2hwQvbijDw/Qr2ddQxrzUE2RQgAxDpePxPF54
02mwkcV22ZT12Vv57QX/+fz21+WXo9hoKyTdhS2WUoZ7bRQvTwl1vLWBF1O2jQLs89p9DhXp+yDb
g6f5FVGARfYGgiEjiWZed2DEG/ABCM6Z8BkVzUlkmjq97TSJUczM9/ixVztLAbeLIOr+g2i2ggV9
gwsjTNxe6WlqGl35fdQZbgyqrZzPRnIIF2PIpqPQcVCs6lp0zfq6AKsRB67alL4jSSSp2A9ceaAN
KODGLTBZRgdNL5zOqpthKUxbuuAeNHNNdXdZm3L/mPlzoBI/AflpMlRn0R9mD3xaAMw2/tN/iwtA
6uVflu36I+9MsDhQP9H+ah5uG46u+8WD6+POI+wlhnLU15U7ZaHfztt7kffHB3SpZn+GlvkPEXNr
xnYKZhkpcGTVOrZWJUfdADpIpL4E5t1pMBpBLP5H2ozyCs0OfBIsTl3oZZAnvAxLgZTiBTp/k4cc
bz/C0LaX+vg2IrE0fMUvoy/Q0Lr4G6ChpVsBgEShIGc3fPDJ2WamTLZPBivluMLymg9t1VINaDpq
61yGukFVLSfQU2IuWuxcCkUIcD2fdX1A+mV8f1tDfTaqS8by634uuBA8ZTuuhRSJiJ1DR89OQxh0
0m/S5bygABN9SxXKCaz1m7+jfy4mrTMKnJJyw1/vsCzftkiLcu7F6YDcbmUBjwS3CxPOqacAcnDj
iwnu3OgZrioCYcOXl7ZMPQHKBkw8RpbV9V5gqWcPiaY6DtKO7KBJrtNEzzFXkqkVLecSpV6dwcal
MPtiqd9F5qxVVvvB9iCOwkloBsKA9qTunMN690hE+MckpY0JjmBoTgS9h7s6kP79uY9EC20LObwd
nD4FjAvWbgtRhXlyt94ljiSUGquVOUoZjwMZ5zKCdF8k3IoKh324gLaKqIegxR2kkNv/Y0+LRQp4
EsfKbT5UmbuuEO1VTSuAVOLsqejdqsDOT+QUv92UGK6Q7HcE6CVkrs0vmGKuyIqDqx43+i2poeeD
5j6Q0QK6eIyD0bIoT6/Wg14nqZ2u3YE45c1l7hAFl5Aqv/RuL/VAQYAp08UPbFpv4vW3Jv/iCKPg
syxywmhpMCLjWL/l6grj/P+YOh63cRaOPjWIU17RgfHg/xg7m0DvMOYwmc8zzavGtytqU9dM3l9Z
OXX4raa0xtaa42N7sA27wJpfiK1OXx3egHunQihRRn5KRwCI5AWBwb9S7Fpp+Rt4HL+qOgZM7vtR
iYME3gHvN3VzF1IWHXn+EpdEWLbNnKC3/iPxlVKUuLptzLjXnEXWariA112g7qMWejz+S2P8FWxu
zknBsDWGIpZWZbYnVeXysxqxTK3odK0R6mLQjnv9Tb7L9d8trP0UzGAmEr5sIRvWJcn7kkDTMfE7
khCvR+kSReMQTS/Y1/m71+LIAZQJH+Nlzt6FjYiCwlXwzeTBF8rSqdWouqBRbxZ/9vs4DCqZkWri
kpMH6jv8zZ0VpZk7glVRf6qRp8bJclIzwjUQ5sCBnrv47mQHjTyYjuoH0ZqkxhTbnKt6AWHR6fV3
PPy8h+M0eodey0l5yZLwUfZzAZ2BtjS56YWrnCgIu3qtt/zDsK6hmp3F8vHaqBgR9EJwVtOxDAec
T4gt4C/Z4DB0gTG+3UjxksL2IPPapoStiNb0hsuybW/dHKpr7mS8irPfNKik6xnuaH1LXfwrKNUI
v7p/m/x9jhHHvdU7+EFpzskpdl4JtFoAJ7mPgFUbT4S0bIAbWq2z+VMHJQxOkAGdVHMyYHwDLFqr
AM82MU6292jz2CtnkvkI0NEbjIvGGQ9r3uaNmbsybm6dZianwSnzh5xStnL7hXm4oskUGdVMbLR6
w1dpciaIqxqa23ul4HPRr5lFhSppqAsyUJJHmXp6QYhXNWLJVpAKpKWudJjxoJ1rXMQ5ZBKwTTpo
l8PTLoYco4QWE22v4koUVU4KQGsffr6c0wUvhlmTQRBmuRXcDY3l88sDU2wYeY5wjOeM5eqTRp12
2TrMYjRPSObqxKSP/7JWdKS/8q51uXhOn9plVWQJbQcXIXW9kmxDNlmTB+1hhf+JylyxTJW0ChsC
AsAF5STcdH85aZKCG6wRf4qM2TG5+5VkKqIC6sryLMV/aHcrRF0at14zZK1qOFlv+QteCcryixNu
/zmC862G+cKRYta7M9wvGTsnLjKIfKj/0kklnoV1jxBi1zx02gHOPQk5FUVFCwWW+YYaRMwCn2BE
furlqajRyoh8D7M2e9HRpuL5zQg67RYyyGb9YLq3athdugEmdoElsNKZJmdjHQdYJWmyZF37Kgsg
ylaubWLrUKWft9i0hd/0quOmKz2fwZtwsDYsRTSUCV2L1EdyIKooxLLRUYwBOVhVIhX68GXTyAOh
5u7fajhvgaj2DItkeJsqtcWvP+C4z8wuPOIISt60m8SWFQIlAmHEBc7s4QrgiLtVxR2JT5xaaGcG
JEEBMYQRlS3ql1WaOwZ2xtyrwYwJqmdF9HltnjTrXKnY4olsJzCOoC3PjbCpdaWeysLv0ymhVAcU
XierwFSgmJYpxjG/SNkos8LMN8ubFlXHylBN8JWaL7SGLh2VD+cFkEymZKH7ibEFZgrkkwP3+mZ3
PiOjtCw5sebJ1vf05WzpTW88ustzxptt6YN/biJKo6aRgylkPlELAYq3ffATrcL/PEP4W76IoSGX
rHOoe4aWrjAjlmgjOaqhPS3CJtF7V86QqM2mXxiafNOCMPg6dktRA0Uu50SlR68mVQyzKRTui2lj
EPj53yt68+ER9o6IWwEs82R3I7Oy1zVxJVGuH8MCoLXrfpMptXD/+GTlvE4SCAu841AGeugCz8+F
RU5qcuFxoejBbe12SPjPZ3WNtlmBLTy3HD+HsrVuxLFq1aTTj/SvUHGHJAXOJuY5CnovHp/tEXDR
Wfe0/K1opOnkfz9O99EzPpHEnuJXsloonwy32nh8d/E4BD2+X5kJKfu6IxNPZV+ZjuYip9meA/VF
TjCzkUHRduHnpcJlkwR+sTf8FjYPjkhTtls00EX3Q34VPEIRLMfWrVPtPwFqOF2cGwzvRUlcj92P
hThlqlUDjYMWrgVYBbOtVfASxJ2NUQdx/pvIwMY+UQMIM0t1eYZKpMjONAwowSaNZg3nQTkyYfxU
qgXBluxKVcs2HUOBNmVY96waHz8e3FW+fI92NR1AARrwiSkzIZqgPLkdH77wCkVZbV3Yj0YdTy9b
y+N1IpWgOgZzlgQZj2KOtORKRJCAmKknEyLZt/F3eGtZ9HqoIY0zLDTOHBFEQvjJ/oaMgACzJtfW
23RqLRqwMIuCgIuiuav0yIOFhTulmLYKCsOBJR39/fChlSKsD+HkFr5LdyJggnQ3U9avQDmSdBwi
kDYL/vCQFJHaryxQ08WegkHgg81QhgU4rdrfGv61uJtuk9xcRNfHb2AbYsmwtxQKg8EjLhB0UPZC
29IVeZaCg4d3fXV6vWfywwmtgIm5tgURO5HUjKnYSOoo4F6bF89p6l2tYgoVv68/NihLH6t51f+d
ZeNxiGU75rwgeQUivjIxxQDBEa5ea3nI6BhupT6IdibolAcH6LFDjl6k7psiaR2fZvwaGdnEfvSM
grXLxEBWDADAZ+YTlEWOJVBY346fiE2taRxpqTWPMa7fR/bUK3sRvFvSY3jpr3/VBnXoDXj48X9L
BZ9mgsnV83tVrt1+E5mAUP5a0OfTdRyN8xmEk9Symll33LaaGI4PIe6E8hAda94GC1Ok6VyCbY7L
fZasCMiTIrNju4qqKNEXqgBV/Fow9Z6Z8QKMgPxo1IVLu7J1EM7/Fqg75xlLzi/vir8Lg4Nx/1Zy
jcf3N/sOCEhatxB7YwHQ/TVUt+6uNbZ22PW35YyjMrOzyqmtkBjNBHIwQx2E8PF+V9Qf/fHETeao
53EsDkdQaxk2EkUSNwbhGKuA9cwjYezMLc/R5ywj1anm22z5BFuKmUd8QrNqXVM3moRKHLqez5Nk
/bNuE/u3sGi+z2PI2SSu5K0s0b6Q1bp35miML8NtP6Y4FCH3C1REITK8iTJjbbaLqC64YkoUyCue
hLFd0udXYGRZad1XWM+bIYeL0Z50wnZB9I02M6xSJxpDSHNbsPLiUFWNToe80LAPWfOK5z7wAtuE
YK/sN/aJ75USexKuPvj7/hBMn3CdgKMPzajs9Ubo4u96hR7fnMndxQUKpkP5dtvAAnOd0rkVUvDC
aSu/1g/7fpN+aqf6Hp5tC72iBRiR75AwXkbUTd7Nia37ucFli5POFI079QAs/USdbB2LcMVh6QCp
L1jNEIJ81G8xck++0/DsQYiojPo4dY654YrS73I0sdSMv/HRcSQrnTdr/rl+zXNVeelassrstYa7
Sg/3cGBsdkcqj7EFTfv33iMgWvfvpTENbf3tnz+pyUYFiut4PyqIaP/Lb4h2HAebHQ7JnaeZ89PQ
dqIYZ9h6osFtPYmvKEFIUYwR5VhBQHAN+N514Nd4vZzICHd/kVai7P6moAQptdRfgq9vRmLKZDEP
/T5u9Fofp+eJAlKqsMKycQE7tmBAFfuAqT+GrlxLEk88DR4Q/KqJd2pOOhTpkQivxcgRMNboRlbA
FZcw0orr1k2/xdsD9OQO3bV7K0Ef/jrnyvQGlWFbZg6ZqdGQGhiM+iKDWrDCXzMT37ZmR/HAf+Ud
AznBjWQBZn6BtOes87i2hyW/B1jN7pRd305r0AVwkc5qX78Bmh2mIJ2ZBZpedmfNC51KPxxWt6QJ
GL1Uv/5QapKjD0OV+do6JKyEOrOM5PODNl6N0hY7rouFrswkzwikpcngKWorQGJ/78MXIVTI02co
V2p0ocYcB+J8Ql9R3SHCFlEMTTQV4F4/61FkpEjkAOpWTS7tbm9WLduOel6F2mpopl4ae03Tv4ma
W2R3UVaMNO2ojpE1WPuFiYA5XERPIHqnLYg5ML+uc6gDMDOIaKxXa6F4xb+Y3ry8y5G3ZHkx+5k6
/rfogQi3IkA6BDg9i8YMUJM7Bla/rafS1hw7XwEW00+QIz/smpHuvukYP3RdXMWFd43cYG3mqQHu
KvL8nGhcR+HXDiGbjcyXEIihf2FM7TLGsXh9qRKl3SBSHEKH6UXMQXNeGSeJLUTBuIQqIDGsXGCa
76fVl3nWChECmtGlD+Pf5SNiHYzG6HUgF/MI0zBYyglILI7r2Z2oDoLfgHF9dLZI3kJENzCgyONe
IvYZ98DkgrYgpqdHUFsU1/96c4ywgmFcKEWf8LK33KKUWJGmV/si2+7rRt9OQxBji6OHa9jLMQkW
DB8LYCV43UcKlKQlEBLFTTUaDeD7KPflkp+7NC7f52SLLd7ru+wxH5jGXkhodicHvT9xjlMixxUH
w3BbDLAgPGWpiN/59A4p3UvmsNV//8iP/pKOs3dkW23wLVVgNMreCsi6c6IgmAfQA7qHrofAkIzN
47NmTQ5Ilq++VXawBFGRUfvxnfVBkUEBJrWpQgjszedDJ/S1n45L5eyiCCOeMNCAjHkd/wZV0O8f
UhuM5wneBB+m5NfbjHthZq12QJi/0xNHaHUsEZ24frU3QH8gyFezB3AXdn5qHUTs18Es2Sby820M
j82ZAqpPSB5ymUtxGKzWmmTQ04SPk4Knj3TaXms6XBkb8aTyjWgFQBGOKT86vmqXwdy7ewilg2gK
1P31lwIQGW3nATJCA2SYKvAUYIka9zU+lxPzFyQjQJ+fYWs3zt2aGT0F1as5VfikldDPUckyuoOi
MOB/9zCTIEC1olJ+oEn0kETTPtcgB2+AKQjcLM71RbqBwAvsFPpVMcfJTuuvU4vQIGt8bYGdEAaD
TKt9/F37VD+AeWypweLLGFLWeiCBCpUg51trsZXm+/BFT66Q4eCHQXAJWQnMO9MPInaqBJY0dNMV
NC2lFu/omVDjQCrQxzpXJg/WNWEHQjrA1CohOyWY5FXI+orinpX4kiVQQeQG1WVQQDeHLrave7sl
Lg/bwwuwrWUG9i6tfEF0T6laSdfW51VFKyCzwMHOS+QayGSpxvT7pMS9CQcD41Vnrlz/S4X0KrZN
jsuad4Bb5fd7Lb/8PWdDfCHaltJ0N6si9wfyQIML4z4PX2VL7Dr47c7xP573j/Tz7nuenJW1NnuO
qP7o8cTcRknuBfRT1l6R5h2ExjFblHaYtNsrFY6zO44rbADi070JRn28WQ1FhCv9c1qJk/XZzxYM
0zShb12LFX6vuB96cMiL1LQVVyHrDv8Oqg7xUHXIYjun7Z5ilNAR/2jaVsE0ICoV49ewaVwnkVQM
lCxa6of0ocIvrYQGEYMAkSCJKSNulhC7W/sIvYu5nRNW5vztncEJsViLKqPpitIMP1Q4ycMVwWsC
vmWzlwuzM1i2dTRncZiA+HktazN0xjH6b/xs0lUBYD/pofwDC4YUFXNscyw896B/xh0eZLoJwoH7
AEwjs79shC6Q4BmFTs6oARoMli7NL37qKfzM/8N1zYd+eKABMMku2CLCM9wG+q2NMPyjtP8RIEgJ
i2AS2Iw+Esm3gJxuAzoNvEQ1Ifvll2GhT6PmXPr3uKqdPJ0onaow/tiXBXLJH37Wp8jhU4wJS1ib
TAV7ShXOS5FY7EHKR9NnqxSZCnlwXTpRX91m5iALTAwnUi7a4apts97fnJQno9GkPNV/g+SbyUBv
ttx1AjjzuM671QXzCKQoz8EjYgDdPH2AVxuP7NpCAmWOnT+FRi2eUZJMwVXHmGcbQWKxmmEWdxaL
SELKssqeV7i2M3BYQ06Qd+aEVbTNxxPzgFqV7nchGYnbWTuQXyhYUVW7bB7XN0jtkff9wJQcyX/D
QljcdLxGS/W9xzMpQMLhB04a6P/HZW3IAWFPIskgtrXAciviqVluOXsCER8cshTDuDJctNNlcdk0
DwdHC9sqf6RMIPVcyZi0ImaTN5jn9IXU0bdDWoISOHENBzUNyF7QrxM9sWMwwOerRvF7bqRjZYVZ
zWRUTeXskwCJFOv7ypNds3fDNc9XJKHmhTS6cesJylocoF7in100daHx8CW3GPFJLqKIpTm4V2IV
qKJvAvv7RkDPR22FB04bSqK3xfaWf3GAr6Ux8H140xgo0Ublgag8uhVbImVzGj5WEszexQA81FIa
rldCVT7cv7v/RuZRFdYqYOu/oIF5XrYFiwZpc7iHgnJEnb/rbblG9Wv/ve283pBfbrpTuLtpGmrM
0acBmIxKop3wXNwaaocdk6LtEF1+1rueGl6i81w2Vi496H8IhoHWP1FxK1mrs/0BNEtZCusb+A2+
32DUTB7s+g+/I8b4DUVetPTu7WvVRTABhaEARoyyxt5LidHZEVPndSh1bdR3BRzpMuLsZm3xJ2Qn
i+9x5vrrSwAUobKeNYyt9e8XU8SrrjgS09FYZy6lqFm0iSBZv9VAUHDGI9n2oyYXxfbEH+GAZaRE
KgmZGzX8ZvMXBGTIsXUDe1SatgS6yQSmooukK3bZrGLYmJBbsu9f53hhACme2HB8DEtLdQHgzgrY
5xoTMsrMeyOY35Td6vsxKSog/4Kbumz/o6raNF/Fha59aR0pA5NMszSZN5CpYmjITgEul+sFtY1U
aLuhx317zaZxj1jy4wJ2Oqszj5xvZaxf2n6dNQE593+xENVoKfjEVJCxgCrithsVVwSWFkyXDYEP
wUc7UyOITqGI+TscnXBwAM5CAfE4rMLZDIfuXuJmL/eCoDRdwSqWRfD1xPk6EYeT4JXLrlE9Egu1
c7Sat1y7thSePtL5QhsE7Kt87TEVF7app4r8wSvjw3cSHnXM2mro5olo7hstnhVRpmQslvsOZcQL
EuxVGExQqmWjMoTH3BZHt8JJ0Rar7qCgXHh+k9q+aLiIUxyEOAoozB+FM2eFgAcQhzuUeHfmyOqE
sdS2wFpHFvTbGWTyvX2nojN+C3GIIwqzTbYTIdKFWTqDM39H2H32hJYIFWmK3OoMHbXzEIeiFyyB
EPZ9NEJVJmlfArlGINvmbkePTu6du6Xoofmf/dlILK7nbMxVTNjFN5He7KqckPRcoFcFr2JG32tU
3wdchuMOgOjBECv/cedLMTWxTtc315IIDi0piTKnwvYNB7U/QfrVqVZYERaRPRQTVAYe9Rjcb1Vk
QvKze2fMEokYRi/OepNaAedlvss/TyqwZ7Lp1FzdcMNlh8s5Y0FXt6Brm7ApK830+Sd8/8wrMQAs
kmr4hVh1y5vOm2EAFumliLRxBmuso5JXwyEG35lkDnFOPr/ATxUX+xdtxH08MYHHyMY4b81qBkPU
DLOVTBobHs/HTe4hukmadsGkVzoqH5C8X8QtzHieWuTzIhKxJq6RQ1ZiLmAy7f4hT8LL3rn9p5UE
5hqBzw37Tiq9SvsTBGTgl9EPrX6uMHeBodMI0PglWFI8QW66PgQVSMtoUCHEII8qpLxSPHPGTHRp
cvUYT9NM3aNCHnyd93o7C3FrWBg7cyLf1nlrNSgRg1VnGvGTEn9sudVm4MOIRt2FDQRdCT06uzvI
SKjSMQtUagNNTwNnVozzu5ZKShXNuXupFJF82GGxHHSUs3TAAMl98+DFJ9GjQicprjkLWqb/QSLD
rjUAgwlDE1w89PtL+JWKH73a/BtLgxSuUBqtHlJ020+KbOSgHbOhpZAJM7mFw1Dzw6e029e81XQo
hMYKvTI2T8elLqGyt6tnWiZmzgCqHllS3Jl14E+VlIRQTxDv0ajkv6r+RL1OmXlROt1nuuyVOqfY
EGgCTAL+ZSucnqJLGylhPFQlyBS3tcFPg4YW9h80IwalacOzJCFWOldVAf2mCHSNdsTQaBlzX7m2
oeYYiVu1XbhKRZBedLv0/dV8WQ2lEt0CWRJE/Q6LE/jcJy2mxig6QdXchr169A9ODciq0lt8cNNN
5Ga5LOoSG9GaQhL3jFk3ZoMA9j7cv3vBaDnspxdsVg9hTVADzb1Ji8nSXOHGHjNsSiQdgRmk8Ri9
riOk2TR5LTK4p2aZHT+LtWWqQPATvIlgcszn4q6Iv0TFccySuFnXLYLJIDnVA7oIz1vbzgtTF02l
QAYr2zIBzGqhvAc38KjsHOPpQcCZC2mPBtPiV6BrmX/PTIq8asCnE8kCw7FkkMSTwnSw1W9ubDVy
powRzHk2BKFbDdYBsIyZQGFocFmCdTmVD76AQQOhs1lciiDjr3OCqCJjIGYmfscUXEcvmRF68Ceb
p2vmeig0POAYlOPZgWGXSdDhkMe8JUzaglnXqPMU9LKjPz0bKByGENCcBQQTymEp/m/+mSlDu9HR
5plabKZHnkBwuNOuoLKqj44qQcnrKSYCL0PbW5jFsMI5yToYzAoe7nUu/aYRqmM+Z5Eo6vjQphDQ
EUZ0ewaXFo6aZ8JhD2VgMfbfggL67yQ7rFWsKzxlqlw9UKjlHPvSa2PjGkNznmUOyD1p2Z411GQP
XwFDL8a/LtI2t2/EjXwZs4t8xfgXX7SjOyiVw/t+gNclp8qyX0SSb4/x7+nHhZevxcDaSO46kOSj
6GTrNSxBgdRPl/7nba7FqR/59bpSUXRQaFdm2hMYagsjwyEocARpCGKrh18RxDop0RAimY3wVkx2
a3su23T5jJEgdsF0JO/Mk/Xhmp0cGOugl2nobf63zJIUtHkm5ifeuDWslHKO+GExMBy3RQ/r2Gzz
OyBQu1BjUXtix+IXh1Oq2Jfs862pAzNud1jG/N8BVrUDZ3lSfBTrvZI79y+5mc+BpzwaAxmQ2nSb
QeSP2SBjGeOEnaeg+iubEQKT+ViEt2VA74qFlrVL7YJhSWMlF1IMvzJLxk9utjRteqXwynRmDB44
pQwg+eXO8IxMpx51qEaKSE59879VT+3MTFIzymJC3QrL1CqjKdlaAkanXc9sWS1u4m8oMZf9t3p+
IulGo78dqnN3oiD1f02EjX124cyVtT2Vv/H9Abrj/6zSQDRWsDaWSKnpzWd2CoHMRkHNQfqPe813
dlNrm7hmnysLd8ZdpTpVYMdCpDoAfInEpNWRj4FPqLuN2BfFpXnrt5ziz7NzyTPVdmqOPg7Vmuro
3slZVff8uDAoYKkJeBvCgodOsDdOoOFNmrfiPQO2m3+4RQRvgL6Lmvs2bVEj8Al0FM4P+xQUspGm
srigd0YysHzu7fSqc3g2Vax8hCxADgrt1BrdsWXbohnk7vwanEZ88sZB0QRUPSFSkAXJf68BYI3G
w6+8R5keiunQQoUl7Shx4Ik/UzSNkaCZ3UqZSYer3YgrpPYfRq6V2oxhtTmkFCkj5St1feuSH/d+
Y+vD8jBNVYle9MXfZxS0dYdNsGH5EUKDuyfTWScDRBxZ0/qB2G9rrzYZV8oN92bDoqQDEgzqQH+z
xZtGSG8LNFamefZ8An3JL4wcjiE4J6wYny1GRqRXmQvXRp2QPkK4Ym5Me22xcqSm5RR4CAk7t8pz
5vfbQB23vKHtiWqMqaCTJ0FUQWzUejTHFcmLnIgReVpr8sRBlcP7oCtdBJ7K1knYQyFLtjUNrH6k
9FJ0EbJCr1gvSVD8cY8/2/5vEuvuJGBJNo1vIVDmBbLYFHiUC6V1e1CGvFohs53uvlzgsRXmNqXs
74U1Brl2KUcRHwAF9NhkRwkeM2dyAVTmXryvSFp7S/yk+p7TjLrOF/u1AHGCRPQXM25t3Y8MOwrP
Uj2mK3ABlGs7wqA3KhmN4cu70nzKVr0uYdedap+qoGAbnx0B6fc9KTSB12CtFnOngPtJKEHJKF4Y
ghkCNYwXL1L6oE1k7VL4h54dlEcI8at0A88naxRPAWl0srnYEC1yGa8QvsyZceM99PysZg2K3Its
C4bw2SsMwZ5imlTTKytfqshA5qGq5ewMDALgBZp3Sz14vnWj2N06iuJcF1N0QSwt5O6a1MfErR1T
AVQr/ftRZ3bJpG4VbGKwepoD0Uh9QDCnrH0R8uZm0J2N0QVyhVUVAynUL5YnS5ycd2/M+tA8V94T
AqNj7UlmC9eWt4u3F4ch3W2DEmKCSopweqlQaOpmjyEK4qyhRPyZDQtnfWtUqEZnSXX0iUviJF3z
paC6DDVHHTJlNlY6cACq27LzGxKoo5QfnBJu9S8KoBjcv6+SaCGa9SMX/OOLVB+kc9WktVR4PqN1
S1sg280I20mGCjEynqDU1vWMXEWRfRU7D63eYvsvZzE8ZxcFJaOgSf91MY4nsPV2UcUMdd00eNBA
JEU/b4T4rHZx6BRL/8E7jkkrozza9H5O8BP5n951BVKAdEccze8cT6bvp/1dYDDcIXbEARgRhkb1
vGiE4E7ami5J3id9tVo4sbBbPH+xNuWJ+ndGNdtw4PfVrvZxjz5IojkO+O12oXR8KDLdb6WRbHEx
tcPnd/StboaM5cz3kk060/dNuGmxPMHUeYc3Ow7JIgaY1+sWGDLHJl9qHkVYQkr3+tS5tfMXarqe
5XWoYOmF14yFGvDVVl99jONcJSvZPH4jmtqDfMJkQxcxc5tQ1RmgcgwcPv8ipJ0v8Lwb8Q3pHOvB
djeGmC6cX2Dw+qj2lawJbbF1TtUsXeL4eDMp4I6BvONoGOtV1pjWmzTb6aXyuDhpCrthnGAxM8KW
KovsC8BZqMlda/sbykADCrhN0ediVjkbIokgT3AR7BmycMe21+jbM0UgYIzbKooiaWctJB5t4fSJ
7PmQf7ie8aWg8n2JhAW4aj0mAqEuOVWgQ3FB65eoX3efGdGLjL6tuQ80oFkP+EWFm7tJoTcBkHfM
h17/fbRUCTTIKIRDbG6xnGZ5VnsJ+/cVu61gsewjHpezcQie9AFwc1OyPIl6a1JHSY+GMLv/S1Qj
I84MWz3PzbjQP/hjB3dFl+YmZU/UFsCAVsD6q3Z3UhbR8aP8innTr7uGJazb7LwlDruybtXpFXk4
Vj/31Rxdgn7JV27xWHeZbacDR8S4ggofCWD3wjevqPZSsEseMXn5vSGT0KsWYFA6KqaNzVAZC2Vk
TyCwOdAAD7ukt2qIIDgmtu4BjAmuVRUGgLg2R7u56XkpbegeWpnVz1YiwX//e/if3MVQ/vVAr621
pL3LB8KvUmTrg9cNdBbE/9kZ9930mbT40mbk0T2QwjPuQMqkAQYilQVYy4m3RRmp0TD+tHhPBtnu
eYyWWQzdPXtWhcnG9o8BGLtQg1VKEBLp/VfqVaXNUlWCi1vE88q0qmRbs2zDInwiUV36CqN6RXsW
WdAjqwbL/JXURDT4IfJOZXnTZQf8peqkr2nRqbtvzAdCjLm7bvAV76L5goUYhZjVRFmIUo5qkX3Y
0KH4fCc/A37n4TWp8i/NcqAK+cJOoXNMvJjuU1/cPKd7o8O0XBcsuInKoEDgI10jD+0mR8VjoI0K
JubzBbpRi49eA1aBNrk4LZAQ2oTFxOI8PnLuqoygPzdHbXnGft83AEqiWwQWsuOO4N1ZdEK4wX3g
AJ+4836z12VF4F2M9XlxwPHRiIxZ45nk4dDR5cdCVvsqgrrI4Z2QeDklIvuSoYkP+Ppf/Zv4EbtT
54J4wh97/G6fSIXpCnB0VYy0wo0MdiVeBQA6/ZR461Scd86Y4oTBpRJe9QtCIIrRqzuoyy9DtRHL
JzhccNjUXmUxRqMMTzyW0UqdU1FyHvbcE43s95jVI+sSX3orHH/iqoDIX55sQoAEtcTW1ht4dahc
um38/im3mtw7pbEnwzqo3ltTwhxSlXf5DYcTQgJBQwLzT4JXRKGRv/kK84gaLRqkj738NOHflBmj
eBaNYhm97K3EAnsZbEfcayk9S5yr/8nSAKGcY+ZlMBkkleIhesCYdq2jEFcLWvRj73Dhi8qbHhd2
zjJMm0I4D3qkTLz750otB7XcLW+iQ9f9JYh9YOIaIufaG2Ek8HLsHfwfyJvVr+vg8o64SCrSBo4Z
DZZnMoZrtvzx8eTZ2ja3oAYM7+5dvxRVWvA0MyL5CBlI15xVejevX4CNE4Pp5qk2wrcy8wE4P2S1
UPCDnISP7sDeUUpFHpfgAx9dgfXpsDC4HcryhEUW9VtHY6IesJ7JTh4/rliQIR3W3zZ+fLbenFVU
yzRbmYEUnadf8jAPSYFg/qVo7ganW0jnfx4q5v1VUdZ5Y48wT1FQACgCgF/6uynvqOP3wJ883x7a
39+20eGxB1IQkoNGabJPNkZqe/EncVQ1D95rKYeR1/z0zH0jCvhesud0aK+xTHYzl1wZs/BNGfqq
NiNapeLmM4QOeYGb021UwKKIb89ryDZZGOIyKk4rZygGcBW9ejd1jMQyfzFrOFL4RUmVuFYc2lag
+n5KiLY73jzfcAdaSWi70GTY29U+/tb71TYZ4qm0CAEkDXQpdC3QQqhi++WDT8I3LbFywwdCf/Pd
kenN3TiuIfOjyyE4JM5GLFburoTTcxEUkTz6D9hhADV5uBiwlan79gXzX721Aer+2Os2U7Ywdd6G
VZ9pCURj3yP7rFKFx0YMvshbcV+rge9YgFUwNkC75MadBIOjyUVpd0kgI4eGY/RVpn5m3BMhK9Xv
7dK17tirISTzVmLt+FbtbGPu/3D1jH3JAwMXXsjDYC+/oLfURaZ5s0Lim83jiyfPE9JObIkUqzBw
N7opp4U9/pi9LmNFfoIL6ez/0ISe6rsjSQMWaDrXbkrlLe7LXIMEIxnNz0+sCFViG0MXTyim78Vk
kO88mHQ/gZIu9l/q1t2zB8hx85x71xFdQK1uNRxxHZZnzjZ7EZKSZKyZQbUI+HNCRB2jwxxcHwAz
SbXoimb0fZDro0lOrMkfurMokPPAmL/eASVsrKBBeVKFE/awaDV44tm1kqdWUxt1Ur4AdFws1CtM
W74fIjZPJFtEUvar6386nye0pQAqYl9LevgpSdTw9uTbfMfBZCwQkJglIB7JgYIZCh6KRNsqbk6q
Vs5TcxkaE8s4izvIPJZWSCyyZtJ+jlLBj1fi9/fdbLReuSgOjPr3hRa/H9JnqT0G9arpgA6UDCm8
mShPAEeN3BPk9ebbW//E+LFGgEwnEUEyt/84/eHS4hC9beMlBwJ3prpDzHPZxKiAKP89jDw8VvqP
ewg9gUk26N33w/HTfd/yytiDM312mgoCZmSkGRiGKE9HRA39VnbcV3Dv0jmJuF+jwNysvVrhO4J6
cNwhj1d/aO2jz1rNYf7MYFYBA6XRhkGWPo/TxfaGEbGsxuv5kdgDCobUY0bTjZ1Z/DPKddKr4SOa
bYmBkQX9ZzRh0qT3crzKyGHW2VcdDdApNUclUu00pq+Kp+A+e2sPwkui4KRYY0diCBNwPbxfXwq+
LKwsM3ajs88WhRwkXAFXSQ9on9FBPFEVaDweerb8NE8fSWpVWv75aWcjq9E+woRT+5jaYUYFyK7f
jdL5jT/O/Xs/1iSeQP7xNX89ZrcDgNK8Xz0GUs0edLHxCjVZcHEO1tPhePwrZx3dInbl7jn/Ilon
gs4wTbKHGOGpNlRjTycogMovPcBz5YW9E3XJ0dmK+ZiAI3He6CJ14DrCJd5MmDlAa8SEk5Kz6NCO
lqU9Gc9PZbs8igpSB7FZLk85weG6rDmJKEk99ddFMzp8+8ycOR/QG1KWjPIo9qaiqIgfkNj3687x
IwLGJiRhBZDlapN8gG7u3K6+dDUwO7qxVxn2lMrpm/fmOtIT7gdRzgqfnL8DC7FbT9gW88VQnzK+
gc9XvcbiUjDlVW2hTVkbAb1L1YDGEhMwGOZeXSbCJ1RvfbNbR+33HGE7Tgi7eRnvGEpaXSqJortf
PVXpFzOBFM8Rn1s/CSq0qVrSPVFIqC009Q+38r/smLGnjLcXh9N+Jyw6Ug//bvbG4AnGByG5Xctm
kwgcBaWg3lbtBZsm1xEc27cy5nZ6fTkmwptf1/zVv9xRMcDE3Q1E7O3+HliP8sl0YLnbA5kHWN8R
wlWTBuORQXXWRCeUdCIp/u+dzxanqR4dkuy9jTI5/kzdFLJMd9A0XCZDD21Boj8vhSU/vhflZAaO
IyBZknJa1p7LDoQ0l5n4tjTPEOfdRV9AFPCB/3LUGkXzPc9HnZWAcQ9d8HAbJVQ/vQO9TSTZdnjw
CVhlQPWnDkK3sU5ppBH02q23kK9dO1y3QmDO/tLPSsVuOx31E2GAxPq5e7lMt5U+m3LEwsQx3PJ7
AVmKeFEBFrKJjyzCdTOCkpUKOPWLpPBD6cW1DKI4eDsvu5BypDFxYFHNACpvrMJQIgOAJSvbQqg8
5HDmbqSE6GM+VHeW7+ePGLTZnxIZtVdmZughsQt0l4qmVRyK9AmF3eoaf3lR6ZPgHACDyxYog4mY
SoFiUbgAwUtk2LqJtEXOSm9CkqKulBzfl26vFqkDb7NB0iysCuj1JeL0E/f0U88g9mfM3biYUxlC
+XaeowRNRlH7a2rZD/S9YYmK5qpV0E5U2+iUO4N+q2bpbK+1thZMccckByUU0bxAT97+tGLkWeMc
S8o0uSSfUhTHo+Kc2ZVVEBFwYxPfzAn2KH3HlWZ8kqNtDO7JmnHAqYgIgXLzCj4cMK1UONnWMMDG
h6xZ3e13adALL5zn5LtUKypTwokgNqnkkJSHY2+uHBgmoU7D0izUsSuoSpBCziByYwCNwA5JQ17C
X7akDpdeLKG7aKgd3Qe3JjZ/zydd/5WnCMk0T79YTvZt3b+kTwQztThWYAVxuNdqkX/DnnVmnA85
I3ri9TGNpQuUJ9vp2ihZLOJqLkrcdlfy3uCVqyzRs11B7YxtBLqlBJ2RMDCG3CUaiqOaEq5KUWRI
hMsjOnQg16zNlK/nClfQB94qxanX6t0D8h1FFtxxk965sOI6f8l/N7RT2NjQ2PEJkI3W9s6Ht3ho
atMsLwCLT2LdgE/y4/VqLaFdIOnVYApON0L05ZEwoPhGERl0E5iJfyB8orcMLYbhoq5sEr+QhIo3
jGBiWIwKUyIuBS3A5xQTs4DrH/H//OI63KUpJk9MHMSvNwsC+iibvL/6tQaw/T2onUIgAdnqDho3
6tmmYk2YJG/iyvjKS11UO3bdlSVVpFYBbgB3ct8wEoG+uz6PjSAUA+I0Pl45rT6r+Hr3G8KASQ+D
jP8+mISDjfahWgoGORiFpFLzpspNVXqA8XP5nFFK7fhz6muQShQheoqku2vg/IYT+ddMxCbuA/Pk
jpl1bj4Jc3RlSpaX/YWw6Yfl4hfNJeSbAK/T6hBY0zxjGWZsvRJzc2eEaJ5akkUREYHM7rlDzuYq
qOsFXI8Rq0l/ILbscXZ4yZfJeTRprNjMyVcBNZMAkIoiW7IRMvOpLYOS5/hUcWrrji96kLccYfMO
o6GQ6yOhfcXly7PG3UlT00Qhz0xJcllGQG1VV/79jVzuIQ9a49s0z1LIDjajNQePsxHZ566Q4Y9h
dt/qEei7r6cIEXAGx8H1N04ytl3O+JWdKVqK5Vs/ItbggclerGaGqjCs9cjpWm4wfkzp3RqIU89T
rggGmCExPc0Hj9i2zutotD7dSCMr68BrMsCIDvUlc4H8XUIY0a5IRQT4T5SjfZfDUWKadlEcjTMF
AShKaOLH/ov8jexjxfy75YrxWzdVGOmNP2AW/Duxiq8OF6Cs6PNcoVI7N/+SxyBslIGc+ljWp4dN
ZyHcaS/A3/D7yLj2Q0UN/eSA3HNikl51iwp2qbLiKmcB4E1EaUgRaomhRSjtrDG5CKq7aJk5sPsT
ENQUPs6Qjq3j8Bsnwidfe4ktMNX6N0DmbL7+3u3z26iQAn84Q4vJJgIbN8M39l9PoFiSnb3wX1C1
vpnZjNIBAXBlHvsSpyfH7Tr5xg9x1n+aky/nbIUJtJ68UKIyzvFLqsz4CQ1Yyv24dK6N3T0SX3gA
cwdNxHrw0GIkDgzJwcH3CDnFcDA+H4je8m2JkOI6/0I1yMzoda0bFYRJfUCTOYBPW4sfYG+NuQnS
ic4av59RegkZZaqpoYuRcPdVTuKISl6ci+hKibJVXM3eDwk20ENqH/h7mVENjCY4Rh5vLp6/vo8W
prTULdA5QKX49jgpguFXu/ChnkU/Aozc+SP+dJhEgLDUXhoaYJ5CV97OrqrDVpX1JiWCt8mpc/YI
rvfbENARaBFufyETQy6ZwEQf9PWx+E9ttNcYHFm8/uZjQdlqnciq0DfMp3FmpI3Bi18AjOE3qlY2
IKoqsQZVfV7AdOxJl/aKDvDIzczl1/HKnvZK56a6eNw86OXoOaQaO+7X88gEogaTDFbjTdBS8MKs
jJPZuRnFN9JxuxPdWW/lJlijlVX540TP7nh3OU6Hc8AHtwqPqsHRlJQdv3atYUfo2Q/x1NN0F/rI
sQD48GPPLaxzJQTQJ1xGk9WOPaDiGYa1zn5doWVbiO+GxUc489XEePi6FMS6ddgjgC27TJfyK+sB
dPfsD79zIupDkCptNSu8/9eNfmL3IJX/eULBRMKfvNbIRyDdRHJ5Cdnvq+zrZu9pcw1x7tdCC+DN
JJ3aERh+syNammxs2JN/dD35xszunt0xi9whN4P3JuJ+BFXUOqm0UmK+Q7vQ6TqhfFvHjeBLznv1
yl7rvVqqv6ksfrI7pw89TBdeBy+4RofESYTg1TRYiEKoSkk6l0cIG4MZuJwZt/uIAa5jW+DMYxMT
TZx6XPmZNPAXVMO8JguG69ONUKWIU3EtMDy/2oK4AQ5fbJsgibr7eKKmEnJznlak1/wQ8f9sF5/5
+JJl/dfr1rfS30grEvLPC7PXblbgx/0dJAWUWBdyvgo18w75j89ypY/IE6Y5EIuUcNIlZ8Rii5yL
TI0V7MEw9tq+b62V18Tt4tKz0d1kLYTvWWYWHTd+CFh7KAZyFKRZBztb+1+bjQ9C0KIcuZzPcpuZ
alOJ+QO4yFOiXKKce+lOCcFetJVspfXnfkB494IuWWgrjY5LVDHNhz09m3M1GBYhgEZhPhpbH6iH
UBBlgJjVHaMFszwTJo+l1BArvMQfjneoweQOnnjcbIQ1XRxY6gCp6LCdI5iR86j0Rz3RziEFDUpG
J/kkJO0l+f/nbFYAze7SPmiDjwlV5WC6B1OWe3dp9C/ajzSNjIX+GFbEEJ64561PN/JQLQk/PpTD
CWDdhZPlxeKDme5Lc+2Mck9amxF8PkhNAxC43pcJvy1Xv8KK1w8NbKlRo0ZxCfT8m9mGzwduRjgi
1mRVqShjyW0EI5tt36f7anjiYCwea9IbYr9oU8WlUYEwUxrkzY/DQrW6vcQgs7ToTfwU7TUAajlN
sVAGnhc0Gasfgyvg/P+SZFWFyLKk0XujY+CvdsRpERkQc49+KYQ6wSookSnp+SRR97gHoKlntiJf
76Xuxl0BnGjVsC2hG0p2FNJOk+J4kx/j+fmFVGyitucslTpub2hz4gPruH24tgoU0kUyuINxZJ8i
8KI3zFH5OTqJv273qE4Qk15NOnvwCFC5+0EYDtG9HQp1ZlnRdwlj69qWufl6YQ6UfPHY+D8UMFk9
qvurOXk6VvmksRT7OcKkJOOdz9CHJJOCyc7um/DNy/4rMqkfU0QZw5l363yWKCMQjVhc+RmWdIOA
pzmSe4KIyW34dCCLj4IgEAotyu/+BGo+fQzHV0cDdPyQaTXVpp0YZU2otYzgy198M7HGiNWDwteR
VL2XeZxVjvfw3T+xaMT3q13TKmsd7FzxND0la8mc7118u1HmX/WYsLPsKvzRpx0zectQKNLcETJk
lHakNM1+CpgfAJkCzU97BqKaitoR9WHgnA/XXMgN27Cgd19gqw2ziAVZERjxmupHb94T1x+Hal7a
Nuy1+1633qcILw01rhYlWUpoXRLtXLEGrX9z1QFoEAKlpES19Vd6/U76utrCPDd8JJS/fpv7Dcd6
BVZpz0pvkLHUVI/8LzUgR2JoCYASj6r1e9dPoIii4BSr/iBhlvOXH2Dt8o1VHHyX6TgOKhJLDoJF
D5K5vcqKEQp8XEZMLYgdQqvAjm29dEstwXi1APkm/cLU3OHH58pdojgO1arBhQeTdZcoM48UOkZ8
03Bn2pUqdsC8B00PNgIWc3up4XiLSzXr/pXCRZiHYrAYfnXx/62b8dxQ1njQmy/Uk1bLdtJWcdJv
p13GKBIe7KyJ5i/60k16nBgQjkASm2gdLRgAIrpvmD2nCp9NlyKiJlo+qN4qtyHSqP/dzy0KeOFF
nPCNXT+LUH8ZGxo/R108dEMQ6jV4utZLAEWl1XsKxSQFvtX56In3j2belBgqByh7xmj3UtWVC/pf
xP0DXVY/qb7asHZ0Q2F50AaNE8M96IKgeeQlt7Ba0qO9nvA91Sl3xZ+TGAJFXLqFL8NMAvIyyhwA
zCOnjj/rVUxQbtvQy7gwfUEHWi+cxPN9c/xhR1BqwFAWNTIlI/lD9XP6nIS6LYCCIuRG/JGc7EXz
uN8g220WnUElkOQTR3VI1WoNRt1Nnp5CYlQR2Ch8njM40oreGhISkcj6qUW1aGQc150HxAtitB1m
YfeDHP5MJRZsw6UNcU5EXalvyKt4A6/EdGfjY/Lk8551KZaQmCJXG6MpLQzAAK0b3VGF2R9sQ9AS
hnO35Y3V+8/AWSRi3St58mlYdxa7Y+FU4mOa95PAbX1TK7Gg8RYGEGITg/m0MCqhHPflcaMfImQF
rC+5yB04sKAQn5VzSxj+Ey2cJjRy6vJlg/F+N5akwksu3x6WoEGOtAG01pSRzCQ78/RgL4Rstwjp
VykISpgWZ4sluBWSJJM61zOhL8MCWLNo+DGwGg99JVx++hg9rr7Kjr6aO6f6riTE+RSNYY0lOmjS
F1pi+EIzqw47L0uEdGMtu2sBcO4xqrwZV9055AmicWe1fnrfbXMRGIuf8FsjBYxZSJ83CNG26B1M
C/DqJIxJFw9wFmfeAByRq12lBcMCz0GLU8QXO5hXhfEUVOv55YF8Vmxiq664dx/vk+PPTsO0Wd+p
YJ8aGutVdmnUxAPqXnAMp5+PvWiCYPmHf0pk83NjiVBA6AwFZolVV1DCeNXwczOxIT7MI0LYZFeL
V71BopNO5SoXYVg52qYxdN+XGNqvs4ttAAcLD9uWDCU6hshQkLo5mZEYkMMAcEncELXcwourOB0F
6PTBvNxFtBIeW4iGodmZsHUDGgDA4xRvTMwOiYzvoElY41OBYEUeSj+92+ni5s1XbXGKPwGh3mW5
R3uFdky5M3BDSYySeUPf16saEzzAVQ6vcRYxxjz9QH/K2xykvjGC4uuh345pq3taYo+HImB0cYxp
44j86Wm7nGNj1zHFOW4WGbEhetJA6medWxbR+uDx3YbaQ2qq4ilRS2odwHdlf1BhANtjauKLQJ6S
K9fF8EbtBS6s2RXLFTTsXPl7rEJcg1szK6+9sCwRfx7dTlzPoqMHhGlbGxBeSU+7Y0h5TiP5FwC8
KT+tna9KnY52Kb1QO5mI5oRFmcl7Ie5lzEZSj+DJ67jLcTvD6VXcblszDAo4a+AUkzfvPnm0RjkC
QE6qdvGBJI8QZINrRGfn4LAfqQhtS0B3RsRAfzTwXIt4oeCOsN4yt5IlXQ9pGZKA23Y/PjfiiN3M
N9AQKtBQdJp9DQZiL7Ou2Pkt7D9hzMznsS8V5HIjPwn4k4Urs/UWYVBPtqdYqfpXXHP7xQujA6OK
92+eE5gLrC6Xq9o+1Pj5nO7SoG0bMy01mIocXEvB0a1FeFcgeKBvhOfFTsy8S70tmlZ3a/0L8vy4
dihnM4HRumI0Mk02GkVuoii9U5rP9YHhFwR2V6CKUXK9QdPTmhQmlodkfJ8K10pG687o8wF75Sp7
cxpzcYKfVZPMaFF5YIf5UQ9Tpr15jIeuz4FCyvJCI6YSjtX/qHPyekXiq4yp1tdYQs36XMsQg8ac
KddMnzGRWkPxpHA7MDrp4V2r6KfLdRY4yJRTkSnn54u7yLj6YwwKrYUnehCAYLdl+OhiBYuIHzJr
UIGhBdKXiyt2sa3kSavWHAXupEf+6nnvIz9mJXf7auEcpEgU9TFdC54x2kNHHZXtohBT7YRlXUHC
ft9f5hwkR7WuF2hmEq1ujkOwX3YnJ5JcWGMfuCsEZVcsPMn5G8833SLpQe1kqUA46YooxjODUnaF
BZoltbJtAiqFH8AskwJxos0SgTbZKyOutAAF/TiLHWdn3COZfbEycgxQlLdVgYFh9q7+D5qsNBYh
xpXRs/eIdl4l4DTQ+EFu6dXKCSBwQS1LHjf9a7wN39P5kaNsnE+JgBXoj1AkndX/9CC75jJa4XhO
zQ+319Qnux6ZzG4KZyaBdA/cP5c7uT3hiIMebOS+9MPqXmsrvrWVO2L2e2mm5tTDrcvZWXjCK6xw
lGqzuAum/8GwUb5uk4V9YcH5UmkjAbOYGoKKhDoxviRs3as0BC7yU4n4QRf7gIbdVi5en1Jk7Us9
lV23CBfokWyUz8gfQCSjxv1kXp0rDYNvyIY6XciYI9IW90hamG/IC6/HPJA5VADK+jhXhqmH0FIE
/CsIifYYlTTGOeREpoe1yN4N9qDz3+VPCLk29BNqYAPf4MuJN+69GXa2N5s4yF9v2N11B+PwoF16
/lF6mWYaHEOUdrkcoDPAsduZwUAGeF+czdVLaNuR9lIAWCQloWrRgXXqMrBUWuUZaJGkCEsG0tO8
lf9FImRGA3fHWvIG/mug1Oz3l9eg2mW4xdOTq/duJ/2dpldqPTUv8SIJPOfsNXa2var+C+39WYt0
yoe7WtrQYxPslHV4DXy0gwJs5XuDBJMmHwS5Vvs0p6v+g+RvHK/4ILgXamVsxVVHW8de+OsiOAM9
xCZ5xzHUWqfe3eoPeH8YwCikMDYIC/mQM/ABbvKx5DLKKy6of19tlfeWv57FGj6Z4+zK1fnF+MY4
HCtRbVaOv4Jol9bXb7a9f4ZKuIBlfH9L5t6aSp/JVzz52SPgziXJ20MJijd2kiTVH5CNuI6t1C7F
IlQr3lKm9P6BjfPmE1e6wyniuZLBQhVLdze5+Zz1EijlAa/0HMwSyXV6P336s4hKiNHsfI6gc47d
NZUb8xM4m8ODVb8VqTCfm+rSu+1ppuRZ5dcOibFI+EOjvSfvW5HEUgsGJZedUpMapAtW7E/cEHe4
akjsuEb4Nl+19zc2NDmSUqF2FX5Ro52rxUALKw5zFFHForOho3fLwoyYF9bAhfzKs5C1gjNzaFBz
gNPk3vQDpE/HBtv/Z1dYn4hVeYriJ9SvLI/cvSJDrAovMZd57o46vexcLVlhEeM5+WMzC/FMJFXM
WJoGc4z36sxNHgYflIX/wWDHOGib41X0+9B9MgG6eLH/yhCiTwkIzd0pdgcrUU1rtEAzms9tHBdL
65noq4WdbuiSrCDqxMnyjbqjx4Sw8RLcParNz3tFEqYQ4yHIueOTILihkYbwoJH1/PKCo04qWz9o
9wE9GsGj4J2k+E5xeOxRAEsML4pnc3hDm3BDYG/7RNzFa/ECiXECvcN0BBJ1Ly3qY6l+rX+x092L
DC+pCDd3rPav6EvAP7dSAjpdGzLnGkkKNiOvmfBqA7me/aUWfqliZqgteY2/eavJ208YrcJRcV6L
LzgushmazvqMHBkwM+ipBqrT3G+c+jc00Qe9GZJGk5ROkiqlBbJ2BfR/K7La+taXzEz3KFMcUfTm
DCO2llhUFIWqemJKr4Puv20ZAWY2qAr/z5nDw/e3U/FyWQfXOdMf9uceQoFJevn0Z54DAgBpBLQE
vH0ayqxcf1hl2ZzZ0vjjTBPXu1ukG86HcZn/SrhfZ5UsEmRSd7lT8Dz+9/PX0czXACekXE/ouox5
Y4nRkuINQEj70htJVYSLvG77KxWhUNFNuDpZPslc4qJ/5s0rv037FajyliORcVZb814jxs01H+tq
tcYQrAW1bSgHw3pwVR4X6HBRiPNkQIcxChvCtXl7q9/jlOqx9YSDfc9dV1cfnRQG8rBBhR0ILDqO
cejMg03nb5B061JNOhWnv6IOoGoY+wRnm3LpITpE0kck+CPSMNKuqt+uuyCV9/dPDKOaeU1fLhD7
eb5H5RwIpRGq7SsH7qS7xoaNCY9FQ9YdVWaEsWESMHrfVgUrDQzxsIV7C9jj7wUAynvpna89dKIq
ynfg1ylPkEOPk70KKRMU11LsiYyxgPbyBuu8twPNLlLVTTQr71UA4LLyFHCAnpkgfnwGdC/wk4P7
mxtjo+1SFO/97n1YOhLq61wWv+sF4/XAxen8JW079LV32QJs9XccIRwJWe/eMAGz23F5H1F/nAgb
BCVbTc4OQ4JmAYwjkyrc0kHKjoHGj3+RP4/Ixsnn67/OK4TMsw/dvdsGTHO65E6q41MQJkl6fC4t
CPVsrgqOX8bb/1ypfFrOzwC/B0vNWau91UMANFyoGAh8THxd2lmmiQGClgChOV88axmabnWKfqfc
da/+1uu5zzDPfEMjgpA32HNyFWJAx4euAQetF1a/GB3iD9zXnzSi1Us+lgEJTKDVKVEXR+CY7Ved
++yKhO3lRQZixUACaczwxNdtWBIB9PNxEpkoCoyixOtH1zhq6DtOacTRilqwvhpo5XXT0IrZPn2E
8GHBeDBU1PUTHj+UXWChNegKO1/J7BR6Q55rmtbjPdggfZbs+yTL7iKwOePOD//Wdn/YhPmcE44O
cQ9F+HGd/VxfxSV/8lVB4MTP0aMicgWN0zvYs4sRHoEJTis75eZTftfvvjZQT6yGaWX9n9aZTfz4
bmkJl7ql/I8XFzGjDO3SF716qJKg0xN4O66fXSxX3kMxx/XabGcZRQm4N1bTp1G0fPav/aMMpHvY
3++tzKMkZcG0ZbmR5dqwdBe+Q/8LAQYSgBW47t5L90qty/m4ti54nKIQMFICdLZSGr5TCx+Jc6W/
Mzf8QbqH2/KuISoNK6bH9zfbCQ7diWNOaF+FMVSbF+AHcW7BJarmg6zGwMQnLN+q2WCN3SIN03TS
t0+p8VKJvpWQi4FRP1A8yGn1ChZyEdt2YDK6nTkXi+uxA1CjvaZxqLR8PB7+IaGjT8uqXDNxGa+x
hz+9Dl+XM5+/1qHx1PxGMfdKTnmWt1Kk3ngL8UuNfMvikCzuKlD0rdlgv2uMPseaK2kLspT+XoxL
OjEK3DXcLSEFfDtDwLECp5i1L1hJNWgqjO/kzlasr8SW28YHG1O9VpI8+sBIYMO2BQFko3jyXDCT
SOOcl4YdJxnImLD4xbN2EAjHFdgepmUY58BsNe8gMdSz2TFogd7/jALCyV0KfPc+ZWrexI/t/FEk
Rel9qEtI6PPl4Iz7gK3aUJIMahZBzt2yA1dP/VRURpteIQTeqVue/wDW2hcYoII0UINBarfJCrOu
1fjxlzB6OdV6H8Il8fehMzVMZsLgPBztkjSnfcpDZpDdNo472Tjchz5Q2yJi1sfFiXBR1KXjH4UM
FbJsA6ULVeU4iZVt+x6TvyRbW/smm5IZF5knM87ZpGJbjzlK683BOgBRK9Iasz3lm5OGq4ef5FEi
yFF8/SX69YZVZGq/gslAR3NkV6TCMMmKYcRlYlHX/oVj5RHOMUMGr9Pm2BpS/fykpqmp5KCvboDJ
GLjzq/dQR8Q2kFbI/LjyAsDVx2ta7uTlAsg8bHDw57PZKI5nD3GjUHPGz20MwxZChdjHYt01gDx2
E2kR1/L7Lsyv5n/wuRftCMSmTHG+zIzlE6dQyITrHP155ctMTFG8t7uH3wyVzsbN119tsvpbCOLR
skou9lQIJ8dmw2LnqAj309edsMXm4ohe6g9qOuFaeKhrD7GIorUOemRLIDzHjb7EYWHoUdzbTjBe
9f1Qwq2M9uhYzySY1rqc2DI+te8f9rTyG3/EhzLU8D4WFOnru6SX9Vzwl7RQk2aV5/iuJDGLRnNf
7N6aFMmes41uXr6LPeT8HZVYYqp3BRZiwyogAmJQeBH9+6m5JNSqg4DGUQmcxRn+6kHvl/oEGsQ8
PtOgDJBFQ/UHb8GBCZL1/rycrLIt2WHXwDiL67XxK3P/5ZhHsejyBB6IlZCzny4F8kdLdH7BIZty
oGtxiPpRLRhthXvlV4sw9KDesO5USWSWsE6rIHL/oxwjRR3eo83LML/cH4HU8JzYbxA7ngJJ5ToI
tEGuTnbc1bjlFsBZQgun8amXfguww4OahnCD/cIIa8DMzJ+2+sLwDQpC8IpM8wcENv/3fYtBrkfj
ekj3/7EfMdzT3uMkuDoGO9fll8NFkWNP6bmrmkCK8rktvj9XiGwjM0CqWfdWOU3WlIZVj53j5znk
t3VmF0HZPItf0mgIxOWxG5s+7ZlN4TRYrMNMcQAxzyVeM4r0mArMeMfIT8CTVnkEHxidJmve9JsH
8F+F2jAybRAQCK/K9D8voq2zuGNx8OZSRjB12ht4I4gphd2pEmy6JZPtW+jEFuBgvk/x3BnG2738
BtuX7g9D4cjZGtoB+SRoAeMBBCG3hI3n2VhHUiisqEfiVLW7YPZy3xF7Uz/PP6/qY9q56XkhHY9j
fPuVouP6NQIkgx8v9gRXHTfRG1mEElWec88/kmuSKPYDmNpEXQKqukT04nLblOhlFotTODcTfqTl
8D5eyf7jur/3xs1KX0GYmSiSjEimr82zVxFEDJAFpzDXHuG4yPYYXySHggtr8Mmqha8BFI+aL+Sd
yHjOONwz8yykp7y/Qn5+DpFhfn0iT6Z1G4EG7odB9Ktklf3Loe+GYD4/CRe1xi84motIFqSydjfa
y1b3sDK1cBbEy0bFsR1RlphL3KodwQxvjtbQmKQVLLrfNLdC2p0vDzTkShGw2IYYvkvx2YEO73jn
ACuEdFaZL2XxFRNL0akIuAdLrd/90gNNZ44YmGwLrKnuV7yN9UmGEDC6ZieweIJZgo5UNIvGZHmv
lDQQXxyRXPXhlFJt0/e01JRh3AHFla6++A3q78nbp8Ij0kFQK0R7kbJdqk4Kc9+5LrLe1gQv4dWs
8rRL7HzPdIGfgXVcpM92U6fYN3LJOTnijXhChKyhPIZ0TOoVqgwgEtD0OYXeixxWM03kHwMS9JZt
YghG3YGP1oxD2mVylnQel7piAE8dv29GwAdXN+6l3A4/htq+gEdgggIeBUEy/BsQ+3RAOIASlqsC
Hme5Q6/QsMP4QPa72Vb1V8uTCMzSs+B0qqEapJsD4riTMkUrtUA2X9vT1spu39L4f5hTlKYcP5/S
XvTY9GDqRivG+D8ol8wxtKJuwk8WOZPcNFIxzrafuNDQYOzSiu5ts8Nps1+s4LLzhAcdi2geGM4y
ODUV/Eo7yKD+XeE1RcYB+tbt4anxaoB102a22Ofsiy7STYh/kMuk4UVUJCxDvg9vThW1IfnxZm+r
aduF77x4vXM9L7DsiR2n9/rs/b4bltfdaJ9/2wIrh2yp0w8oV4cxmJMD3fnJa/V0sRVXkFWsc0rt
kv7SEWNkTf2zsgju0gwmhr2mV/lMlS7rXNOKxn5qBbFP2PK0v9sW2qSUKXTQO/nAk210ZmVbC1nD
HWhVA2vV32f/iEtDkU1ebeAnpsak4KqItFgkpdqWdtfJG0oM1AhrwCtIFAxFU/hP5kPrp/Yic/2E
KjzcWJP7edFL8I4pRa/2KT09dpmYGulK791Hcs8N7xXzrUhL5Y0hdESSc4LB1HcZEqmMUVTIozGF
0aCxx6vdqnepH+A1EsQViGNy84goHKyRNcriy5tX5+OVGb7PCaLZPIGHb/v8q2uXqtiKMDADxTSg
WimAoJlkD6nP0pznygnfJp/5GRiOpR7EKMvmZ28vFMnFDkVLIYt8TfQZdPVobK/BcLwoko7LwYkr
JKDFvoYUH7fbSJ85RqK0vE9hh2C6GKqYvgBuLOoFL8lkzHl5HBP4wTnYOG6lFZofSCxvHY8+ImrO
SLv0bUB6P6RftyM7AqClK3eoogPySQJhsBa+uw1/smogJ1jq654ylO7j2rZbwQL6INbTCB3HqCPD
xfhETFqCsXJXeENL2ray8aMw3Ru8FhE6WAOo5xF5zg40Kq7SMPbxqtZQPBYVfd+UbWCd/1kCj+QX
/9yN8izJgn8kVKp+UJgxkhOo+JDREWd7e1wyO0WI25VwZ9/aWd7nf25frVU34j3INv/8iL4jW84J
lbOyKP9XQjrhFJbh2tW1D6yw5rmW+4dRFRfD11IlTGJMvtj6x8jJbYAEjEReD0Pys9IDjhf4xTku
N5mC3KXMogT7287fIoaJJ3JI9sSMODCxNvAgqOQv2oarSdULAAY5xEvW2pRlVR9nG2HYaeRGMeIm
wuxAUoZANpXlE1XPPY/TqljsnAIV6/3cLHHyo19Hv0HzPyrHYPGwDGJYKTUrjJUatHucdcgUuDUH
AOjD9nCIuKiQ89IHvqaX8qh76zg7CN4Ryvhpzi6g4u5QYNPSmw4rzT42L8W6fnuw3lTJKhrUfVgD
8LgWpNF0CezQoO0gCmIYidXrOJV8jko8xaRqDvXqGe0Ozhn60F8e1nUGvJZT8zX4qaVH0rZdP2Hw
d2GMqInzBOrgnY4Yz4YNEtDZOjw25f8lAcufoJHp/+LXans8fD5fIENyA41vA5jeYkSJhCR+f2su
fRncc8mQe22aimDCJUFnYMdh+10vKIgCYEGP7TOvoOBz9mZc//T5X4oPajpF1HOrDqK7L1OhclIR
s4CJXPMGWb1nL3FLwro+sJ1Cyn2F9UORBmWyeSV/+nhuoLHUXLqawwfCMcb9sakcag9o2NTupx9z
1zMVdRxPz37LrOFmI17l/mMOQUqzZgOIHqiD74fOKJzpriDa2Ai7FLAJYOyWIeI4Q0oSBZdWnNVW
lvRvC+hq/ehgk7zShWxTyoenEYcEUvYvwxB+qmK6QbQngYYX77ift+0W1laNuAGcKyw9v6kkWFxt
oaf5h1xdQnFS6Q962QaWK4V3feVYht7kSgtQnII5EQcPOsaM5dILS6XS+l5c9zm6M774DcprWeBy
kstE7UfGWfQN2SgFHIibo8IWtVCI29ZrDCG1bR/v0KnU3tYoQrE/yxGF1ackombjqvMCGAPObL+b
dutSq2xREBWbBcK22eSnTPVj14+aiHvOSjcAxDR/VvBEA2QTj90D7gkF9759AB5WWUVMyCzO5OZf
3K/pKTz9rPHF9IZ15s+I/zwnLVQ06qBvLh2an16bciylGYBRTUDk3neQnISK4xSiUtfZvTwPRoXd
kp+U3Bp+JtLt8QWTQTgqGGNvG7H2UH1j2yE9TxOy008VMixICf9t12hjKQ3RFD+cWCY7w9WGGjEx
/ENcfjTL9St6ivUtB5NxG7+USTLzVsxO8gsXZaachX4xCEjr7EspBJ9yG8r1RRdMyHVb6Gn8o0Y1
3OHENtSyPdTXv10afrTRiMzrM3vk08KAi9FduCnvF+V3eVEwPV1iQinb7vFDQ/Cj5e5GbkKK5EIp
nZcNNAPAjSJ1kBXZdGDtTX3jaN9PsEUQvm7KqWmd1LmdRbeKlR2so6bCwcKTHPjjuAZJdOJHcQep
sC4ay5ToQu8FJVO78VNntLFQfTzfTI86pUkxUMoh8m/okOoyEvqXlrYrBMUTQPRba83Iqf87siN0
1h1plZgPGNDvZNbd1bSeu+TU59VRKdLZahOk7w5hEYBYxFNUEhOPHGfkCBd1Eqi31UUi3WpdHrB7
tppVBBjqXBFcppzKBGFfb4Cavl8YfiglHHX/dabj/efh4NScvHz0c7x6JlCJ0jjMJvGUgix3v/aD
afrx5jaddQPhXkGjstpw1GcAmTEG+gR5Kvi5ImcLZcQJddkh4XaB5SOcd7D8Oh6Ed+nnc7GDtZxb
teVuEdLcDdbY3C+fpD16e+eGnvD0gY9I0x7Cc/CCdpcTa3Adt6IjqwKz6TffszAhvsZiKnAxBIqx
rUqVSjRnFy7qKvG/4JMmntTEM1YQPxEd/iK64RvXTCumMNiCxhNl+uctFy83eOZ77mIfeh8Ojure
QzCsSEGpaQRs3+QYLYRNSRNcTcMeK5LTOtT+Jm6vf9bVSFf8YOO6ClxdK5sUTmZOHJEP3WoUthsK
Owprgd2mjKZ5S4eKDqZDrop9cLaChZrI/nHZnBaTNiHaD+NXeNxDfclZlFBt6KyC5zrJP6viCdl2
Eyu+QsEi1SBIq4t/OYB+kV7LLYZMDt4urh3asZ/nukX5qV8QqdY9tUWLMqmLsQJHgpW1tFkK+UBv
xx5S8ENl82xn2zCfb1VTtVKSzTjE3iy/6xEKchDAj9aYPU+x3BqenGxDHmk86nr5iyr/e+GfnVhH
6xCUhR3xmcUT9TXZGdtQ9O6ii8HueR4wAMh9M/b0ByyF0+x7M6QmNyp3A5vYlupQiVvsZRHqLtUz
Z3OBgMXzCLxODCTpCsMtL03a5ZX2HCCS4Z6yEMTbA4S7wIk6TC/zsks8Q6gPnUX32SJzHwa9OfhL
PclKBClL9aTZ7nYVBM6LrDJOQtvJoq2W/eQWvS+v8fS4ADVDJTjTO8KmaHIMInBtboBZc0hpNa+n
JiBYdnIYQnsmjxCFF6B4BpRiOVFzLbO2UOnvDzpfwjJkVz8hXa2rONBbCBH7EM7NR7bdqYepA1SE
Q+wj128ZT8uZAg8hN47tVn8WlzZmV+cKMtsjtniOJZYU9mpWOl9Lot0zp6afosbWjydLK+Z7H/2b
Ck7URjqtUDBHtRMw0oNOQu98uhQSgDVo00Zkti0sXUIPKp4NoghW9h/ctEhnfvQQxGLui6CCWgpM
m/fD+TVfHo75fTE8ddoNzkDorBVfe3UB5YeEzj3KMlpcQvHbwGOItHCKNDyJg7dbYrkEtjSst1Yg
Bf95Ws6TvaGt1cnfR8/VmsUV1FqQmsu273qv6lbHunJ2HPTRKOV/zI2QL+Q8VrM2O3LY9EZ6R7aG
8UydDJBOAuBSF+CHMbny3J092Cxo2nlYZNKTjEDo5klo5vtBnDDhMwTjyKPsxk6aJELI1YYPVFdG
pszY6g80gk6ibEkzfgUqvljIn4aNbCW4niXHcbbSsOr5eRqyGmIVv/mf8TwvIaH/gdwFfJ7WaCAi
fg/9OBn0ni4WFNFcVF5cf23zGDDFozBgXeW0LkWPpAhUN5e11qawYxKcRMvnhBoYfXMZAyVTCnMZ
GJMWOowF8a5ZYDMpijJFeokOEjkisy0oNZmHbKp+vf8GeGKU+cZ3Rq6FsgdUy8YnkWGJp2aCSERt
LHUWkgbrJwaK7XNEd6KADUfNe75noDCtISgwVYm11EfWHSkT3uU1D1K+i+n6n7OYZCecCTWe2HqH
OKfoiRaLoqWDoeKjkFCQYIJ4F+vRUoo5+D3dKC8JIztGxz2/Le3xz45bS/Z1VeUkiqa/T4DrJThU
7H+jLY4YkVGvo0soRdPXMSwWIA0UwcaTX+tjJfwGybjpxNINWFvNp4/91GPNvFJoGQ/YaN01MKfb
z19k1i/IzEU0SWPizzuOX+wcwBxAHjRq9sEl0PZE39nWwCCwhuxv0KMnSH4QnChJIROdhA9gct+U
Jr65B7W4tvv97Mw0topXU/EwljUERBeBoa7eVjfy/OEgRxUD6zuToJquMJ397aDHNCNFkIQlAfX/
S0JH5b9z9SZ52wLluiU/Kb1h+x2vRcW4o9+VzBPJqO5tEnwy+vBx6hzcC7StZXqxoTu/d2Px6l2T
LKqEQ7GV5pyDpbh2g6RuHi5ZtZlTsj9BDoY5HM07o6ie9rVt0etrnrUjCgIKBr9gujNwN3M8NgSO
jpP238rLPhqumt6aqg1MbgrUvSPw3DHIeCWzWilGjFvKHko0W++dhgvYFx5MZJnQmWRECrfx7lt+
M7D150G3Jjp6fkzZi1jQhjT3Ruuv5O7obXoXnnluR5Uwp7IHuZ2KjEuXteQCmm/BaA2yPsr6hnu+
ftXH/tmEaaXM3bhrUB1VdEsNcI177/W23KfPoIr2WP1gThd5yej1ypdLftLz/m/sNJpnDfl4hVpI
9gq56so+KnsdVJURJT3g4mtOU2ujwBPm7my2jCwFByg7bivLIeIhstDE4beIE+17GqAv+hmi6PsH
3pXos2MXuc0TQfpS9IIXloSzBObB4hJbRxx5aTjNnW8xMK3pcJl31HMeqdOxfxFwUNfHWNguvmbc
9WGirhPIJpuFImcUVwv9zW7DMgEbRhv5smib7ArqqoWZ0EKjdgjnzCyw5uNttf5qcfYEmJb8YCE2
mX6pSJfMNfrCfwJ/hkVIonC94D3lwrILlyR1LjXJ63Rgq4nL7y0cqe4yMIfv3F57VGR8VXZWEc6K
Mi0pZOLQ1wWwfDY3e4y4WPYMq8fhdp6NfephaWoPL96Wr+Tn5c3l3MsYnh6krAJKgtoy15P2W7nL
3iI531QFTdjebeybhRdYl3tkmpUNQrWqZbstWLCf6xbnV9WAubjtEdfw6k0/kcjleojj02KP8SFK
ueUVkzVsu0bNGY0LwgHZ3mz1hKlM8n6eMC497Hx5tBMGk7v/Hm5Pp2IQI0qZpaAV4N6uLaiTf9NH
OR3icAAXVIayM2961JF7AgUuuHJTSNzPwfS7NHoSayEEEmmSyhOqG4/k+R7T6AqwVawTJ0pWcM/8
f8f77joQBDRLvhCcnFVH0JfZhd/ohDZwYoJh1xy4JZ8BdhyNQAONeB02YwZbmD56SLgq0Toyokzv
TaFDwEY3FroyhwNQuFA4YqhheCZpWvM490pV6NWBskjDoEKXM/LC7JwNAhBSCdOfkJEUdvA2dL7D
jq0x0uetjuPfD+DC1F9cJEb3OS+Qb0+UtEPMDlgpi1wBFgb9u/s8SU1UTRtemhPaMJWsFLLxYzR8
yLTVyKwY6HZ9gk4gFPmBeTzj1GgBy7ZD1LyGRv24c9jWqRztEDWih6IyY9H8yJdmWf3pm/v3lLXs
ODGUcUaCQ2WeXZjPA13cF9rTR/J6YtnMOTzHvCWhjGIslD/XjqyuyM/IpySJ733fY+n7UGpNf3h0
FufQL5M+n95lXwJtKPI2QVDtLe+8YrkabxYH0wI/SRlLbbElUTViAxJHPpUTyI3/mStpK4vsvFUk
C4OYHEgv4tNU4xq/W86Pejt9auR/obZynLc5IcOWAoPZ7MhXBQ4FDhbcBHrx01ktGDAFhTRiuKxF
KK7OX+l63SA3WDihVltow9iU8CqV7dlVqMwU5Y4/CDKuUa42DhD6QJQgv6qculSZN9Q1HPoZXA/T
LqOU2byNW2VJOYMtHvFbOS1cnpIBTq7Rjew8mqFlXL3hvbLHIB/Py8RHd/1fWvJB5nCkaSasX7HS
BmkG7GbIf3pnxfubvdIWcAGXlf8u+qcuRRDV1CzNVRGSQnQY/Dz6QVKiu4hckJNMkimB8QMQgYZk
+vSarGv2F4Nucz6t/ivNtCd3bXK/9+AaUg9Vw0PE2a0YxI/8oLKrByqg1P/i2Yc42w27JzLSxcf7
A2jmuye4vbrLRujY6JXl8gbFNW6b9f83rKP4obkn1/tM+ITkD/oMvcc6AGppcQlPmf3fEnF4CJCd
IiPUCTqoD+LKF4fsSnwBEF0BLqUOH+eN2Ny2iRFFoVnSygVfGnzCFgqc9DwrPeBaJYBvJj+NTdz/
YADRY73yxmjNowFUlpb0uA9CFvbZL0+utFrVKkvsv+MnxS/NNogRp1MniAhcf8RVlBli+GXk7vfK
17ZXXjbmRC/rSphrIgsVPlo8KC2Ph6bwZwz1QrFoBmxT61hxwmCgBtRIb/MKkLTt2oKP3FWdYLtQ
8zHJe91vAoVhc7c2TqlrnBkIElshfltvSKZ99EbQspG6NktDhH4WJbRpXCceTel0xC0IRBzVwK/1
628zuK33Ruthh+LX6AxR3tEetODTbQVm7vw5KA4m/6cW5LOMK7qBlyxrruQ903/Xp0JeP+sv+n0k
Vz2bT8NC/7bTVQ0RlyA7ZEP8DyLs2VlSXMFaY+2zxQqybphZFuhJy7nCYHF5oCeRpzhXZGYZ3iUQ
6Q2S7WIQmcvTZv5kTbJgcAWW3F37XY+NXuAcHqak84RjwUtHvmr25+tg3bMjs8JHWXfZcyV2Dgxe
+xxD1hT/f8tybwUSP7LOMd3eUhO5NCWSkziHM8qpZ+k4dAwU16L+JQsrPplUz2pf9BjvQpLdcuyg
aAHdXhKmH/JBtN5g9J21X8rrChu5ChUdQN2EL+aO77J8NTtj19yi25v4zuy7xL8sbDAX48OrkNeo
xsy/u+3222QoPVJNUkmQVhv3+fH3092yNcmky1rpboxx8aArw2EBgI7UoqioxvhCVkCexe4I1RAh
PK8xAOuIb+yYh1VrR3C2zrv+06lo1dBXMFTSmss/kLhs83v/03kTCMV/vkjKOmE1Ji+EqFebndTH
+/4RLwN8pxx8Y7dhvw/HAWy04ZdqnYDQ0fHYOCJVquziQ+kvqV9DztzZD4TE9+bhDTOE/4N2ALb3
qoZB66mkOW1CmQTCpeZb286xijRVTQ5Wp+MNglCKkeGMwoojl6aEKN6COxfk+KZgnTNPTM+xVMnO
rQPco1uh55FobjgEcMbtLA9fWwq6SeTE611dNMbSX7paeGJWLTz1tbd1T2cfZLfk1Qy7AnM4lwZ2
oxrJYPs7efAcO/P5NXMM45bHvflW/XEqlndYDdRrSYETYLv1fmIsiVLKL5Zhwzyn+MGNmtCAHvqc
80IGdmO9ex9z3JErgbcEQQjYCdZ8aGq76eXp5lLkK0/9fi6hMM4+FkagvmSQNmy6gqJSrr4ZUn/g
hzWhW029T1SaSedfh4i7SKL79Ycmj2QqJmf5HQPEmBhzezBGMaRC+NepIikNiyjhUV/eOQrQw/58
xjh6n+IQ+aJgHTv9/yjL/QuijgQbooKewQsEFvGhSGFMOdXcBd4zExsLfuSODhy5gmEni++pr1xV
rMcYl/cO8cLXUuomO9z30z0zTFoHVmrxOhBaAmD4ZC62rq4PbymQ1/A07X+KOswkQitUhCnADjI+
OSgCMXa1pnzaw3sbcitpjF6lVdYi+UwBeW87Zl8NQCR56INB3zr5b70qYUKc9MnUQlMzciohe1ix
iPFBV4SSTaXJC7p4xmwofBMEVR71IoOH8ESFKLHfxLSFF3/CCIOXnNeLwpQwsbfj+6kXoBWCq1Ag
1Zr/Vztd9vY8PrHAtE9XMew0BakowgyFzbRWWgdDMRGpVpNQMvM9QwoMDX8juMOdnk336dli9Psk
PSCwHKdbHbtIa7+u+8VvJJqoPzxVHwxZDZ/jTF4XHYIS/TMiFAnO1u/6OxlAPrWquLAPXJcuWI64
s8NgHueR7ub7K1NQeNemNPE8QxMduoQ0Rv2rfFeX2E9Rn1rFgKvsUYjiHXwlST2RQ+3oJeUNHk69
wDjcCT1yoOWfA/HMjYdy1hu7rJ/jijr5Hah+QElY+2aNdG14o95nmcjFfCZt0+Zut2M74+sgmG90
7sfTQxZtAFlsvx8otdzvJU0kPF591uUnpjRxIGd/B9Yvq/2y81ftTbcykiauomOR+NBfzYpJfNOA
i0sDMksqVpQItPwoH/OBTF5g2Hghx3kbxZoh4AZ1kPNrZudynNxh1YVRC+rf8pmUroIcMxkVdKCR
dAAsF6jZ7kZcThSjs/UqLza5G8Jc4O6FVH6XibYdmcxk9H+dKf2hpsArbaqTy4OIq9faAy6R7G5H
rNY715rIpwGvPGmKCSwseq/1D2EB3W5H4Yq1rHakwI1MA6EV6nl3givyAYsyEQkvd6tDsCQLkpL3
+SC+uCbvNoF+B/M7eWICcKPrRW8CXEiK95rtgqGK0lO+K9TixrrSncQhtGRxZAkizn6ITW8R54i7
QJCqgI3rctUOYiuhh1MeXDMIE2d6Mz0Vc9JZZN1/C20J48/V6kmE8dB3yN8hHXfOdRfRu83rNOwY
347nG+BJCT7Xsx4Jpx5q+m8F5060hskyP13fr4ZxCP3MXEJGO0g38jmKmheplQvmC7S9TQu2Z4hd
8vvBpQNRMHYSKH3ZCi1ZnPd3q3APRI0YjJnCLDiPzfh50U6ZZCZchptwe1rxhfgAE3ynae2F9rvr
IsB7lG+sAl05rJLaJm8q+89OFSj68IkZvyaxwCfMxhAHHqiG/lm5wHYHQA6rpgODmyWxJVxpbf8x
MX9/cSiuuRHcgITBjH3pR/onsW/fnRKFkj3xWpTFH3zdsHQAgZk5oX/PUthJMYpgUqGloEGdi4pG
vxcQPqOQi7fVl2dRw95/wM842iR6YE5caLQLsBLAa8hTzhrlRS1n2TMRegM08MleeYOr5Hl58J6N
KGoTdKKeUA1wLJ9EqWv7gz+7cK86O22ySOb+lRVoFosuzIcd4ximNxarFKzwzWQ8iU0HzQTrmEZb
J1n08XXuomHkcszn97dlHC2LB0rPsMpX98rjgdegD6/RvVp9M0P088PtZSA9wZIn+XEv1HSHtf6/
LRaeqvt5W/E9eKDvvcGFKde+u+lvDFW0zfhNEvYAtoBvTxgjUzNm0cE6q6SJDSevWZuFKFDJxZOb
bBOj4xHn3y6Lzn8GcD0EReCX+1wlZEN67ZpVEENM/a/zZSHg8txzK1Ey3GLDPqF5thyX4sjYEXH6
1q7d/cybKHVJT3E6kvQ/Zt5G+4K4cXf8EDskNV0S1ZgYbtAdtMWBDgmUiiRCMgQ3zn/OShA0Gk+5
FeHhRQu0vfmgBCMWWryrHiqrJftHukxUI6Rjn0WiHQnd0j1i2Qf3pLHuqcFKZZXDbnSmRDCMAdN1
Te0j5U9U9hgE64Pvr2FajSOh0UL7b74VfghTPsKZ6dTdSbz94IRe3KSMAZsfaGaz80KyjceM8+Pb
lnmqZhGx7BgquUI6lkruY5UD5pSJgilCS2wvlK9bEW0jNhDh8pMZHQqVeTqfCatxi+lsNX/iVDlK
rZ0n50evmHQsiSHimzSuZEo54UtZdL78GFCim+tii4qYZF0Y+748bjWdKjyVGS5TaXcqV46v5Lel
/7XavTfuvuszHVozyQjZhWvE6FupCoP5tGdhqoOfMwTnP5b+y0yhFKy3LG5yprK01+fxy1GJQZVt
lp9Cg560j+p1wsJbbJtsh6apXo9+gptzO63p3ttxiCI5Wakdd0D5iXcdJSvmobCPmFlFqbVfXvVU
6Q2B41VCHs7c+ccdYDOJsaLRzyErfvuEPLWDSDC70PYihHdaOhW+efVR/87x2nY9cL2O+J+ouBoX
y/Wve0NLOKm5hadyGoxtDtCrp+w2SbrICNII9f7qoEWS49dBR2d6fxnXuK4TW306szbCwZgKh7MR
qUp+bZwSGHD4FZewuY5bv1mlbGxgB9EBtDEh9IH6vqv2NPe2fP0MGPhloSmEMipFZc5YcYzFC6Ew
jKIFsfVxGP0xoyjOTlJntbLJMojCrGzSEHhxIkiH8Rn34Zbf3N4Nqae7TLFObz5ab/Rx5Nx2O/ev
+Ox2/sfxxYrpcUVvJ6P/kppF2Zk4/Ebdw2XwlFOoB1sXHatLj1xZleAVhvdy1yXuYwEQ7LWX5C60
Zznl84S0HnP4I/wAL8K1pIT09Z29C7V1cIlSdTDq7ZVttG3aVz8bHmZPa9aScWy/tMkOKMKnEjX6
sU1bryafjU88UOBzNeuh7ouep+nA9KWBEJwCClOx1RS6q/9OZzEx2jxmbwtkznkesHo/kRF36FMC
7WGzktaCNm68vj43I6rOCNw76Mb7sgetxmYfiwcyoqZRYYQHPE9lYtTsq01IpAajoQVDYweSYGf7
6sVm6u8bjrp15RyRBH8JvVPH0MEnKVaPEVrgy6Zuh71a8Hvqa2JwVEudyLYbawIr/1E51O+EBJuI
q4/BJlnNF7KnZ/EI5Dq19rhTVTbP1Ii/CAObiIOyGPZBHJ1vlXuqXU+g2JfpnM3BP2b2CI2moqvb
3d3ta3+JB6+iHnNFkR9hGoU8B9ZDbISVZeMKdHpjmws4JqZ4XcjecRuBnEkNjJS1NItIxdf08HLu
CW3AL2XyOzLvqBZu37MGuyOzC3KZxkplewd6K0yBF3XCYYyF2xzxdi20k6nGfd3x68NvJZcG0n5n
c9iQmkXL52Vyw2RvWqV9dYefeefJim0/GSSvvKkcuFZu3J0hEXgkf7SudlGlxmYLItNIF33a+MyM
AQ5a9/mWfIFyoxrvJJdkUQcjHnAPumrsCDBAZlklKhPKM1jd+Sja83I4gRq2MBTnORDoRfIvxH31
tkXTmRHoPV/S8D3W2lXzNtThqnh8TU+3w26u/SoRL4+ob77nTtuL6jI9NK8rxNkFcvdRi4HG6ovU
ktDBRjEqwuO8gNbs8TaWghyGRXIazAT7MZ3147h2G+/mP+vBJHfJKkxP2tIJ2CuCnGN8Hexg4ZOV
dtqnDEJcyyQs93clMGSpZty0KlKGZ8ZexfpXu/uajP1f85Z81ZTkjKvurjmF+kmpW8Xb+Udthe+f
z1Mm2Qovj1eEoN0wx+/BWAEKqjig7d53GgU5UR6Q2/9OSnFQSR+bMplwVpitYK6MFChDHXsrP62S
YVtOPtQf7JKAuPqF0BsjQuQM3Ur0iCQDyDVXdtJOwnKAog+Ce40i6iuVOtfv0NHOtWaF3FzQvQo8
plq0pdZlj/RdmCqeV9LUrPmFUCa8Zu3enEWxeJQ/P+zVcmCyG/faFYfnUCRIMlr6FBF32LuoX1jv
garXfpOx1r+uR3sS4YZ+omhrdOatSPM0ZwsvTge0urvJ+/5IlIFTqijHB3Lor+v0KLHw0Aw+Aiur
KkxJwuHIAlwDHmW6Gw/DZtszLgpVWJMSWko75tRgt9sR1Rw9535H0J+oXKhUZy167MNlGUwY9bAo
ydIWQyC8R9rd1AFE3ceMwwO7O3aDY+13aS+zI45+S6GwDH4hNjpjPtESZvCWyi3DAMsjsNNCHqpw
zPfllT4EnBO7ycnxOBI9EuMlQ1RjWuzHyKaT3gEy/E7EMHAWuSvsykPtTqGnkO4bTfku3FEdOzgq
pvqhXop8yA81W3pKIXXaOgMRGKRvc9IrjyaXJ6GPsoMHJlX6ZypeiK4z8R4tOR84OpG0dEAJohJg
Exo8tm5BHSF18xnsNzUAqIXnHPkjeAPyzwXC3HN1dIiJCHPze/lUkB5QFyda7Nlem1uJ3c0wqhzP
qay4aSZUOR1V4yrJZsSDDp7TMi32CCW3SGFOc0TYXL1rZtPHU1P2liql0AbIvuKpxPbm5Ls/052v
rCDshckpXEzEMCef9X9lSzZirmTqmZV5zZ9DnUr6LiHl1Uq8O2JfCMj1KpyyAY63tLiih6HbUYAA
Z8aB3CsWwXiZLjDlzNYGCcDzE1ZlTvQaXRNx/Ya1WFQhKw4kmScxRrGdDeYDjEV5ouiGKOzUNHBC
U3i1E9MCuzAXI+EHTg9Mq7z5KHSk2qGEax8sqeOW9uJsyh6rNEbz9hmFVQQL86N7lM3Bu9N/Jioj
+1potb8AIjMKrVsCeGYqemVSAXHrbDQIlRQ72zNhxLV4zYGfUKXw5fDxA7849gfmtT8xMaPOlMmY
31v8Wa0JMTZFLrtJZUp1Kkdaz1xRxecsdH92j7WHVFJpKsTWu1/pIAsoacoARqbhE6rKY9aMPFXT
gsDT/kt8/7TAZCivWfnvi6Sh21WMAvD2+YeFbnF722HB5/mv85idQ51JlOYm6s3qt0zFEdAO8s34
wMn/Fl890aUYoLhO5AbPZg1U2MHzn5VUZkwI0sbJt0RKEwzhsWhx+E7RXq5F57MSBoaIbK4oLEbv
zUI06pDCSraBYu5rUQebT6PjBywVIjrr0jzwyQ5kLJ7thahlwr7sQW7ZDowzYZXOcsSwnHSFXLTy
deR2jKQiyBor3psO7P7nQBPxPFe4H7cGnYb1mX9MNoR8+XJIqFgKeGLfN3J+ht1bjWxPKawdY9Hs
MD3L1AkSurtkCadWoruxPV0odnopaQSSsmMYqBxVusR1vnTezydlTgexlCT83L14bLNlGEg0ocDs
QpnS60O1AICZuKBAEEHseSwhONoWqf+9JE2VlOti+EUXkzLDp4RLuTY6XnQr2gwZDCxiid2Luo9Z
64xWjzruNs9uKj25Ja6kcynvLP557X22Gowx8hHHrHJy+19nsUx2mezE8lKdL2XzWSCrXNJDrizy
uC/zIldQj+vo9Zg+83rNPBaKiMYXbjOlyGw0QHWGoG7xryfoSV9JLBBTIH416lo6dGD2/Axw1TxS
L1Zm5kgX67jKcuIecsyhWfrPdkSXJFp5d8XKY/TpPWqT1Y1N7168tLaaBIgzn1FpuwjaMoR2mMQi
LqEBZdGUM8awjs+VpMxUzECE37CYTcVf0w/DITYRretOAh0xO3UD4YyoDH2ysIQIsIMSshpidY7L
ED2AueqWPavFROEwzk3FlbNGfJ0DYxgwi35RnBoG+r0iaIAzpwHlpD7YjI8zoengR0fngCR4bCHQ
qt7M3Y+tsJz47S91sfPHeMcKWxIA6cUcETDEaPbkZwpmLwc7bh4Q5no4lyNeck4fzKabIoVKiE5Z
uxoeIIigBQF5ZqthvaERFcdTD3U2JsMNgwDDVpctdHg8TcQFv910ltL1SLRPXPaD4EJUJFUvxnt3
ZTpr3znTtZz+BHJnqDurd92cX9tovlrC/UJN6slUcuYJHraGW46U1/6XuWrgtu6zzMPgOkBxNfpN
xv+JOnxHOPhvLjdcVlYO2Gz/qtEieQrJ7W3t7z4VUVQuuA6MMUckURZL0FnlzGWdt9oi5x9i2pwu
jPQbqhBvxJETKEYm8zUNH3MUq1TC1/yVedMAsnWuUo11ZwYL9g+t+Kc4lXjfh+Pqksa0L77ksWA4
NYtc+F+BfrlA7/eUPonH/IOmAS/VDvJgjVceqOBDj9JLGeJAw6rj5MeSyWhcmddq/Ei8epl7pw7p
16sKuzYJSK9JrJVMkImwOsZi2AIMrImfovO8p9U+4zVPZYKUoXpsJW/laxJujTCxcSUqPYVe7OEy
NpeTbZdf2eMacid8gp4yEWIM4WtqJF7/PYq+UbMEfKs2E+/jwQBR0TXjveXIxj3j8ol1daNfC7lj
rTg89eVzUIiBvpqhyJUyWsg7XBFolybS1CI71khdyVIHTfUXHmiWq4Mm+tX2i28hJSEnK+kwfpaz
j6KCNYlkfJ48qcGR2kkbMyFpuexYeTvohZsu0C+r/5mP4WunD1Q/9gpylafpnTFuRg2TNBHnKLwv
rPI2G+7G4BEt2qA8eBs2r21SaTUYYV3C+CQqVu6f5hp0UF2Ee5pCw2goLCgi+m9p0cDcbX6zOzTc
5hPU5gje1WGhcjNdoeAl/dLGjorc0+47nGOcwTs8pSemjBzvG5oINKXekbRh6dW1oIOsanvZYdQs
dKpkQyFPRC39koh6jofxvQiLZAxjB1FkOwgxf1aaxC1/bJYXTYkNIrKFQxd7ZFmX4twdOLplSxu5
mMDT2BrXNMlNmBClxDzbvF0lmc8AH3S1z+oJlS54PmPJTITqgRRaArU8xpempAsqAOgONkMfU0z5
NfqdkWPHL/v2hOpuiI3hkkH8zN8Ka8x8zz/eHMdyCFOvXUZ2qPUllCJYlFpNmzpS43A543aosp0g
Av8Ele1xKllb4i0rJfXFwBD+91M6x8eYTlBQhDKGQk3NSHy1U3UCoLgfcUXmLOBYfq3PxhCVRxos
YgJoccjsSXT/LWRbXQ/xrI062r20TW0g8BoyBk/gbtwr21vNI9bS12UHQApxOah2P7adPHyv7M9A
KgkwPK1OVRZDGW3ap8PrbZ/TvTketOdEiCUsfNQfR0Wkgb+Ol9jI9fhQPUI3p7hyPd7JUpOnW59R
JXCkY6F4D8nIvdl+WGQ9bebHwtGJKLP1D92B/KLgGsFIzInKlZgCapDDUQSQNZQXVVpFotjbTqg8
p1uplQZu89hl9aXVuy3o3OAp6ghKowaKyGWhIuEHEIv39O6WR09wrg/FNHZGAff3Yf1qmZTkB10S
/lz63ELA6YXfhVVe80EwY0yPInrjOodKGykWrFioKveXvAKjK1iYrz0gdWAKnfKIHtljx+OZW0x8
Uw0YuVfQIVaL0VZkr+4hhSRadPYke6BuHaUU4NFchfzXJCl/0TUZcnEmFqmz7j5VWCk6ofJsxPOn
goQWLH9e+ztMvvvkvgE7V6VIGtkF+aQrrIFlOCblCoBM5/mXd4P+sxPgiIMR7S1A6ctQBNbu1QuS
XSVDf/pKpVLJBtQ8VHGU5O7CsLtsLmnXy3o3GVHnHZzWEFMIvUyWjH2ekNRsIkLDb3vno/EwkpCj
9Db6HvZ5cUCJXF/OCBnx8LIvvzYrQh0D42O70BOSW4ASj+o8yAAILJgV+bOnPX7UOWN//xvSfL43
6/owYLqQ1WrNLn8GUcIEEw9uS99Xqiqfuo26peZ4FGvfOdtV/hy7ng0fT1fbyNfCB2Xt8Xz1F4d6
wpECHHzNbnIthXfJ0mfBn8GHONiaU57jzmmppvistojwocEaljOBywZ+qPJwiooN2gm5+sFFCDaY
RUFSPzlG8BhqEj4mz0Gt8VuvvOVyWBBMfjFLov1YwgKk3iCNIw8NWMUU8pGqe3Vs2mqpfWHp97Z5
yd8zOKoZenPy5mtgH8E7/Z7CMbTkqhnLbnXLB0aSSJCWAZb+1Lstjilpawt38zfv99Qhn0KHZLqc
qWR9tWFYLy3vpSKKI+LeFGM/x02iPsu4Qj+gJER/zPNZmem6tmvgBHS0hvpNJ8A734IS1MO6xWmS
smr/76J5ZXxHbTJEVv9X6tCTZZRh+16B2WJBxSXjt3DuLtqSLhbeD5QVzZV20Ghk0Afa/DFUyKG2
HEaaKhljLQMu2k9YIz8Cvy3P3dcteUglmnTVF6ml7sKiQPzVlRe6M+RnvkR7GVk680W6Sd4A3hTL
FfmnNaOOE35io81OoIqxC23FyfjT+5ErcT2KQ4DKWEufRaiIjC9MMjlyuL3EeX9qjMdPaMMb+zyl
r6VT12dhMOOryQmtRfJu+3LjkwDZeFsG+8Tg2tZmx+DMg7aUNdAuYXUm/Mz+6SRqDybIgpUkJze0
u+uvq6pRDDFaASCKPIjjtbBs+bWROtb9mpaAypD7RRgEwRjhN5WXKp/KkdwlCGtgBw4lR0Z+32WA
nhd9SGyeQaq/Vm/xGFucQimWuN69/6pe8nHYQStubGrzmKiO17Ou81dsQSliEv3EnuqlMywoLwGn
WExEdocHUSpCwfV9lXrMzVEiu0ZKfLNk3zJ1GHQRKz6wugtAh7Am2NL91xXhiECaTHxdG5NOSDZ5
rtDZDPIlWdDVRQwkVzkFgsB1Eq02eR2uxp9q21WbmpVh6nAbDLg5IQ4gYCqF2xLMEWSs/OWvh/ig
aWkgcpNa4+tdjamz7mZZwHLWThc9XzT/vMYdJgtMOEBQFLl3rgKBAPBZNcJmmQHd3D0o7/MKmaje
F/iRfJrpHf6lgg2Dcj2PoBCfoiJVopkx/wolhNSvcvbr0qKjH2bpea579qkGqYXz5hGrhrfjkiJD
rMkSt31ICNV0qgXU6yrWhQJBLhfPxb+7PH6Jfz3myJRMRgs92P4NgPCFbjU2LPlCgOnzrNfXH77Y
RKJEAMKh8lBNEjhBUvTxIl2D9j8Z64QBqq+j44VvlKpp8dQK7bF60cvn+ry//AW1vS8xmQu5qYou
fio2Dkxj27bqrgnxxmxRTsmuiueApn6tbXYwmR/HISkGhGy/E2QD+Tc7W2voHBiipPLDoPjNyGns
XCVIyAkcSnsXU3RrSdSRHVQNO5RgGv5ao7GPU7NmobwBZebyjcWs2QfUegSpZJPHD/76MskwfSvt
jqrXfOFJTr1WsJqp7AAJfvJuqZk7dMopQk7JhmkKTVyD++EphUN28Z2/IHJGqt1g0ijkFENlR7CS
zr+in/98/65MWfSD5DqgrKKqB0lqzaDLCiAWMrRPiJqe4bAkz1A3SvaRbr5JN1EsPL9/4z6ebP13
aexrBBSsZreRuN5NcfBV/+Gs9bH1sOvvREtDE4IkRmzFXl4xuJsQ1dejfipLBOZ7mmUlcKrqhiZ1
lwanA7+K6hgOrkMoM7xMGVg2Y73BWdCdRLEbhoq6pyF1rzdlzDqGNdjTodIE6kT8mM9maOZEwHPg
u/k4b4Kn0BSLYsfD7rKOhJFxxbGED89VL2PVp4OX5SDEBrOt5MiMd171My81JCE6o7Wo5+dBpOB6
ca4poMmcBuDrRaVJA92bw5KgtYxBtpoSXbapfJQX7EWpHh+kkrYXxHU/QsFiuL47MOLmpoHTP3Ao
bPVwi5H1CPZEFh7NEt9L7+N+Wap9WsYfDUwwIsYFnEa1fEAuu+zlY0NdYPMcBWC/mh82mcG20mB5
Qs5BOJDSHrFaqE3nDDueS0bKc3HQ0N6Ncd6MSBx9oIdRIsIPUinsiDQpzMoFP5DG8ZtzA7iS6HAw
kmgAqyEdA1GLHK3wmzZngN8YQJr5DmnQC3zn/7lZzIYlcaP+oNWFJmbd65/5x0iy37h97KW4fCQ/
QVCIQlHFq1m9O1W/A0Wz0r33FYWHhSq2Krp+7L6q1CQTgFdSnx0w4q5tIe+aObaKziBPEeuB8Cht
5S21EpvfFDBpCFpRpyYXzPkZESLpyjV4RnMTC1jj2g6PQTFeSJHYFrWbUgeQrOx8P2aBWOBswfaw
5Q/BnHlZFufidH0PTRK8gLQPXOZn0J0nJqig696JSQoBglo/AOVa7b9r12f3XvsecGIVoo9j9S+T
0Z19AC23QDCo5TJRCHjVATs31wjlXxwua+V1BB27hTkdtVAJ43BaDPZrvaO8nWV25eTc2W7fX9aN
7FXUjBaWnD4P7tOGbcu92L92PIcQmaAZ1Eyjo3D2fcou2RU+i9zYBl+iOcpslnwZnmuko9WMgNm7
FBH1nK7C9C/qKtWeA6+9C5HXBWR4Yr9s77TwsKlN01mrmabPZDs4TcZFhzTri513qwCAAfAI/JXB
cGKeCklT6tIklEiU/vj2srE1PcWlbsG5/aVAYXPYrU7/KMoIzDj+nvB/n1EOLFtkjmSN7HhmBJLV
vmKBhPK9qzw2HS+pq3hWwu75V+1ps0rkKZqQyYrvGW1Ih9bCtY+5cM7CKPPH1bm48t2gNnutR17n
OFR3nSougf6rb/ali97aQFYDKesbXwRhVjKkdIQeEpZETSRob4NihABWdJ2JjyU+6mjzlV4dXn6m
A8VDJq4qQqECdv6GdPkOSrepPSuFJR2ImfYBlYB0Pp99EjMewoowQfluJlmFniZVawl59nCEfwR6
cSw6WcEb2Zbm8STLnfnlySMuyRF4RXqcDYtDcwrEs6e24Sek+FmIVvCAIPpUJZothoPEV+guZvaU
hDYfr8g3t55Pq0E0j2vCsXwNjLrvMDqUuNopkl60hQcs4Wr3PISB3p6dgbPPr6W9xH8xN5zn/Y6X
kLtAKstbsA5/iAz2uHV+QrUDtdpcj/XGnoZDXyOrvC47FmYYxVtbSTfh+/cBvpJIHvi3eKggRjTX
e8kCENmTsQURYgFNrrPIjqJ97yVpIvF9wmpI5/KW6y+95vIWiCUrAB+6mvaeAqdhm3n7PHMl2Z67
Qk9uPzRUbqOk0FkfrB9NIhpFSew5V28W4l2zXKEUbO4GKiB/jgmZoefwMwNhH/n3OmIR/hnkMUWy
SmOuZ1mrS6W0pMRAZxFKQ4333OV5r7/am1qEcebl+hWIlXYeFYk4h13H41j0XRow4ResxdDrwYay
4qYfMvnrFFZjbkYUAplFCoQtzhljeah2+zdRQPDa8ANlC5QOCuDFLSQKX6JRxOP6X+BMSGJyHey9
qUuHQ13jVwRIW8LHlvZDqxlUFyKmHQ4yMQSx0z91XxSUfRJVrLEyVPFTR8KM48cRjFIP3j0SuRvP
DvB+zDp0JZMvz4eJwQlMLyHTsRciP1rZl1UAbxkhxra4vTyzVgCj5qrSqGXL32AXTzZUvZDx5tab
PyYhqzNKFXT0YnEeiy/atme0iyrXzsVq8XHHcohVeQZD6Pn3Xdxjlcnk6vdnC15CJhuDQpasBEN8
3fWuS0oaclNqV3jG+ndAqBqKwP9LU05ctm6AdCfJEcmOjwN1IWASIu8330LQEWu4hEixA9gcP8Fq
t34ajMVz9M9zkti2pYJ6n/4Kx3p7CR8btqDcGIIV+3PtYX8hUtsfg4spZnGgDmW4BJszmVsef+6J
btpmzjJnIgbdfolDu4rPVa1dRsGLUzlSd1hEeXg1M6S+tW+vhX6uUNsU167RxQfTXKCarFHQlMEo
pPmahy73bCaBAWuOzKc6z/riHiI0YuceELDVVPLwzv2RIpIAlRtyVxt4brrKEj/1cxcyk7e05p4X
1XBeeZJmZ+qeNR10iaNN9CM8hK5YI09zr9S6ISaA+1lwEAn7esL80fgCqBJNmTSaSPrHFMzoKiP9
UZgogv2v4mziqskM0VCpKbdOWYrxiWmmWscA/KsigGPYJnakneP56+utfKb6fKtEmYjabLiEbhwX
EGk/naBoTnSeF+h3YmucTYTHApWuvfKAp3l1SiuVcqg1/kBFboAmc+98BLE2Ta/zk7ABsuywrO/a
VVz8nGQGyak9aYMl3KOgKzaFpSm9Sp+vlBGuXCFzZ5Zb0k3Z1G1JziE8HFY7FeQct1233eCtpAT7
5szwnXR4dCL5tdcLiPukba8qg/l1HzBVWx/7oxphZf0FcQ6DHLJ8zf9P0shz4vmbVfewSIgSJ4AT
ThjRNB/S8jdqfZ25vuE3dKjOipfyFuXaLJMTzdm+wt0kY2ZaKdlQZPrE46K6rZRdzyToIwfBzV9X
C5LabSdoBM2k2kjPrKTwjQjZBpnxk9c7NpuMGBGMpcTv3IpNDj3HvE+nJaU4mpWyEWEDmJmn8uFE
kaZv/VAp2m9w6/6d7D/iuR3tCP9fiKR75W6hd3dX4XSxH0pTau9r/zdtjyvTL6mGqCBJhNVzwu3Q
pb2AxxtPUmXY1Jwd/QJ0GIcsD9gxEHSDJPzz8Br1CQatkBN5y4ilO8qEyNV1xw9/1fTJ+2Ol3G7Y
bZsayOF9PIYPk4yPH+MYr2WcUCXoxtvjB5k9dEkqapUyJHmlquexry3a8Lva7iwoPe0iv+d8dspb
0ohwPpL6nABJv8kPJr8Uwh7QtsFQ1WNFYW7H/jdF61nImH4BmIw/77Nvw6iZkq6fM8yUj6cgDnjL
Q10KwQMYlIByKaJenl7pOjx87wIFZ5haF7kTtvcI1MOeOGIwD7zZFEaikjQPy1lpB56GVZkNIquC
nK/L8a96VQEXMkkVOMxx/dQlr6rysHGzooRC8mTROveutv5OIOJhC88Lp+gjJQcQhyqG5OQQddAu
YS/Tw7wiZXSw3Z9/UBV2WcDJaO0v1j4Fy6iawGnc+fGevRX2+zQz3Kr3GVWrxbb9x5RWzd0JB6+7
GtVh81i0frTDjRpug626/bxzDr7EB198YW436Q2tDwYXbv2jahRCiR9vbS7KWZRTfKF+g0FS+WVR
WmBjj5A3W9aGGBbQvpIn+XYJjO4rQgwewXunGF17R+2OUMadzEyG6iuM0G6AabgbVxbYXbK4Y7NF
HtyhzS9IP5dm5ehCZrIvcM8dICpnoASTeQdQCd/BiAIPbIjZc/YoFnce/sK1jjO4lzQTKIbCsPIl
sN7FR9G+iFlq+WV78D2+4mSra5toLi+Q5QuixmiifoFnLoaEGK30dOn8SQmYs6xYVEWHK4MaoXjD
b51YuLMyK2oKGX0sET64ZiB+VF/VxLvdBFWqOg0uxU0jQJb/zcFJF9jg/BsbWX1CyaVD/xkU97jb
EeR+qbnQqcSWy2ZYiMTO/cI6Q2DSihUn+9MwCWaR++yR5lfk64SY9XpFIF1+rT+5lJ8DLa74kCsR
oZOYblLhZCP78HU/pfKjc2OGf0XrB+E0IA5t7ptug/x3a//9aybhmGtpe9MdGuQofFgaThu2XXtt
v3FX66SpqAv+l5zniZXgo80yw5U9Q2b9LIUtU9Lkh3qgFlsLrvKeVKiddGTiZTvfOLIOIixe67RO
DSHJy+N05sX4l9MMDxO2bcSrFfSab5OZkOSOlqQJb7HuwG6Ys2S1ajUGRV91OobS9RNA0Jr927Jg
wcd1s4lU95fpgQNTBvUFpR5hH1baLBiodT5FrfGxyNrD0Kj09wlRPwUQt8OeczcYMvnB1T1lqCR+
GnV4ArLcbrdsUs7nC+tiCbBypvdrmUaVFJrWa9uN9QRSqjtZheGHJ/8GouEkeIuf9nvLBoCq8ju0
V2/8Kzy12wT5MCNmTsEMYfjOXNdW+HvBuvWFZvtm8G4woOBLFcgT8ks65i8pfyBxeVCRa0CPTbsl
/33U6s39t9D4k7aYx667olKaGA4nbQxlpgOICmCkqnjVehj4TpEKcAZJaq/7XF6ngLVe6cVoVfkQ
TtLgN1gXZy7zvGdCcwnf0QztO65vLcWyBhkAT9MEwSibOEAvNIFdYbRNxX+tSW9mTGG+8sGhZjp9
7Q0F4oJCVYszz/IvnDDphjBUlbUBc3R2A8vGasgvQWUwhf5d8Wztot2dcCxcPIfi7YG6PV1v0L5g
SKEIxKkQfJ/osNoZoAiw3hrt24YTeer9dc3WQdwZRoDTwiZKV/PCxNySjXpNnsgveiWBc8Tf0IjF
BS7nZ0unIyyM7sXe7BlARA+LT+KRDAxpblUPgZX92V/31dbSADplSftpMU8fBtc2iTiS7OknclJV
/8Iz3OeWucUI3aQxUvSVYUXrGO/45on+K9JFtgWL4Ct5UmyUaXiwY/slpZThuyKiH/1aXaerhXBd
ElInn2GBFI7KEvUV15iB/ypayE498WFmXV4ag6r3EVIuztgMLSmeWo0u5h4lLuXQ8cBHVOtO63Hl
DjJ22NjKxOlMh+NQgLhUgKc0p8Os4Oi0Bi/MjO7h5QRa7/Umu5r5SQc99nI82FJLL38xHit0+2lP
roLHMZhhp+fr5oMk1z1QZF5bMfmZruBd2wOvl5/3m+zr1NX+CvPVCS2LOd5ywMpLglMlb6IanN0f
n0cAyArY3kHpEVE2gRcbHRs4n9hSeEkXjqDIlMY/7tTeVe34HdtGfEAbdejZ9Wd6J52g4kIvtoEe
wYOlI2bVmP9kdw65Kp+lNvdu+cINovA4gKOhMnOxksi0Qs12uLALasI9Gpf3OaaLPPLY5jdIezhb
/3OMtEAdmUNFO0Nwf46qwQgt7GRCxoGYr4Cc6lXB0bzVTTYeJQrdoa5+OLDL3DGtMNLuCyktduoL
2ehm0ni45NMY9BLf6sg5MTF1NFui8TINd6YEk3KslFg9ZfK7OlEJwatXM8qPeTNp7W4AjlsQwIZI
jlI4hGECizdg5EhfCvGeeoU1HPuii7txgpcW8V3bBou24w3CFtVFG2oNihqqZfg9brvvirfBjEK5
kna7z2onMTdKiBYB1rdrdnbVAv1ctRxTzLlLrqI9Zb26QZLp6aONBBOfQzcMA9Md+X52jat2+wPI
RgxXq86CIJXweVB1DnhTkJJlHVScuY9wqesyto7K+f9knSn9lsNHXCi7skAHPLGTPNIrgcSrE30a
oD2uADW3dalmib7sz6vJQGb72JsaxReDVkygo7vg4c0DleS/vQezq37LNxZcGLdWwQXTj72H9kgp
dJBEbalA6/SpMbwg1Nk3w/T7pfpCJmSgvupsAj9emaQ/Jm+HEl/WUBXu3VYSPNTV7hmdjHe4xsSl
NJi4LRE7epuXHLq76lQP2UBI3a+koqGMm0vEqPs0/UTGoBj+nKo8O2bUTaiM2bi2T0tHKMdTidhB
8ovYNsyS21Q87EAUetZLZJg01Lq92Kjlqf3Q7ujCIgyMpICtXe4GWdDUlOGlG2jsuB/3+Zo9hbM4
6RP7WFtJQw7TlUirZZasZBB1+KC2Eqg1MyFrS2iDNmRIXAOuq41kIQW37Nhdfb7konj/sLYFQcIE
9O4vXwZuw3F8t2r1C0jCrmodHhpiv5HFpJfgYO+/xczoXiaGYDXnqXHCTE408DGywv8XdonxKK3L
0ZVy3O+D1C1QGjPbu050Vt+Bu/Snx7vqzZXPOGC2QpqVuKb56G0iZ4ytYAQj6JUUIcJH7aA4ifSS
KjiGTX8GHFFtSJavyFhIi9+nOFiZpVX2/fVV8zyU4jQZGUVUVYkZdrCMSGAcRyuUc/U9fkGC3UUY
z/tPPmkscBH15TwUHFD6+wJaVCkCxVZIRx4r1/ygBfBdMHbZsCbdDerOy7U65FRErpPLQLnaVTAF
KCaOFaSDpXJqMKrpLYvcE0/UFrvTJHdTPmGQQYGpkB/u7SxMiZQgLqhpNRCT6hfjsDIZUreIeiTi
AbZtukpqGsLNRAWI6VNQRy+XmZkCE8unLmMi0jm5kcFS8NFQDyrSLC9WudonkeXnwrWBXit/zrJM
CC2JTM40gQpd9P1mzFnqDnFmnNmB+Rok8iGY1HzSXEhPtriw7FdMb8u2s/we2aWhlYVFHpMtncWK
MOrjXyv9374NFa1GA9VWCKwv7RsB1lZFxTja1HcNvK1em8PGTBLE0MqJl114N9KePqE5igW0iOe1
tOS54jyXCkCXlu/dbJmaZKihOLyDhB51Yy5qUINnmwNFimPyXnp8uI6zd0YBcldkA+yxct4+zD9w
XN9pmDVzU3VCuGMSmDkpkIV6uhU/juWfjqeWyFoSb65sw4y4gqmnWei80TWPwOSHipK4x6Eb7gJH
sPzDxUmeJB7P0SQuKbOaSC8t2znRI0qOcwvs6beYqYue2OnwlZxktKDbG2LFE6KCyGFECo/1zjHA
1lg56ujYNJv/xA0AwTvyI+ZNendFtEDZbhaoxoJGfoYX0+r3eod8s9dc2kdeYOEW5AALn9a4wTBU
hS0DFsdLbWg/uaZZyqR4cFzyuX8rCUM8KdtzmthNjvfgFzDKQ43uEsDh6AGhrj3GBIo9RJzC44JI
AFgefTHp6zOCyne0i1wCYF/GQM56c5rr2EVFwuNJ6G5ny399h3JkIc48x/o1fsCFH6O96SHBeUsa
n6QIg9y0I4TpN6ttDkAjIOxs/tawjJ9vgfTIxJUyemQiJtTDPqlxhGCfh63HZoF0e26igHgAasg0
dq02e13/qvagmb/WgVINVMIIxqijkNTkCjCDSsW6B2XHZHvoy7XtCv1N02eBZRFTWlb0aYoKGv24
L9uHWZwF6FbuisZ6Ox2KsXC3R1WBN6q9qnigEyyiFYNkQOtN/84hiq1WcUUR0ZHF6lBZfll5NjIU
lkcWD84FQLB/2e16JyxgY0xUjk69OW19TVePPvSShahqXUt2Qy0TCBWxvPclDAKEjrDU8cq23q6P
Fb3jDggLYOBd2NCyPamNpmuKjNNTM3m2rnGERaSuv2meMW45y6wTD7zijzosgGTnpPk7M59vrQWC
HQrSOpou0jP0cGNIzhd/nk+l1zEFGgj97OP9IIIIXNlg5c+2vGkfaHkttJ0YDhCyUpU7dkeZ9Swa
IIoMfBgOQOV0CBquAqP5OXGY8bp6WUtBOMHaCWO+vZjJhNjvB6wPvJkJsCsknkHY5bm+eSvK0YOM
dp+Tzn9m/FfpzRy59reXAUbx3osQj6iykozs869fkknGOtclPFAuWbbYWh75jB2vNQL4SNyKsECu
+wAai+Bg3ytuI5g0r3R5DJ7Oq1iS5L3T6JYO1gpxusKcfADbqjQLyGAQKphpLWSjZ+SGERaJ/8qc
4XRv71ZGMDIgFrQtfGyYmwZH7R2vYntrr93c7lwT5ZVfiNLLHSgjHDdocwwX2DkOhtdmTL3Tz0EG
FoySzHNr8YJvdSvxEmLzE/mmae8m2TJQkSJhWxz1MlUtHakQvjeRXksYKdBNMphV8v9JCCmxV/X1
qLoh4SFHrX7njVRNtGA+K0Y0J/ptC3g4Ul/eisO21GmKMmeAO2Ysh7hnYz601oG6Y/7XynBGMd6i
gHnHoat/9Iv6odAgSBTUkxx9l7onURMZmAoC59m0fA4bR8JjQKgynGSpqqdZXWYxcgghW5Wua0Gj
+aQgLYvOMPuuY6eL/Q6FxWHYaZj/fldfawGSRZtKZBVmMteRG23ncpnqRYskX48wGJfwJL3Ku35l
mD9mghFlEj9SzofL+lLgrubjp3asp2Ja+vWf5iECmx0oW8+e/3vy6PPGmz4TGB6rMYD+n4edj8P5
Pvpb0p15PdnUDNvw2WTvSXGTBuA8RqwlYLWBPGRR0N2SDUF+8h94p/SafAZcimV9FQkQ/gV3YW+d
rv8/FPMmhvbHEqSgsZh1XlrGe2IAf7TJ1+PUTa1FboPg8WdRFXgrxrIePlS2F7XYuCHwsD5PN1I0
CidWpTSidRcCCzDp7lbxRg93aHl7E1BQQvFyxbrNbMfCbk3q5Dzn5yWX/dyi5xdd/OKDU0no39Mw
qs07S92Y4JM7mZGbkvawAAU9Edg0AdoB4LImfETBEMIgepI4uPn1rG6oizHC3IVbOSC7ECy2AQsF
KFrIo6cEYQyt2ebe+mA+jgs18dXjvX0znJ+BnRmBhPe6bAl7VOTyYchLd+cvH6avOtd3EGOUfh1Z
m92WBbYcBly8kEfoTUlfAS5pvfRZmLq/sviU1FW+9Jquof8nmII8s2tdj3jr1zmXxanp62l5xkrW
m0od5Ca4Zt0uCbkbSj4tYorgxxEuwmyTnuKyzON2fPOb8GQmEkVBxpo4X4jtnW/lMZbfBaNuVMVn
WYuPPyVHMTHYXUom0fVmQma3vSBI+jxG64RN3bjE9CVC0zHugE4NwY+yfKxPqTvaR7kfSN5yy+xV
MiprGbT44xrxt+wDC73NJ8Z9PtSLppLCdEV9bYGsTPuY7cK9N2SEVxVgj5FbL0vkSMsHvyQFr5GZ
8sbHkfke5RII1rOwBPX2bd4Z7RHsFmH0x6fBezlEHbW2eWRA4Xi6cPXeqH3YziXkuyr06dRwoJSv
AwMdFvdD0/GuMlzboDmlkpyfvoyJATVVh0bN6VQFz2mZ6R70+sqPw+eQVXwkXae+fueK2UQQIDPB
+ixJ5MRwt/EicJYLwpTZA5U6Htdvf8Rxib0R0Lxx9BEgikNYyenNOKegId/Qsq2zjPfJBfrcxVhY
vp993nVfh27Z5rwYmecLA0HchPhfFINwPwpS+qmQWz7aaiVJ4aN85mmljDuwJy/u/0ECA1owN1aT
o4X0c+VxQch31ljklX32P1fdOkiIa7Ir50S9OczKsUWWR/rB618yUaVpHNrGdUmQm7ag7M0mgNR6
AKwlP0uZnSo0GbI7YtOCd6N+6pir2CuKZ2WTLaijHCYKPBEscZuNa5/y/t5KRu7UanGF1PoCQAGd
tKFuq4/DSoHGsXXIIllClTAlaW68ZWee4f68tMn9zTSNEetrVO8ZjpxRjvuxqFPbpiT2rHwe65eC
JRjISpTHB5buVtq9rt/oZAr4VXJlmmsR8q5hcfqr4U3u6qcFHsF9RU8fZFH3wH49ldFB8TfKVdI6
DZGpEJnLSB0mIHYOKtzljNL8AffVwdeGv8cQUtpes/pbI9/a4rq3wixtCoOdBOL97VOgDZMpUPsZ
RM2PadqNujGmMP4+6MpoBMqndRLKPkTEMXMDlFwd1lAKTzMaj8z0w2sH8WK6rqniB+IkWy4lk3IA
EoxelTlacqDYYX82VuEYsA8i5OPytK8Z4lnR9xWzEH372CR/imG6qlB0yEPCUxINJDAuX5zEAsgy
R2rLidi9W9MYOEObKzxtfHIipnTMtckKyiEDeCxlzCpU5M8r4NPVvwnX6boAXSJWpJ4GkAjUonHD
M3cmwFQ2kQVSbjVashHSRnmTw2b4WvtYcm909v8BruWsKhjDQtmJMBfR5L6uKwyFYiz3d+oVSNXT
MlnPTPCQMObvbcj5PvpCj8NrKnFMVV9r6E5jSGxMtktjIOQS5MfO4RbVWZHrxiz7/w/FK6WMeoDV
pJz7MYjc32LKUI036MV98Cb/E0udlD4IJBBwm3kp47J1ij4YBzOsVgWV1RJZf/ES4jZUnoYtsIhB
hpCxSI6kpgskILLxAeDc2lacWd01u1oUip8pBGkNTdPa37mUafGOXzcp6aXZJJtqamBdrZcNFphO
d7Grq2wKcjtXNFeTA84P24ucZZqmK43gvTEz4q/AP+cGoZjBVR9rRqE/FmfEUiTbAGAi9Ui0pVpx
DzJhNrlQ8gxAELPm2O8sMsXGuscOdz8vrDWKcd4avysRElt7hrDNiKezSxtNqThUKJT14aZ2WJ79
Eb3QqAne1+Y8bzimZCIqEW+ptKJGhKadvufBXRp/kQzUWJVmGJeHDPeje7ycH6dqc2f695s7+Nt4
6xHo7QvnD+SUMzCSIX5do3E5Hf/rGNqP0+5w9zM3X3x3LQTMspSGzhVjTYGp/OdmW1m6bL09fZfk
RsJQtPCt7B+GdF/M/FLUOcFU05gltM7eizFfiksRl81/dzCGTXLDM1Ba/J45y+ME6OM8j/mzjp15
ANmsrEOuiGwsK+i0qasFrU3cZaraZ+5Ll/WJM1hvHyw7H/OSmew8+1C0xr+pQGfyj67Uizu+IijU
ROzEXtFnItD0IcZBP2/AtuShkRsnYQxqA9PBy8zQsE5r6/PmqO8t/2KYapyyXmiOqKoKHUjF6O3T
n5lhXWviLOZYYWJ/sO8y1l/bNQzWWGi7emtXp80JlWPOYysKZ8terCFoaupzpYdm1x1lgB842emO
ntSg787dLBoNnHnYsTvnVoVq9MYeyvqsSfpy3KPqACktOOUiOoHoolqJF29gyysYkSg+NTbuj2kl
hnAttL4LQhcyBA0/AUJ1C44OUqFJgGcgafiwcayiDjG5xJsN5EayM9kl30LuEYM8u+I1eY7ws3qL
fl+yOoXYIEsE97NrB6xCbmmEwgLij65CXsatZqj2rsnSYhlDnu9AzS2ec5XLDWRFn1dyZAPmjdy7
nwF2Cal1GILUNfzdbOmveIjDwGlNmvIcPCpbpkn9Og/Ct+yXkMfCrTx6QT1BswaKCieBrsziWlBw
otkW32ZWT/7TKzDdKx/WfsSgca5bQnEUoZaSsK8Zhb+Lj+WMXLN54q+cCSJAlAWkrFZlZIZL7lQx
krX3X9dlaoi44/Ef1wS1hwLgh/UbjuXwR59fpx1NzjbPC1j1WgcRc6LOPK7z4HeT87aZ6mFTCqYL
KkrsopnURlUuGv9srROQ2k3w6M9TiuVDIL1QJi/UUikr78eygvm6vUt0O1Q3lLe+X5jCuhP4obi4
sr01PfYFdWojQI8kFDLwqRw1hbzd6QhY6oIj82NADjK8Wz4PFUYGEPOMfzdbAwQFFpsfgSnqEvXv
KRHLSq/Ce8gC+EfWvW/3dywTHPEpRMy03yMqWbJoiWWbBkZ7HR7lpCC9y2V30yjcSQvFmnLFXJGZ
AZJzJnPlm8KKxZhwOxizgNVOjq7Zdh8BCsRP625hP0C868H7hykPdkIZLk4dhGvWI+Qz6A+UUZWj
snpFX6zBo7R3lZJAi0T1lMjp82Qo/HjxGXlZaP11FyQwOAqZUPnBnxxDe9k0fslke8CiNxAWvy4f
SpLMI4C79eILexHpZ35krWvHc6iUiOBKLnBfQFFg+oE91HNRIcA9RT93tX8sUZf0xBtQxDzGRb0C
PzVo4Ime0Kg/SY04MN9zQtHKjaAcNg+AKWwd31ZuDPvN42Val5HtHBkqvxqpXos46qQzpo5pPGgl
QWtg5zdbdnS4Rl7tY4oqfKfv1FUQikkrKOijaiP9ug7+pgcT9VSSxGCMk/U7ebFXFSzw2iZljqFI
k5N4KRqAKnzSYEV8KvI7zLJ3SDmeQaJww63cbwYwkYwEhiXw7mImUFA2JLPJjCZLTqeU7qyJijbL
jmPKVsKQx9eXAR2ez41wf7vyZancsZwlsgJP0+DCgUPxHLj21s4AaMiEkRjySNDPXt4AUaQ0TP2p
dI6yPZ24oQn6ZHpjCc+0AAgEihMQkiUjHpWa3qggaPyAzXRUiJhru3q9zWkhPFa8MNKWjHDGPY42
OrUx6RjAPG1N0C65E7ES6ZxJthEDPzaKg+o0fRAAOlqTOBpfO9nibBrtnYzIHCwCoFpp1fjCbyC/
1kJ3R/tg/cAN44Tj6UEmJeVh1FM2GTk2fdQveYCAEXR4XgEJlPQcmbtT1q5FHrGXkBR5hntI3S+N
jHKpVtlPezPxHgC6qvdsAw3vemCpfyzClmEvBWqnU6CQbRXpVpe6GcYk/D9enRTLSIrhovKCePMy
oKZytNbbOJsTJi13nEjvAt93JD1varxbQVODCJeF7HVFIxJt3kZf0+A4oJRFnbDvISAuuUCIvRck
MNljCsKhmCRzTdRQmLCuqxtEomoSuMqFXaOK/HIe+Rhb09t4Y7DhuBiA5AsYlT0oQOzmIZbCQkg4
/aYP3/2tUUE/F1NjwFc8gmO70n+UKsklAznuVMFlFeJWQ0D75OfVCFH4x1jnn7Z6zp3RbRZShhMB
1/qffmoCHoe86u0pbHSmFwWs0ySHACkX4ST4WyyP2PAzzppwjTFsSP77KpnnGHvBEwQc/1W2gAtB
jXWNZMgvSvQQl9CUi9cYKCS0JkCRs19hRZjQmARFAczh1NEanT+qkpSoKAGuSmr/n3hAXwZ0wlDv
JNQTxyulyR+6W8X91EafJMDhaGQYPafX3u46wTV4INWvp6eGuruatb8IHq2UzGZeDDc7hY06rPjE
HEV8YGzuPzc6GvE85yNtJkR9/BUTrOLW5PuEk5XLr/OlFv0KnIE2GTN/HO39T6E8E6Mct7LuuoU2
R2SxlTRsDDEj8JUScfemyCqz7u59f7U1Vn5oNUAlVmQhbRKwVpQnGwxMMx0L06dk9DmIN5MxdJUs
wWlhEMayQKsjkiDMnXj0v5nmnLgvj/v1WoZtuJGJtIT4/fCohk6g+LcmIbFRcE/7mJhkqzQxycbA
CGtRAldEtqXCcpxoZJQPK5o14bQIdEdcqJ7Eo+oq611YWZrgSAWKQaKFFuSoB3gP825Nvjs/jurO
f+E+5OqvSsCg9vMDVJFGb5cG5F5dKZQmWblkOyyTDG9YGSSiGpJkf4S/p9UDxTpqByghMcT5Zyji
dJ6qRKTbNx9097q5tYYSPDDA+ooxEEFC1NZ5f4iMyIdFWmhDdra30z3jX0JtLdDQMZ/24/UJu1dU
AXzyEm3M3NbtjhRdrpaJ3+b1HiAgIdHeUSa2wtCO5ZArPJoXleKEgLyMjWAbJ1eMjv4zbP3xVJbh
f/4eX1nf3eviYkKDXVuexCedHz0teJM14fze67dmn5ygZ7u/Bdq/ukzBBEXDAoq72tdqd0PAjHcE
iDp3+Frlz8u7Jm6ax/SuY4xbtk5853slVbQCbOdG0B5HUaCIehz7YVoch96Lm40RlGfiF0gtMtGR
6J56yCLwqhYEQdFAQDkaY4tNqDLzE4NGjbYuWi6F7BFQfjQcSX5by34YLHFOHNwFQfNdJh9d/of7
uNf+iPaTv+79a/6R04u/Assd3n9ZkEuiHBiCjHSeHGjOD77vUunVGiza/Z+TSQ5uBzbhuny6fCrz
Q/vpl/BWz0oDS6jATo61kUA/sVyQeE5VO9V2xAs1pObk3S4QqY0QDqhduSf7zRe52k13C8sloec5
pQE9z1XcupRUUIf5FAIISV9c6S9Sa9bGCkadfjWJWRJJEtlo0cTlNbXIEFiyzfeoWlrSzC+FuDiU
CCO1OHzGWua1mzD87LcyEeGmql08QBT76kjBM8A20O1VoBdY2pgNQ1HD9zAa1vRi4wDF2kEGMThE
cuzZqyiwRPiggIuwhB3Ar5GDzjLO4+dt51jMwqV8ekazefS1YFNkCX+i40V2YQfMbQBgiaytOBWE
BgbLO+6BzbgtD47svMN73U84Ww8Fg29kDJZBGFiCtWu45anmS9x1PlSOIClP79U1u8PPITL1LnxP
n+etuh/2t3qq2cOx4YbBw24jkBaDJkRUO/Yv+1pI/Igy9MGmUZrhSoVhvbGH+VBbxNYH/sAfvmRR
Kp9i0nWpaXE+0ZlITd0/0leWGeQkvd1kzE1xmpSSBO6zgxwUZiVKFFDL7lbPO8S5DJDhTgtSYM1i
IknsnvWci7k/++8L1XT/Ju59aDMLeVWO35z9Dz0LDK7CMDn+bMkMMJcd/Uv8m7pe4KrSkdfU3YgH
STbEXhGu2nOq7XsqSmoQXlrr4jQxyyPugf+kGbTz0IQPEqJ3ovBp3VYKvfqlQcnbtPxzczTUGrot
fUfDubXdVQ9I5zNiU62HNlm9ke7vQ2bUiMOytUnjEFRPxiHbo73+tE2ORRpbdfVw0DMpmhgTQ7eV
7yKvlpoV5C+kh4lh5LgusuFKE00+o2zD1b1XgbN1uEpG5SQws71iy4YcRrz6ZWuFtE2zgpi2m+7q
y2ztfkIfeP6OHd5T0ooeSq/GA1peACoyJhXfFcSQfCMX8AkjUW0ygqXlhtHf9/19u95DSdDeIfyy
ze9DBq2zDFDHRcb88vNyeTJUiOy6iV4Uu/Z9go1zmkGF2L/iomujjwKLxoAbESmUD7NTZ1Q173WN
1r5Ah6iakqLNCRz4/8pm0zQSrUaeQh1DzPJl/RiiCjjADhTZziGU1rQYk7txhEuT8ReloLlRQnlv
hxaS7Ywfrqo+jOvfDpw0HIoys+CzOyyC8z67LMpKgkiWh73T3d3kpVu0bwFBbFbqZHLjBELPGx5V
dAkPt6H6do1HkuqqEyn21YajwBNHj20eXUclKznExriFaMMvNG3bTVwkKbhf44AVyeDuD6dDWhba
HqJP3NHMjKqVF1AnxNRdoNqabsq6tGS+uVONimWJgXwiKdBDAKfob0MqjUvTBeGuU8kY+vh1SmaY
C3ZvB6kGNb9RD5BwhnFwHTXFGiRhtOo2OIHf4gnxs+hPN4pVZe2+YQWuXN9AuLdaspILPi52e1fh
PJHW2qwnHTGFuxl16F1gaaTxFgur+6/cjqSpixWtbUlS7w4rMM2m7lPa7uWA77Ch/U+zOLjbgXEs
aMpj7ff1QfngLkgGl1X97f9eFKjpTF8ap9yfO1nff2qDW1trYmLYxaDcAR3O9unGJj8IaAv7LqxM
H0lY/Wy/F6EyKQHk4uzEuFu+HJz6FOyLp6WXR2SeBnbHpTjyQxhSnlX/Qw/xx/4tbYQGtdP1V5fj
1jlSdpp56pA/Q8LkCrdCqLVsdtslSvbJda/QVriWZDCbXF7bVyZPyJ1edmQgGD46NB8c6wtOuxnX
m8CFpSdYxW//itHrEt5i5gOL+W2bLjswiPLkdA+XPGM+Obq3DcY7MATIs8mFuacP+QnD+UtKoia5
PSGzUlcPgx9iTtO8pkfU0v50MWbGWwisz8puVuq2DdR9pWiPDGVfDp/wyVFDmFBfIjSr9Iv5pD/m
nIibTYBalI2FjcXwa7JqAmI4Rs8METIOKH3veiywktW340VyuVMjmUo2PlZ76x1GzkG0dlytO1CM
9IxbHVQne4V6l9QQpcuE4MJ+mrJoI3xrRN5g1Q+fpNK2ME6WOUi2QC4iOrK8glv5eGp2HubKYNJM
RZkEOfihPctEz5MetJIKUqwxHGr1+vUn/PCi50Nu58uzvQK1qdVoITAQPljsLMa3hZ9bLSws+zqe
i/DDCeGFiZbb/ZJW/vNpk2TfbOLrYxKOdK+N2o7EZNlo0z0rovVGDuFUVwEyNxYkdSGLZBbZFHLc
auAHdDA27RhODlXNPv77LQw6QPIN5AU7AuzvbTbN336OjFDriQdonB2Y+kiKc8eIP47kgeb29MCM
QSbltkZ85f/N2B4L9MPy2hBjTsgNzXt/xwWaxoiHOmFo4tk4h8g/XtpNybEAeexdYy9BY//6Nz48
+07srlSKho2hwA9ESL/uLXZB+/m7r6rfQj86EbeVEIQFiU//MkH5VjHK/dFUHp66/LplYRSRBINe
NZhHk8586RgNB/efAKeepwS1qhpalOA6AHFtXKhmOmwMSgvHNz8U/kyxDY4+PuQVPH4NINRHcYA7
lw2lRrdkIQL+FHLX4sSXdX+BDnA262N5sBdlaEVZRF5g9r9cyFtGz737axlacfY2Lya/ERQh5A1n
uKqFPqCGvFKARjgk2DmNelfJ9MWqVFLYesPpWskiQ9FmuKNcuEztsAOQX84DpJYAPum4sNicObVb
Up38rBk0kZLu39+rYpHRWP/FJhyq1NGC8l8oGNGfrCRTrJypW6pRWYrYkUtNftVdje/9ihbWVkZS
b1SuXntv7nwbHOSeaDlv8NOhOlQkIzgQqyfZcKMenTuPJOt19LrvoZKJJ7SKXccqZ7zvHqiCu4SZ
+uc0VEOQsucvE1NyKkGNn9jPoTsDvrez6JGJ48C56fgyUvDCYVfCEeYJaAtq09hpE/Nx5rcBrgJE
MhTzzunXMbjdK3ogWyAmf8kbLOL5P1egAV8X/SYdtrLGPqnUVB8tFcMzhK0qCUAqZd/l64aNdYmf
0ue28c+0dAQMMVJ3/pr9690i5oFO6TV0moFpJFgswPpfUX0H1cDDQ5hg8GEctqQ5eE/6sBA6pjDO
ogT519eIQg61GL9pOBiJlLmD11xe8kVNIcv8VKCx3AIr2klWsecI8BhL3ZYdvPRpXpPzIFuqoAT3
brl7CFS0YbswmWnOE7egAS6BhnfdzegcU1hlB/9RQXsfCfiTBgDr5SjS7cm+I/Na9+67QytERvFj
uRh+5H9Q2Ci8s/MGqdiOaZN5R/Xpi2DKxjNcnmig09q0q9+RiDuvQegxoXNdcMPzZfZGH21kLFP8
Tx/tTywqPFagGrwcAfEotO7okUwyaGeZ2mnzY4Ff87kN8fu2VGkoitarU4AqOoi1YP4ZXl22G+pk
RiuV07fZPUb+OB2FHSoTlmQ6oAxadfTg6Q9i6f1UPf9BDmpgNyU/DUfzJWKQtHTK+UyCGsN4MqPI
ruwFDgdRZUFUyDfUNq5d8Ipa9Pi6/AUrOkDurFS9VN5TO8dTiMbsXePigBVYXQLhKO0cx+sDvcfG
2feHusrUyQn+RG5Fx+wAg+QRYAE3AtcoCixdHYn4Rh2lVNYSMEHAW/nCwfBnYUO3KNoTcBN3jz4H
ao0fv91Cf73PDvc16M175pbvt96voJVanAnwwTQt3NjAkS0hhKaizqY5MXV3QLbZ3xxzuqXI1mf2
2v31gRk/IGXqgYuAB+7NOfr+r9L2sHZZ0sfj2pEYOdZyZXHFWGGgJWYc1gQRoY4GAamg5yrRw2gN
N6ORugddQB3mrZvAY9b9jQfLvWO+EkDMYkPtDtEvOIgzTgew23u4YCDTEcwQ5ETr0yEllOs9g98w
h6ZsM9XGY9KulUZQBVeRf8EtXAJO3Jq8b3saXn0jykDiF7BeAcwyrhYla7PFce8MfKHGfZgOlQVK
M0pAwxOhodjoFx2E89AGbog4Hh+3zXiyccnYcptCgXT9PCSgNaCTcgSBUWZYfP7TftxL86edaWy5
RhlT5CfIsJ3APARzLjgDd2zZaVWxoo2z++CRGbx2UHlJl9KKhYd8rQvBierE3Hy5TVdn0cLiZqO6
Jaw6dWoJV8/MXdoe442bU9Ivzc9RYyUayzcdq2LQ9wQjv2Y+BVV+/o3g0QPljm0sPDvD6gltJHeW
FhM6k2qa686eUEfNxR3L0o4JoPcM/1GPuLPuaqVUfSEmufVR1wzzEDHHSafT/QfP7by+xkaRuQY4
zmj/yHQ+gf2mJvB+i5AJN+PeUF5XDv3UH2mm2+lkWDGVhtcmLi/J6s1hXTvSUwZ8o7nZqT8fgoEy
Jy8lUxjvXuKpARu7TtrbhM1OBtHBLagAkJcXiZV646CumlnfiiUVzJMZnkrhZgMRYXyqa+C9Pa7G
V8fMfHcL8s6KAtN5btEHTMy198io8BsSUoKVvDD95RPzirwrVA/klXJP9L4inuECVgLn64lH2VWo
ylaJGvuvUcPMenUoRXTPQd1RSJ71IH1aal8xJsH7p0LgMcK9ULTV7lV54ARsLeSDz0h6hYwVoYFH
6vaBjo19vi3nnSvEzvQwBhXhvzGQmlM5ROexN/HcPloNpEw4G6O/9zDnzuEiHpsXUDoC/Cqf7U7w
D9CtwlRI45kShXkQtY4cWy79S8wlIvUmqJqx9f0mGlJgFi6ou3Xkq7ZMzElkASR76t/UaZfSUDrf
iQEm41HwYV3ZSVXzJFbLafJXEAeyKzgBvoppuIpN4EblPL87mCLxv/D9HIBRh3Ygn+FMnJuaKXUi
P2zBOMjQTL6QXsPTvvs1vGcpdYr5ABJFIra6DvM7u9wRoJZZOviRdAe5Pfrrm2WAvYvSVCwCJGnd
DBA52OB3XBYFjoprsQlFes0Jm5Fd4EayxMHNlBaAB1IpTME2jFqsNdJfuHeMWvw/BGfm/226Pigo
ltD3VJ3TT4W2PwbgK0bj51PFFdj8KfoRn3v2AfnHMag0dxqP68HruXiYlGiOUim9Pdt29Fsl/cld
/yjwKfCILDD9Le0lPu9XFer/Rv5rNK5LpOGpHii5krgQP1dp3j95AjzyhZaRTmaCCJR5dwsj6UTr
Dq3LlWFBsEfrEQeiRL0z8e9xl2omk7ucwbyvJABCVtPbj3thQpD/mE5VGQbyyO02Hy3iX9O9VzHi
eg7BYBiPS6GHiVTnrE+2CpdWrrYM/h7LlJwZVxetEWOO/Az8iw1TIcOYuPr2LIGk7FPU9WtWmKmy
cgLwNBQfzyg8pp+OeVrWiC01LUWieffVepSFIRuuRddyC8MG+W9PlXa3SWdaUpraJUDnK67wIeOm
VMmeo5Qz/fmBKEeEJTKqDGMrNUR3kYQpH0eoepxYjrU8j9S8bsyZRW5mvw1aG2foBuJafOTCGoAE
ECsw4eW9hCx7sgRDLD9I1fx2MmwT0bUL5h14py/uK9PUDVgnpVOCBvqUXdkSmCQ+YvBcP+QhKwIU
yT/cR1RQ4hZ8XolRO1hPli4M1oOYmXSW34Jcbm8vdI9Emp+9rQbDXoyNJgxqntqQsea0QrpIBlGJ
Ij6aMdApCq4npYtQx7yOVKOlqoTZP4Pot4HjNTL33TrxrcVNqbodzlHfLPaXR+s931vXDv58bkPB
kh1wSwKE9+blJecMXTCxdKjfyX6RVJoUkuKyDtLviZmqdRBz9ORaiaGpBxF9VpCB/5cpmjs7hgp/
7cBzmRQb1uI7feR20vaxzU1A7825PIzE9BFgBdKs2UvRRLqOycmfugtniLNbgSel7NAzU4eDgkgS
ybNeefhgXZdY3kcvBfjpHOhJDZdOUNNR2vRdPuGbWRg3IMKHVVvqIjk4Rd5wJ2X7KbJV4Nj/mjRG
yMKUQ5BVmc4lUgUQ2YaD+7ycjH+qgYvpg1DqjTjmUyUoaaxTH/z56c4xPsfD6GkkNa/B7mKeZdwP
WhMxzJZGqZ4tHt7ZVS6LuPazYPLw5FeEZk8RYvAlfttf2BDPwebipH8tjVZYuNGFO2I3XO87J2sP
+Oo7/dDAiJYV/s63d+aiF6Oc9cY5T69DIonCxLAo80ysRLUuB4p8huGlXVQvIoBPHlg5GHGD+jLw
yUeXQWflAu7AhzpY/9N6kA2aamF0Lhu2v9jK9Qk0jWFU0fEJBvTWMajT+nUCQaydXYUKOePKLrr3
Ip+PzPo27SAGnapjKsaxO0Mhqr1g1JabysWNJsEQjhqJh/fBEmEpxmi//tpdaVzfSpH6Avy9qAnQ
tlchPIzoeEJG5oMdcKe9zzV0ogbFTV1MimJqgvRQNrM5sNyt49XxiA/TB6qA5y0krmz/MZlCcpZ0
Qx2mDOxphIL3rxTirWL08t3+TjeS00YRvooaUd2yURardg72BrbEp7TIdu2tFP9vqoXBSbIUvIVZ
zo2GB7s09HYXsvNV/5S9RXz5DU8tkT3/d8NRKN3dqI7ZyAHQvFRCVtjKjJI1MJNY8mj2MHXYQdr3
WxARkprM3u8zCHrx9aek5Xx76pGDpskuZsoKsi1fmbOvkrLt8+yZWEx4bWdOLVhykMIt8HIV251Q
J/7bQqfU99x5IGsZW4k9akPa2WcBXikLkmbzhxiVjsudXfA0y6rbD3ASXn7VnR/XvXQKhXqtcqd9
0uQnMkuI52CvBkeqjdAlQnyEc0tylpHZhkToqm2lI2VFist/6m4Xt2c+3o3qnC1e76zIsU5v/sdG
Fq7F3lWa4/Zmjvz2ByqznUYBLJ+MLWfkfPcJuykUKrz/G3BidUOYae5Lejz5uKEcTNhYDcUh477j
m5V+2j6C6JOz7EmR759St0D84EAarkQBykVxS15wvZigNrDZWYYTqQ8hwsX3skgZnzXy35AfSD24
ByFkXI3Kt/6yakog8mtaDvgnUL+w/X+y047bJDrtQEXFaEZAF7Yf68ISs3k6drC+Mjp5whHF+5LL
c0y4zG9DQlfBhFjMWbKJCRX+6EhCnoYUO0BilHmyaiYEQUTf82G2uFa3TIyj6S42+zLgxn0uiLjS
zo0z0Lb+/PJ4jT9F0jtqegX8VEDbQvoIB4DoLkQl/1fZHB8ECu3Yg6pdFJoW9Zfz5q6cokE8D0eU
ZykuIznEvN34d/lH4E9nql3R2+S2/EfQiTKumRC8yc+XdnxKUFzw/QtjW2NGadLDHFFjTW1HDrMg
zzMFFMWXaG0u7izBrga/vRWmhtK/Ke3VqsDcLwG1/ATS+7stZnnVKN6laHdRXdJKoOanEkxExzze
liW3b0QPI+qZzEvuDT4ndVsQ9qcEWAYdeJHzBhcGoqBCvUF175Wl3e/BbuscYAGiqecsDd2eQlt9
vbS+D4PhCZoSayEpJBDJ4fOghqWfFb6HFITTbkqDFYVfVfEDd4zbW3dziUOOwFJ60KyD5Trdh9ox
LXVkY+pGBPuvPNbHiNoVBI8fb8puKdbPck4TokngnHaUevX1hsn07UTCBelerb+Qp/bWs4SAZ2mx
LmDVbBUeC/jHRGI/29FBQ/YpMCCTDtlpT4uOdEObhM3D7qQK7TEW9B2kpLk99xYP3UtvYjUlfOnK
qx8x9Ns3DZoC5ZE264ShMRnzdEpPTEC95LO9I7pQ51AyWhaC2vfWDykD1KAaWES1Z0jBvoZiAiK3
npbvu+BTZJQ4vzsPWWGZ8v+kLwiZZr4uDaz6HHOuIMFk8FzBG6Bhl8g+/CBiseeyybADEuHs9PMP
p/sLMFl2kJ4fSOMKUhQllUVI4CoyJfw3Wt7tp8NMJtRI371BN5/OTli2q37QwJ3oqmV9fkUt6KrY
jvDpGV4VCFfqBCDI0pcSBXmAR08nMJ6oev8c98dkAURpEJYP1jjW8EX3o/ZyI7tpv2TUmYdt7U7L
EEHfePrWw3tQ9aZjV6yA5crNX5TkXcDWBNzDM5TlB3wJNU0dT8vVqlyhGNgahTUKhgCQR2hj5sNC
UmOPuUxjjtBjHjtufCliOIsyEjk17H6UZYjb4g8JfA93Xkdx5z5otl30OVrdjGgOHM68iw8tWEFe
4NXUGyhavjQUviP/6m31v3dCHgXlY0Mxc68j1hyHR0cpa9TzGk4fi14+tHe730NEWJUUFqOLki+8
EBIzEO61TsZ3MF9MZ1D3h8lgopR7uWFx+Qu71OcAShmUwu/+92yTwhI3wL8Qt2R0Y5LcMbf8UEfC
PNCA5oQWiKyJVqwPEbJ0udZBxOnBLTELb0gUMRNODpKmVw4W3MNk9uCLOYR9dbm4IfSXd9Q1foXV
Q40bnx1GibzpjsJwThlz1DEhQRv7J5fm+Jfg+LRDtTylgxS9mt586lj8va/j1B21rvWQRyygP4zh
GESf2XWk7urF5DxJMGoB3BN17w6O0bGvMwuEuyKinzPBxkOa6rGfABzfNKTA6LNSQRPH1p5pT2Zs
rhrCw/M4U9yLtngOSJICtwRvEK89Mzh4sgi6gVra7tBQuKr7PgQvPULOvBBRUQ76Uv6Ar3CsDUcI
PVAeSJ5YGasJ1S97EUhlWKSEVTzPOl7yfb3gUnwboB8ddVjQvOrQcH2TTQ1D7atLKlByY2e8iQiG
6hQE73+QVXK9cgP1XSYVAAEzT47Fj7SUnIlZp9Re67UQa1YZW0biNSOtZ8AHmy271iisaB/zw9XV
UFywuMoXwN7u6jvlDlh5Y2P37isrC0nq0VEdrrSkkUbf9fZxrBB0UEtjxZcocoay6UqCWb8sQTuo
iPgtBD/boRS9j9RNoG+HE2bwA26lvxOAO73LGX4MzYn1oMfu8lfcxYuwTC1GaOMB1kNPU2S0CHSE
RusZOxXxopyvgbbdXUsTDfSXgm1e+XTKs5SbQo3NtctOgbFQFkbO557LYxrxtLXH4bJfp2xzHIvV
PFkf+HpVYsx8K05EcADywVce2AVevdHCI6rZ6Ce4qf0ZeSS4mjeL1O2ZP45ND7DR14WDZlTEK5H6
52M2VzMpjlG/mg+ls9wAhoxKEtXkNB+c6+MGBo0pTFN2vYjFyoX8DT7ZkDl4h0s7Ye9+IPAPef3J
ssRb0U2K+THSfC/TgTlihjH0TZicsQ+3fRDyEiBlAwgiHjd+KyAVWQCbkhAbHXqG6LXw1YgM3b0s
T+77yISom4xPE/+15nksgAWd1xGyv2qLeWYI2fBHJyU19LOSU5Kx7e8jPuuhh4jVzSV2uhDb8JhG
FyWuEM6m/mFcBqKjkLzU2nBQvCgHlKkuStVsksdLo4hvu09wpAE38F+3airgMMLMqSp+QT40eRtK
I0W9EN8lThqdUYaZxPc4C7qjHSiVfh4IC/yRF+PUpNIOf3pAFbC5vmJLBLEH5uB3bLiihc0C5g9Q
7IsHl6uapOqwAzpxbRUDxGRlhZ/IeRdJKRusszYOvZPI8eVxUTVHKXZBTz/PaT466ZFEdKx4UK4d
FECLIWb9gMOFFFcsm6hnzG92sdD5Vv5R5pxkP7YjndAT1Wp3Phh0cwA6LMpgplJRhzII5+UsJET9
vxw7bHd83ifURSqseLTemzkI28hA9U1MOJt9khh8CFPJJbsUQq64J1nsft9sBCh0CTvMvkBGiqxu
YmKFKENLgbBXQLfe7Qk+JYBYNib7LO/fxSHPWKR6BFqw2BOYpaN3SIHfA5SNZCrZ95tZJ6T6JCME
Q3xqzfH6vhx0zwwqsLbgzUkg3IuWct+Y2z/OPvUgxuf3tdlado1b7DxNz2k8g/vYBz5b/LsPCkOQ
fcZL8cXyJ97Fm3JDfYrJUSpKjWyUIAHyLlQXyK8YACwvzCzaMQB5Lg5y8p0gqjy6UgKkRnQYQOR1
gkti4v12Z5a2/zfaJr60RPnZuWS3O/1QUOCaZ0qFrPNE1WC4R7tkfzSQUCws4l1JhXt/ZXTIo+r/
Xxk3abOTIc4/pyhIfzxpmOnMMW6xf+X2wBfm+E/n0tkTBxkYq9CzlTNtyEjc4nhkeGvGyoTpcK9y
Csg4Ln0V/HAeJSCstV01jdNaUvJrcozDVNBK90UH9sV7WfnECLftcu21TgdWpbYvpeJbvYSv0ep9
zBVUNgUCV8zKgJE61mAHTZn0AdbcPO/K9bOdtvd5QRkOE1s8Hy9UoVQCOZgzsJw1h2tfz2u/Qm32
WmJKVPeChijsEmcVZblkwiXI5bPDoLll1nzAXfUrk0WAcW8ASBFAD5xLLA2dnpMXzIKveXGvCO5K
FD6GhPAWcQRtwRhhFJAK3KIrbEOcmH7z92vIOOExiL2Gf5M6bhyQ/xv9hKt73DcbpJUNenii/ngV
0oss29oKb2H5JJtivUbgmb0wNxDV7owZ+mqrFP3k5tud+sOun6FCQ/FXe0V3xCOWsYz6R7ueP0TG
vVznkuxFQV4di9lUb8cFMa8+7SwmwYc8F7jNYk6IUI0RFiE/zcQcubyXso7qfl4HpcIKgB6vnfcG
gw4useyBPti6beRjFk2vgKwgsYq4wXrfP8K+mQJK13VAfHkh25KRh9+X28omvucKPwf9TXDSYPNr
absLhXzmAMQjw/eIpc7YDnCei/ooFn5XRP4G1BU3RY1wJIIctbikPTfGimSGPynl1d6Ecb3mJ7/b
ZjX1zlwU/LzcOBkBDwHpU4oy5t/t54cNha7UUIDZihRvnOZt2W7O5lfP0JaqefNddE0QLXQrvnXU
xBOubPxejUe6Skg4Kfze1hyU+ttDf7VeNmfKlnm3MdBzcP+tVPh6HmgOSmpEXQJeWpsXWpgKNv3g
LwVySxmoKOhMi5hM370AJAHhIdHoZVqdwhyXg8KHkksA81EQiuDdgeO8ET0OkpLZmh4kljq4T8iy
EZ7jD8qLLvzuNnwrD9l+2H79fgjDmEpPrWrwv7N9BrAYgL3aCKX0vz2N6uzP+xLXsoxu01xoEM4E
6bin8Eo0OyGiArEJ9S6nrfNoD/hEPaTThnMc3gCqAEJ28qNG2yeSdU//jHWkeIke9sKpz6RnWXEW
rkrytC2A2XvwKAte1m0JV8nWcgKnauznQAY/5nUyBh8JdVRmby2FGKbZaJYgyCiL7cJPHBledwgD
UIYMYRBJurywMIuOPO7tnz9TmxxUNHQ4s4DrHmpVPvHoOTr49Mh0/Wiy7cnyFuPj1hMdCnOTgEtD
5yp4oKyKBLORUIL9Nfs9La7UG/u7bM0qWbhT6W52qVHRmcuZpdEhsscVbUhrDtVpvyVVIY1jP2Zc
+gUona/bx4VsJAc2s0eO+udj5ipVfbmnvzj+8ie3yLprEWZp2LgGQQZzF8e/SnffgigQvRSY+S/O
+Zyvo+I63Qri6tBrGoSwenGpLh/JXJBh9RUKD6W0O+fPEF3wMjLjAIWO1pMAdasyUbHAAVg5uakJ
lThkPXQ1DHzeJTRDFcaxuMZkgm0dvPf7ThAdHGfZPeEvAvIjDugNbJttCtEaFgNSmev/DXaGcEhV
8xIibf94Vns1jSaSKFJ2Qk7P2vRoAJdbNNcaneSOwuXADbfpQqxKw53vK8pFsr8NyezS+DttRwF+
UVT1KnzQHGlwrJ331/4AtOyJjyhH9fmyMLqML/AM4ILMncmrkaPWHkWGsdZWBQS1SeHubh5M7/1d
Gzifva4mVn6m9oG7TMSa8QXBnuwav1LdeUsLctT0LFslmw/p3bjXSi6bfdttEwMPTMQG6G4YvNri
zjxd9oWnuccbbs3oSt5S6knhaBHCYPI3/080I+RxV10uNJPT1SxMWEqfL3pKxIG8mbpgU0+GXcdV
azIrrrcmeZ7Nc6YPiAYQQ7brQ1dpr+Oe4NZ/P7Ja7N1+G/K5doU6U5Tky99QcmchyBOg4lDurJWX
XJbkGnpJx6T/0t4UEi4fdmA2bXo/xlmZShK34+vwJN12K6s2nphMSgRs5LEAaz8d2FulJy2Nc+dv
KKho8AS8x+mmNn74Zo1L6PcNp/msJc9mWxlfWMAYha/nhibBwqD7filWFJsYbEUTloMExrF7Yyq5
9rjihWEp6JjfDa7A+RvUEOjlxjcgNywPGHDk+lsIoKT5LHH/AXzNUNec85979LreCrrDaudOKzaQ
ArRbJ1K+9a0X+5uQDHJ1CyeAPN5UqOlcmBWcCxWvr0PWMG2bTYobEkssy53KxSefyTxmPcDWt0tJ
cCLRiD17vk4Ew9eHftBQRv31tG5XK4y7Vbq7MfDQY/8+snvRhMa4ZmhOEgY0G6/Zv1hdOSpLokeV
ZBvMx/J9JSKCtAQkyip09yPoBOoE1fAjx/62/Gh1DGoacYTIJqB+fWMufSoGr5K4T85dknWdbzxo
R1+OVgf19FX49B7XOTItvLvwl8HKs/B7+Tzox5BBkitpkbjldUE6UfYfPMoDYbfIUi5nN0ZwARvI
RO3EqQ5/PmuWo+EB5AyLbJ5Yu6oEos9LykL89BS9dxWVK2CF9egnPy097BmUaLkX7Z70bcPceF/1
6bS8sPafdH2Tj3ZA1XYrmiVOBlPgfzCcW/Q8dUTsi3PvcbGkoLuX/7di8qA5OIWPpUGB53ApHvmg
FaXf3McoXNyK6r+TrZLYe2IO3quTup0LtWld2itq6NGK9pnuO9htKC8Q821zZ17E3I+tdzBbQeas
GacW3o5J+Gaept2sVXKRWEi9eFMyMjzrx53CP32Bt+eidE72A3zG2YMfP61yjbW3Nkjg7VZXeaEx
H1ASMGQtoYIJy5pjrQz19OVTZqFtFTJy1KO3hNb63sxiM8PpUKiPOLKzPh2+a+IzF8l9F+MjzUia
gAepKAacXna3qqh9Yq8bSknHKtCXbvrWf3+A0m3o3GhMOjyvMjca7DvNujBT96s9961RIa4SbXzB
4kWekbjAI0FFJeVM4GJx3tHt0zklrdZzB2JJIUJh9JBhpu5ajaMDUgl76DDZzJRZdkTNOPIuKIm8
PoQIWNQ51e0eHyWEF2c3TRPgrZzvaeQyxO+gZNGlGqJHVCZjL7kcBvvAIvlCBjmwcarqE7QGELCN
pzLhHV5YT86u7JKu8gThnNLWgzoc66KBfCm5psDClgTfXT+/zicb33xUSM2hgdAkJxSk+MfjWjts
LrWkb6+EsrfywffeWwlEMtUP7ESFQOTrnI/JxhA3rsvu6ZYsaZeXXVjohD5ISKIiC9NHfYiJoIEn
oQHFY7VQLYAlMDGWZjsIPqlPZN/KKSsZ9R0upbAllKYJXysclyRBwnz887ew5h9ZOAxZD93grmdx
rLe0B8fmnk3vQRVWvGooseBpZHCDao28z/c7t13o9Dq7ll4QjZuXEdAA7Bpa/ro26mOxAEhVX42R
Tfv64J3UR12Aid03AcXsU8SN6utFNXN9lN7awpCyWv7Z3idn6csZwzj70FUi4zKb93ouo6Wd4umP
5+O4xfdre4AY3xnqAuBcZsb8bjLN5cHspZv0uRu+ne1cvJq+j4Sh9m2gYS0XHfvmf7DjSWBKU7Rj
7sLlOl5+d8WzunVyjly9fI4ZIhyAzOnTUwOPNZvz4lQDyvssg9fxy7XUkaS6+PYbxSh1wRG/uJJI
ZFhYLrfvRX1TtXelkaJotcWl9r0k6WCKAx6D0pEyYG8tfteyzUBTCav6ubQTdKJRbRQQtW7nYEPs
Y6kn+pNO/S1L9gHG8rMUdAbQDMLhddxSymXbAlNJamyQaCnu4xWGMfIj/+tq+tvqScJyjg2mnoos
Ekj4/j06+4OHIFOAFcBMsppXmS0jGRdzQzExc2SXp4K52O7NRbXeIWQs1q+Yce8zBzzi2ntm/hvC
LXuVGO6/VxCdwLseohJpcYfAbovnCBRUl3JWpNgHYKrCRGGJESecKIqXAj8ea1tv0d/gWX7bimYY
QmcWZgZYGXlveuPSOeEwhdQJRJMrjgTyi+wsQJsF8TTzzADEBVkuuRPeJ/ZSRTRNMyRmVhnh1+4f
PI/v2wzrNMZHElZ/2QgdtvyZm5xWFmMorpqn/NHdu63+M1J4xQdC3I3FwR+SdZ3IL57P0MwtYUQY
WV60R9i+jO/QNqM6L8YLzsW0PFG2JP3MKg3f40auHJKL9bi92pND/s36KG/EJyZDIMQhO+CZ0DnY
TxULtaDIlUukJ6u0TjiBOHa3lqGNefc7Q8e2KrxGbeDvufMYnSksEMN+jsMNB6JuiJdbLeyPN8EY
hptgJN7zzqMyab/081xkio5Vc6OZE7jmk+WwH7RrmPRT7ns1a4Bo5MPBQWQ8tlrc8oBmYsRt4q76
0KqVfkZNcO1LuSP9Jt4NEkUEf5Q0DtukXlY0hM2J/iJb8c9ZNt8xj5htJJC1S0SFZZUNHIyfvyhC
M8xeswpEUpFCQrBrfwmavoZbIwhNPp6I7Vi+2wbnUi+zbOfrPWFz19rdfG3p/7C+SzV4nGjGuDSN
Gujg61bp18PHnd/sVkwaJLjgrm3qm97U+vWXXYkPhCJh7Z8hrRe+a9NXfNlEJnkG2CtOKvhWCpA0
4vVz5FYouE6pp2oukBczlivJp+WUgVE0/JwV1wI4tZyUNC10e7HitDkRzhkJFh896XYtCuOGUKq7
16e+1jigUqur4R9BeqcCy394Qk2fEVkDyfleDbJ8bVHoO81IPsgOdoSWvult1Ru+hyK8yMuNcMC/
XHpfrJc7GL1TMoM8dXuH9b2IUkRNk02B4T97BC9/uGot3WtqDkGM7qWylC2T/Qmo7gsayMiE4ohD
aPDdAbktjeiYF0kstxTXtyKivCqHpDl+XonzjF2jEHm4poXrSl9H3ZCnNMkQmb1XPD02a6Nh5LKL
foS8pxIa5QEFzBFIj0BvVArG8gMUEHfYAsWhW0kJjH07Qsd8u/3h/ohhhWcJnUINExhZtVxejTiD
3WbRCL1qFeUAgYAxczRIuzt+daCEgOcM7PN2wOGf07yymKOec37IRSD7nTDcS9TxgcbVyxGlDEk0
fwRWq75lK80EtkKveFsOk51vJleN7Vqmb5aa83JuOHkwprGjzmCnpObb5SMhAfFvLJMt5iOxwpwk
qHjSME5qlMaB90f1nKT5g1o1L7yWx/w2M35SD9sfixnAXITQiL+LO0aRqFnGH/vW8wpkvDSBRzwP
OUpXja1a7YyqWmnPQ71PXv2U/wmLfaBKBFXXRG9wkJP0JjvTQbGdrt7f+P+OW3bSAXwycvXtYxsw
RzhQhmgoCvry6KvJvgISe+HL2JDBK6UC4yMu2DACThsMTs9PmUm7gCycW9dl7AX0tpmvJtYyZ7ll
WI32yUM3iTYL/Tci/nlyPnBajneC4+Wt/gEQ6LNPW4Gf4Uvb2aSBp7ODXBkoxz+44O7NjXZW5kr7
/TghSk1kAS+YzAxQKi1RpOCiAUA7BBmY9qOkDWk+xj2JQlC99tjAwfZ7jDyqKGE94m7RoVrWAykH
38ugeyDk4VC1s99vLeTzL0dOsp23NMH+YlW67xsbIw9Xp81oiMbyM/7ADdk9OboaZtqj6KO82OGx
IprLzWw+brI1wHqamSGOO/DwCGAAjOAqR/zpaIboqfFSa7QcSJKApfW5AoQc57mVA1m20uhPNNrf
CskP/b//hXG2DIwLzc9pSlo2Qe/DLJeBmfympQyJkYq/uSn6oe4rFErgFdoEwmc429LdICJFbVKY
iciYleHdaE/IVGQJLJgkjBkapW0wdOp7bBT6FMIYA/XQUWMg6fR7LlGS6jp3NwBmcQfSWV/CfoyN
uaOE/foZXbn+ixca+GxEX0Q08U0FFWIDn4xqP7wdr9MBs8rKovfsMG7mllSBElZ/1hvDtGZgBXrx
TNqgMvncZrPp36tESYFcY+nvwX2ZKdm4oA4NAL2tW8PybWLmPd2xoHv788TPuX1MODC8X6yKAJM1
xtglVOIdzDkJ8nkmB5cO+WfaIRpOKz71dW8K3dugjqmFfSCfK2wxynbMTs3DFfRFO4YTPVpyH0mA
qszw64XDgaOST+oDVpflGwNRvuFWrRxGfxVMIppwx7nTkgpT9YDCmnGuUB3lSPb3Gw6c5EUFti7u
DOPQ2VB73HumB3Y0mE7AdBBaMkcTcUIlVNG8tAeLf1bo+kLSt4rW2Ysac4MzfFql93XZHINz/SW/
pHNmGk7fbjwAz3APV5I2zpPf61wW5/kFFoeyKCUpoMs5V8kCaPJkomj+hRKsGwfX5Vvk/XWkK2tW
dsHWv+XmRXb0Y6dy8Jbd8pWec97NdOtPym+qWTo/m0Ee9QeicyQI7Ipln9mXdVroxcJctSbjGrxs
d/h4Q0qH2ui6Wrbs156C7iS6BJdX5/ZHeJlNTFs540C4Fq7dQHVujr0naec6wWP4vd9Vf0o+uwUh
XsBjZGHiCUsaUTmmfakED0R5Cp5yFanCXUfo+heei3/Z1Uoa3QV9OKOYg9zdMwg6Zb2Vh62vxk0s
PY+7kAedOdRRo9xfQQHn3KckaoT9BYAMbhU/NSqHi1oSJWY65mCOKZsAyKnIX52/TS2xfQyL1oOc
FxizOUU/berhVL4LGULhehVhdX/4mLuECMH9VS8EanEYPm3k0m0NjaPDju3MkWTOwACAAmZcZpKP
ZwNMHXlRNJloVZkswKUqnMX9AiyaHnnjnOQUzZfkr70P2bCrxrRlsXThKBurfKtm+8SjwFhOEUpc
6SSHikZX82KxBHDc4bWBs61xFUBu4a2zgFNBdehhMiiyMOko/cLFcsIdaMA7EfUPp2AT78YqJ63A
BtptbnFKMxl58LW8ua2SSESZquOZLcKqdP2oectaL4R6X7/qkiOEIIUAkdLWLOtb5sAo/taSByKk
xvKV0F+2Xz06Qz0hz88j/xZNf2OxDyO3hVij9du7BAI3yjzho6AyIQ6ws0BvwxDXnefhRRE/nUGa
6RFRi/ltKPsu8CXA0aEl6ppzMZ+YF7jsPSNFY6I9Kgem2OXgiSy8PWf+YHdqP+4jXwDIpX8+6bYC
PJKehBZDSARyGq37UrBj4RUv5TJRMessbB16g3cK7TDnveaBR4U6iPqgY/3JsupBVTZ1X3GMfDvM
MOv0gdKIscEIjoiMtrAucu+3KOlyTd5YOMBzuYuw+NaBVlZSn2vBGd+xapwmqE/k3HoCB2VCRJhE
hT/hKpH+yRLbm6U8+kuIsVedpEVoBdoNFJjWd9ZH2AQrp8h3VBc430OLHVkCkVU1ef09G3UAOjj0
zFg8L9W6ZSQi6J9f/X/bKRdKs+51H5Mi1g0lplu5o72scjEv4l8F2yjobIRRPwBbFhwqEB2DDRfV
kBK9DRYLVG0yguo2YxITji+w0FutLsJBlmL3qItERrTzFSXw0n6Av2jXWdtHF8MfsUclaAPS5UnN
08uQ7+GJQ1Lb2oK5Gm2fosg7eXi5stc9T4BwVnRNoq6JEyV822UihaZ2LCD1hmuWWbwuO+EuqroS
Jpedc/Ovd3Ft8gsWuNDSirgAOqP944pYv/S4vE16J88Q49rBFj8Wo//ljw/F/ps6eiwXNvKIWwfK
oXRmZA3PN5KYByw4jyGHiZFrxtuXLDd25cNvgKBnxEnD15pyfNMsN5p80zjnfRu2szTDJUyqcswq
ZPPmGkmzq0YHcn49wEYG/fI1p30B/gSzijMEmKBjmxUpoiP03rV5yBCIyuAWcBY4uWmHdL/hLpKg
ZRmeeISDWZ+qGbLvY+i8BDeVHn76cagzo2Xgju/KOaJ1DCef9OXY2e9iNCiWAR7V7055px2/R+10
VG4+fCpyZUUV1d2W+lA0CUY63mD1aTEN+nMywYN6r3LbkeR3cRBdLPQAuoOx6s4PZ/yh++4C5mRh
ZwBDtCmGkS00z4WsBqlljVxCz4yAh1Y/tIRUC2ws2R/u6eCMCGLTvJv3V26jElQYcM817y20iJhv
NXhQTU2yM9nMsDTpBmiOwgZQFs09dj4qupo5LHP9c2/GY6AW+jiIhVYfxUr4/DHoE2xbwHdD0z6l
SY7miIglfwFMXpg6USQG7PMKlFkbiOtjIhKOutaaWX3j7xgHjeYFab52hn1f5AxKot7844cII8Cu
jd+BcNVJGpRFfQlpxodUxJIgMDxy6rweFhgNb86Hh1zasrJF/BL9BTc4ZxUUAoSRloc4KE3XoThh
BxN/X3IMT9i7qRSBk0HijkmAdMgKB996qb8O+nKNTHPoZjGASXYu3waBOgHWpJZerb4mZqoJp7J7
7bk6fCHzad5xjhwDSkF71XSDSr2gkXwrzDEzeoxbIrY+vSb3J3JbhdE7TPb7wuH+S/jtaKZZbsrI
+DD2dCgFY/s4AeX3EDpEpaG69HLk8NwjSmNGa9Nep8kdjT8UUHG1LaobkCKn00ha0DCPT0YxbeNb
PCeYm+xw6+ghrBYvC45lgnKAqmi0ut7X1q7g6tvwP4SW7Au80m1AuNzBxT7YD2E6/GORO/jl9okn
iX0GzdzJXiwGm7w+xJmBO4fNsyiSJu4blYhRathFFfAFDQdX8Ndn6Y4i6dln5/2ofOsr99fpJjKw
FsHfZqWnj1DEEV6K9j7x+gFAHWwShb4MqZKepRjkOX6Q9Gq6NbmQmxhTz5Gouwu5+74npaIP/7Nl
WT4iR9EQatNw3ZPTGsU6tudBKsIW9v7rBfN/+DftlGFwVJJXRteFqPHV+bdLSRLqkv3iKyhQFnLZ
4rju3JA+86UxL3+iglAaTDSIB99B/03ZkXfhIo/DJwi8H/eIIwOYb+9kNnnJT5OVhCD+ZEs6TU0O
+3uvf74+Keh5+aaRaz/wPhOe4uHpBK5hEmAIZJWk8gmqK3CqSrZOZF6ZKsY5bPg4FUpmdpdLTon7
/8R1K0l3QlU3YdlNhjxjhbdNaC5O7va7mnxaruyg2ZbCFM27AWNWwF6/EBgvjEu6kn+z7BECrtau
mLYEHy+vbzUbDVq9r+yvbqRhZJ2ky2RN11mJIWCl0Gv58VxwcYSmxJQQLq9WjPFottL7LR11hY2E
l/UXuw0ughNzkTFBmBoWIbtJuqmRbqKu6EUjxie9yC26QcA0pFJTjqj89kAfAtFr5K4/BhdfI+7h
aKcpGektPQTHVUHsbEplQpX31qDb60dHOBX6GnYpjh4I62b3dqqObr7XCHVbw+d/T4/2DnlKebUq
Uuiby4nQ81k2obUdZ51sFkU50m5LscspjbT5f1ay9ld5zRhB6eweBXtZ5kJKHTLsCr0hAVoUa+r9
qPGEwnBa1SYg0R6ClGcoits6PghorvSNiH2vHr54UubWD4glUKtXaLvc1L3F734ukMmwbLyZjqB/
21VaAmw1w6LfyFzc5qQViNDYDgVsrd0M1c/j5rZZVymolFYnDBLbmdTyoY7jgm58kQJMz+1LSxRz
X90FJ3bj38YG++pAIIlrR1Dnsk4NxM7Wk4RzHjRAGqDaOmqkbBOVpUodZ1azhxXI//4ewZv9Yj/5
GRMtKfwM3FVbT2V4+7PhmjQvzNrjeX6pUfQahk7YLcY8pc4DeH/envQnZ2V7KmuwzMN/wrJxg4o9
7U18X2F7+LPI8puWk9NIG8iFimhBethuSKsMRyWjWkdjmzSMMAZKxBn04hkpRAZ2gFhQPcnkLw5o
MQGTh326b6sDaaLY7iQSeINCyUlGeBJZKVlrLntiGylSa/2pxYlMiHyC+dmdJCpVwv++q409GosW
f+Np0/t7g5pYzg8/iqNi9RDXrOWo1FOK0NucDsBGTUYxd6z6K7BQduKZsttyrb5ZGaCWG6Uo1qTT
IkXzazCxPNu2Q/6pSPw9blgY3HHC8BtvVEGJga9CvFwCDXrNF9eePmDqx7evQIhMegmzaOd2AGtJ
HXgXrx9dWsCgAbMQfXrnwSTik5/4GKlVLMQPJJh6lkudbcKSpWwQNsWf3Ih/DKjL9qozAUBjM+CW
FqDwjAprFfn7SfWMC9Lv/VryXXOQX5SrWwroEGFG3BcwwvRo8axnYt5zjdTfIBsh2Esur74k3k7w
Pai6w9g6mMY0BIWm4ZYJwsmEAwnJXx/ZiVjADS/N7BJZHpGpzVDSG3/TgUjUyOmNJD0LioKXhk2U
T1Xc4GS3l7oLsDzmbw7RVm8GEtJVOvnFnZ8+dnzmBp6UldT8lc/wvAMij+uEcZ6+j5bCTG87bkwy
RVt7IxxWmmzkSZFfqcNwJSYaaXwySVrORq0s7iQsjAuoIcVQH8qAh3ThmmTFI0v7shLyddV98Qyd
Vwx+KYJkIEoKWH0Lb+M3ugddiiWmirNye1iaWDMdMvePIJnWc+tgY9Cfy+3Oqg6uextXYjfjw7VX
gZXrpzgPOZQGJUDJsPcH6/o2rmqWspmoHrAyae+hycWTPldEXyIsK0ew/ecDl7nSLmWL5O+IHaa8
JvqKaSSNNk6N02iKp3txjhBVpZgVEX1hgGbbNCFq0IMoNydKmwXpSwWTXgeGM+sHq0sdUe4Qcgp7
4DHi7bEfgZmS1WwDyxQd6xWCwKIEc5OMjXF/jn+Xu6vJLw0Zy6uUSmzyW3+vzceEzvUA04msFHwN
KTa9NPAPz8PxFKdo90UpPjiLEmxfN9hauMfLzQ4M2dqqMdKO0GileaBEirmX5HkFEWDMEL8MOnqG
yoWi1ZqRxw3JEUcuxxdfoaw9SBSKBiQu3k43WON0ifqxF3pmNiPSusKXiU3nDdGtwJBm+KP5Z9jx
tiYQ9vlGMjqvP1CW987mc553IRLIpu7s3eYvxbEztnGWT/iMLoNBsxDRQL95aIsIu7pYmMXB24JV
nfKiME1S1+Fv+jw2Fc0efKWEZQ4s4qhC728KV2INhlf2R5yKp6Lmqyl2FAFiTlzvWwEnBDMb7M1S
Vd06H70gjLIE1CsXoY74gB40rhYdIedH5E2fy6Aidrjzrvhry7EUdoQhzB9iVBhbk80NuOr/nvcJ
FEO29M1sBawtjJejwum05s4+1sANPRkAKS2FloofBHvwG0BlAqOIW4IIgzbVa5Uot3GObYX9jd0a
8RaGJa77OondQKOkpi/Qh5kMoM2GpSeihszfZFfb51Y7eCu4fdpDah2Hgb1Lm2/obpd15Po3rvZ2
zGNniAlavztkY1fCI9nyND3OWvN8WVvYpR21V7yffd3Q4b5NXMbK0OQbCv+qPcsEb+e9e7FBmkkL
IUpvtOd8PtZKJdHloa13h44dtYOjA54rP0FXvlshqL84eJL8897xHzNvC2UvIx1pAlnTlc9Xzq8h
FBJQeHYcM7ZKwOxOYSOP1jPhIf6qPtkEYORz2huRPirTfOLR0lTstYm695e940ML9DjXDFlOpmhg
mtDXxXPlnIkyAlCalxARu0qSsUxLrpvVskIhqXdk2ZFLi5LIBUEvT9B/Q2Ux97GeaKM0yNk8UEir
/gJ9atg3hZV6mwiTmh1/cCYs5XhhhZ5RdFK3CFIL36qMxigteDG7eSNO8BP41icJI+xcnTN+e0EH
CLekkEkINImvBwAOvwSG1rwTOIfmH4ngpgMC6h7JoCx2zRTQqtLBUBJOLvlJ032xiapUN2KV7PWR
3zm45HnPcSwlBwvbfIyaidxfPPDbuFrk/WqBV0GjTgI/fUB0VRzjqokKzq4EmzR7pY07JhG2BTUc
Im/fgcQNG0JT+NO1q0C0wu5QFmtRI3R/YbXGsT3tmnuHBS41MuXSXi5LwSvEXQssKtXLqws2chFn
9GTkUhQaWuLH27KNPZevB83P4YANxckbZZrJqABOwdS/YiudoBSL7xJKpeVcBluWBq1+SLkKHM1M
+JKkvo5Vw2O7jXveyBJOgjFEHlyUtIPRIcLPK+7vyHI2tJL0sboAjv7/iNmR4c/YP01dE6qcF96p
WYSAuBZok+bGUDrLw8MoCtQfyUnm3Dny6Qe0YnDLDcQFoB7vJsHJmYN1N1I/5aEizQdcZa6ymWpR
Y6db5VF4gyo8YU9w8zMqRLiIha9cNzlQdm4WBG/y/Qq4249onYn5DytrbVyzfJuze566j9HIcdJO
bJfUPSi3qMgP8dtTqy3fTA6CqqmYPY4wGQ5hRBpmGevtJK1G8eThtpt1y3+3I0wm3QhwY+6kfJa6
64RIUxQvX4LQ2TKsYWhmJPNZWN4kino6yFxfUMI0t8sP4nl12vv7vsvKkxlGMCjcJCEVT6ZjccYW
oSUS9DNr/GwyWpKu+gujGrHZEiQzPtqw1hUomvZQkuZ0DMu3A/EbGHOxyXdvBISMwOrMgThkMlhJ
R8miLPoierVNvw0bBsUCCvqshW+wr9R3lXkPKMk6VzDbY3Koeo06ypI3PQ1ajuJDmhcg3V7ek4eD
tceQF/pKELpW9LsSFrv8GNM7s5MCDR+RhQWSQYbDi8czigbRE+Xdoip5Fc220sa1uyUb0tb2eCkT
LJdT//BtvfFMrDycYNAsLh0w7Cj7Mu2Kn1CF7qbYEy9oQpmEp78VGZYwE2Vcb5Q6tGKw6x6iEK57
qsxw5oO+HtZzlAzrN3D+uo7zeT8xi/npHmwLTyjx69V2vAC5/9fgrs0fYhL749ly/wyy16OjARMN
p+5hMXnmuOoedE90lY36UytSqANSiDsLMj01+SB8Tkz9lLAMsvT42KppiNPhvpkOndLMZ5JjEbdG
as5YE7DDStth/Ix+MVkQXPnEhkTycmmdCyjVFvvia/KOlq/bFEMsM83pP9gZv88pinBhtvdeUUFt
Hvbpo7hgvP4mLLNTftR9cHBwbM4OBhg3X4sDr93etmZfn6Jve8Y8CcS8ESk6wuAhVsZzNb3rmAHe
n3QC3AVP3sUV7UjaD6T5f2/bXG3/n3eIhr0f8x2hpiuwO20azCQv1a0wfs/h8BmxJPJ7qqMge9Ew
5mA908DvVj8z7UlbFjhNS/RQq0Qlg9mm8iqSYwpmeZknMU6c+g6RingHLNCkhrR7uwrxMlwp+pln
u8L4M9szLCyX2YWEFQZTJKQZajlJu0aY4spwHSF+PVXOydNbTZz6lDbVIWfnOtGXGh7iLqVwV9K1
cq4uXp9a1Ql33RwvCkIK3MlIZQXwfZIPs3+7qupeX+eyCvtpTXrLIp/8FGie4sBaMim/cbRD2ReI
HHeomIiaCONoQQrT+q4Iq3IOr/zCSmJlT4csfJ5jhBEXjaHnl9oGjgMEfZaG/xgQBGm6OzoiJO8v
WKAdPkRj3ywFVjWgPijRpbWZuBYJU4MfwphhvWkRze5WhQWRGFv1+3J8/rvOyWqUlOelcOkOFR8v
yi+liZ5Py2W2ct3vC3HKjhCkH5sA8ITD9GkVFQIJ+edW0oxeDOcA6kc6gVhTk8qr/oAhVOYasZed
PYxdtVgw8/K4hHJbXhx/ndJ3Q8OAk4VP7At5VAKTg8p9MPnhGSVXmFfPvclq8dj6jtL1diJgkkdQ
UOy9AgzDIGUCrccH4NvMIBcVQD3ReYd04HMFK68s5TUBETh8DDUyWkNsllBWAvNJaJFQQb1KhMgm
K5Iy/r9iMhozLiIrj5sTCPz5+akv5B1a80w47E2s3tppA5i+zBJNzbrwRMoKPiAOidOpRNwOnJo2
mGzj26mV8yHCGO1jWvfbf+pD3OLztHV3Nm176eM4XF0YeHiufIf34sx0F652FRIxCDiN4HGv4UqC
M59gVaG6HCdQRTXNxQ/G4KF8jPQe2Cds61qAyhO9hBcVV7t6D6mqcgmLldGAzMjdXt2jwQ99q6Hw
JrQnnFKOi2h5WIm8lSwPj3LjF2lMUp20lBqrCt5m6aQTkNtt5jAk9MRFmvYJmP65XUMwcwSwIhmk
sQU9KxILsfjYJGnoEYqbHuUkJSWKNN3UUQxv3e0YMyyjC761hZ99d3ZBJ7jg8jwRvhRrWqHrYBwR
vN78bsNmG8bd1Kp0qp9kOQH/JSDlGrQAoUBXv3lieGlyNFknxEJSppGHbMlQhhhimV9FFQ6RM06n
8sGIWjuwJl8S5cnvjY4uXb4NWHwtwzfVXDqL/fxn3trsYSsQsgpF7DwxNlnJ8uyQDtX+4egYvAlC
EUMoct0nZnGmLyNtRa5WrVu2q8BvLsk4me639Jq4dzLwRzpBgaPVTaIhsZrQv3ZZFSxEgCnf8Geo
dX/zgfnHDHhRW3EhGap7NelIO0eBaj5sK+DRdWelDMRE7OHOF+1Cz4jiwvNxdS52LCOgWi0ENrGV
WkJ/6nZw1Hw4ZN5IpGGAiiMLgxjeJxkD1D2gDd0Cik8eWiEvKvYreYyGjqZMf6PpIKnpKD9TzBpt
MBgHFZfefmE1hbtoSKogEzBkR2B7F0Kj55/WB/2KS9f+X1Iaih0APfm4Q+3bgLV4q7jlmwQpezb1
kob+dGyAvbN/Rm9mahxIwY73stMFHSxoIff/KADz3WuEi8FFzmIMjOfJt/cYl9Fei/kdOCK3hfZA
xkW1wDlwG6GwhjML8PrCG8omrhSt0ZQbHpAJ7E+zDx8drsbnDJYGJI5wM8xJIWG6EYgBgn7vNDeB
f9zVbU5KI7NzSjBsiQquDVYTYlsB7jY4saJN+USWLEakE36hBkC7US6yzYIujePlt1GgO3F4ynYu
ox9J4FCcLin8k64TcVFtRFsW60+sySLE+igLE5ldZf6RbQLm7yThchwHI8Kbj8wEWr761LEIMFgG
FE3pLCYf4vH7e3IOOEOXwDbrNhsM8lIjIgO4u500o+QzTm/Qg3Nt8xSoglYNNEVTAvjnDwFaLusg
RQg5YahvE/6ukfOct+aou+6d+/N0kRbng6OdHQJaUwYPFNzI/hi/0m5lVGSfPIlvQmeFX7QlTysy
3vUkg+qJo+W79YFUyPElRGosoxwZJREcSUXb5E7RdyPsbO+lse1NtOdUvjlMJELHdf+PvF3EfBaY
sU75ntgmdv/Z6e4lR0vtAtNb83N0aBlwd6r3+bplhr8FHhHVJ0BhfAEfXrBn2a4Xj6yz3en+Y//G
XWXgb2l/ZoOYiQlgFsJA3ZzVePPmNCYdQSpI0/bs7tTiJTg3kA9Pde1mgWZ/8uVDynVCktXNCISE
o7FKf54LuOU3qzB2DDd0Oy8e2DeEmfJm/iADMjRDedAXLzrPBOSTlipYtFvzNpXacwxVFLx5xHSZ
YUN1g7RufJFgihIqCx8rYPS8oFgJW8yejtRGVVm6B6OYTxoCeOrPJtvGkV7VvBJLCKbv6uAXIxOm
AKqvxzAITBCFwNYN6xMYtc3VoPkKPVQbdX5G4G5nxj6MwNaZYUK/fanXNbfbozRKp/BLAhoA5+QC
C2n23DAJJy6FTnsqFb8zM8YDma5Bu26pXSeormnsD17M5gJ1nbNhJaH6g6X9K1B0c8w4bVJlRQfo
4S0fglu+jyuTc4MkQwdipCsHWc+OJyanoADYSjUc3/ixQxY/rQp2jxQ+OODTzBXGDKxJmH1tajPc
ctaKLU45f2G2omYCRiSwKLdQL3YW/wHF/+HM4FcxZ2aaHWLw9Y04TYGyF5dW2fcaea06VHbGd0Sl
290lc+giEyho2n191OWmTtlmNtxh7aKMfggGnH0PcaXaQYmLJ5zBmiyUxBYcDUynAA363UnbDYaM
21FgDJdclVrStJ/erpfAxbBJFu1uPNQR/oZj9cffaxRVTZHlJ2mtXoSO647m41l3IEIqI84K+1xA
JnRUTK4p9CVTB0m1ENADgSwK1s/pXNiD6YVrgsE0HhPQW/GUKFbfVmXZlyAhE5R82eaxljdqZsZU
vJvdceY5zB4UpJL5QpZnOsXpkDb6ipa5Y9pVitwalY+XJmyqC+ug+NdD1B057Eows0ofYJ8Cs7Sg
PDBuyF2X0YCD/JHlqJZNP5+b3WM/9XaAs7tX/1EktMQusSvgwaw7gO28ViG9bhhMo0y0Xqu7iHxa
3IUBHNVMZoq8R1LQzzBoKbXCj9nrHYCJvMzYPOYZ1XMX/xSk9cj3GW7K0Bi0Grkpd0BLxP1wkHuL
COV7aT5CYD5ywrnlhNzI6rFdzK9GVCvYnwP60gzR+hY412J2V1Vl0go6gRHgTFjWOnM2kTXmpV+r
py6gmuwp8LL79k3klQwibmO7ZadGRr3W0ZtiKR2M8mEhfRgbVQq6fdQ6WJJzvnkfqrysYBDVk4ik
NzSrKBtLnsdSpyXZbSVdWaD1FPBPlxbLCzrD8G+du7lwONdWlSoG/2MkSK4NFfYXET46IUNXleIw
3ESOmIqQIJG82O5S06+HcfYMALiFjLvWr2+6Gzg3D/BFmoVS0LXF9NI5PTmvC407xtWogvD1O4p1
AwqQqS1gfCVBKfChJpKFjI3MLTZ8w/f44O7ivKhc8/rdP891zjZEFNtY32kRg6r/XnbRwdubQDK5
aylRu1wTaCHcuULuw5k7Y4w6jz4Mse8+1J1JUzUcK3oETDFEI7pjCUDrIZuCLqvezkrgKy1fa1Pf
WXabe1dCoRVHuCL3xnqTW5RTDxrAHOmQI9/68D3bbhDPdx1gBNos7go7cBNddO8Ysy6Fowcp/6AK
m36D19j1/IdeVc53ZKmdhsSGxD/3OEbaa3yuvahXReUnVo+WHQb1zLzEwejczJf3YMtqB2+NgETG
9T979p3MT39c1VNwRuFEhc7ZDbklVL53sbkiTClTtAiUThKHP5fQLlogLJAbn7pS28TQp85M0UUY
OYMRAfIFWZD4aUEGb4Oxnx2d/NdLW4xXITLLQhhqE53LnUGjPJqZ7y/JEHe26Tm66gHP/9uHpkeB
iOlEzZkZHg0PXub2vtECz6xi/ZvOtoUcg2WMkPWe0exgv/27SodUC2aGmm2NVpAr2iW4GlENroxH
+7TA8J59siz/ByYzdUU1aGsyltWnC7/TvPpVhh6zlc3a2GWeEt9yuTFLELzRfFhLSLMh+20A3L0e
p7Uawu/Px+Afp4zRdAXENCFX3U2FKQz+gxLFTLOU19b4jxR6Od8m5XjIOCFeq7w6EuftHH8WXKgJ
MOQMv599VlICHHoIgJR/WKv9qNrOYirK3YJVEY/tFK4rpFdXMvdtgPPYe0FCIf/S162c8ZJLEru0
ePUSOUaMF7eShscuNmej4wahb7vj+8HO9Y6mYwEhjYt0SZgJiwg7s6tpoawivqsESDyCHFZqSnFl
fARQ3XVkD6/+lYU8hB9/DdlsiDlt73DeTh4Kq2QJhKNf+pEZhQ8Qo61Rd1I0BUhqS26wUlc7jDCe
bhF7d2qQlXaR0uibSinUBIBDtU4iNLJ/GzeFUURJoXZfTBFwIlR7tt+X1PYJeCO2JJ3oB577kEEp
QSxWYW9MuMCCG+R0e3Ne7D26ghyyDBjPezxK/Yg2K6OusotTrkLvu6+GkheRzJc5L7jJSmyQxC3w
4NiC9NaMamKth2TjmuYFoOevg+yCKbldEtxpkmW7ViU47kZljxXRP7UC6b8z5S7yHiG+Lct+TRhk
O6Ric57YzoEissgFm1SOTAbml9ScW7gEO84C4LM2UB+pjRn+KFeXwTLshpI+WWb9XiAgFIDOk4yZ
H1OCtcgddlTpKOS7LSeMCERNykpAKcm/0iFbU2g10akNjxsNBMcf1gIN/V1VdWPWStZVOGa72gXo
L8xc5e2k5YlKXTJch+ekjYNlTNqx5LeERBiEY6J9DK3z0JNUETM4ilNd3Wfy2Fs0jPmK12ndO9z3
mJeWaiTCbPoHFqe0s+nSOxcQ5QJW7wvpPzHVciOtMydvtpavYkpS84Mf01xZkKXwnyanwsVpIiaV
BYlCfwyvWpvF1bXP1BSwlgH+ELW7DUX+C0y9fz5mlx/5+1k1CyiJT5r7C8/aaIYD1KI8JTWEqRHD
RlkSmue03AYVNKZ6PJhEfM821GoBetmYZe7ofCPjexa0HsIkoeEIhshyKMsfcFDgHFgD8BDhe/iF
wKc1um5ItXCsRL4zLlNmtS/eW6nwBzKjxtrjM/FMeI/sF+I9Xd+r9Zb03kL/ztd9JcbeFTRu+/XD
PhQmceC3Y845456ctixqfbsaIORa+1Ym614KYpyYj7Dg08vPwr5VugdXQa6PcidFhkUeQdodCPxp
U87wUL41fKJV3H7oG/R4A2iCrX3NHzG/RkohjyLTHcO555HVUqBVuFVIaAQY2JIYhEgV+3yF1W4A
nYfaGHVYbqi42vLnJw1brXsgi8wt3H+DRYWgtisno5LwUBP4oB9SX0pbATRmltpuZYZotUfaTWzb
stVoeXe2RqP2kOryWBXvTYI80RlFAC+BaotHG/Ak9Cw43r+pyVolSCpj3FOMUdSavSE9biUGiUux
o7jPs6O4pLzXCn7+1zcvSse8KmfNWiqVbkfMhqm+ExyTNzuCyhI9Nbiol3jEAD9gqwEu3sCZSqGj
dKgPxGJCvSDiZDFaoAqEQ+f2m6bZ5w5QJe/JLSwidmh5SmzFVm5LBqvJXJ2fDkwnhco3uNabxHYy
NAAraZnSs1116EbOHJsedZ4Fu2t3CXPug7l5B9dCn6oVx3xbCdCKt930NrMwB3x1FzQcD5jB2wne
5zx42K/W9AYDzQLg6Edj3Gb6N7S4bi5kw77PgFRY3u+suDemQPZcyq+PY74MBpWv3iGS6oy5RhqR
O4zeAXwvEW3dPahRuHgNlOEPu7dt39NiqGzHou5VG0Zub6LG50oh3qAiLf2Nd3Oy8TJQ7ColAu0s
AKCpzU0ayDaF5al5T0JE28tHt3IpTi7043aF7jExdFd0yhAkD56cNuMWyalfAKRUBVRotmT5tPHx
4ZnXiFdJJC/HEndeNoo45H8DmG8ECkvl12onitLQZluTa2olJADgIMJLLlfLramoV1LzPmwcuPCx
zS1qztK1ZV7Wd1yujwcSIkzTbpVHD650Zqs/RveIIOFizgmbwf3JNDsVVFI+Wy0WUk3IUXuVksGa
Hfc8GvcZ4+yryKHqLNRlpMZFSa2LgvXz7mS2Ixjg00CHgNV+bGMNVtz8oYAkrv8ruo4mgsAuZOOV
e3OdUFb1gbGHweBL0bXOci9l0tXqUFPd80qCOx9DeDjYyG/lsQCQZXJUhpSEHBN+8WA7+GxdXNV9
QXEes1NO1dYg5a08LHM8mVNstXDDK1/dyUM1APBLpNDnru+p+2UPD0Xs8xitfWqMZRi1LPRdDdqf
VUZVpLGsGySgkmCJV0zCg6UZfVAAiqZQRZZAYfjd0NH+83/tKPwHUmL7gh6tuHDByJkbOwB0OHq5
GJ1WzH+uI4hLmmtaRTXNc+Xb07bB6N9A4UcKbJT5vrcZ2bHJKNZDd+2KVpD3zjTc79wTkSpAAmyq
pP6zml2rVqs38fC8e6kU5D3J3LUVHnhVJeerQouKWjPCMEyuNl9cO/ZndZV5EWvd4BL0USxaDyFG
OL6PtuZ8FWLEayxSBy8Q/G83YG1PFUHrbpP/y2PJzWAUtyWVRSjUMH0XsTtGS2HgUdX0ZAwVaUqG
rJIhkLBdQ9JFuDU26OmqIh2OJkfH+gbcH3eCu2/TDeElZBzNIBZ5eoBd+TWIqaSqTJ0VFhnTmCqN
FC8UkInAdF1CXCotnPNdEWkf/GE+xT1dQmUvwnVyxr2L1VlhBWm8B+nGe9tRhyXDfvRW0TIGaIcV
4YqMJyvWTXgBObLIXCsC5idP8mDWwsPiRs3cCKKotrivnyUiVzc0rnBP/uKe/iKsaavkfPpvagcI
2OEA+I8leNvk5pMlHQ57MrGioMdzns6zwxOaazsRRODothJA2g937vd4VjrLl0uUaXLWSOtvvjCb
/Y8Nuyvd2jVzdat94GG0jsiNFNFLdCeiahhfEnm8BMOxv/yTppK6bzxLXnCvheXg6lMhOeU4yMc5
KoaGVDkVlMW77sbJrpZHGqiRF0y4DNqqM+Ov/arLP/pen8P+o8zhGFAEg2uhzUhrqBymYGe+Ue7m
gNtN3suoIFwLX0c2KxHtMz9JUgRMhxc/mkUqdifDKCAez9ZsLoLpibxfweNBdDiw8rnzG36TRmT5
W46+Qk9VVmhdfyBcB+tZCmeY4VNTiiQRKt9xMrz7BGFtKXEpMBLMiGV3tBy1v1ny7dDz9tWN2hvd
9CQK+oZ6lt8OGEvyIYEt0yWit8NbgptAEQb0Xjjvm9bIP90g4b5p92v5GUg+Bs+JSaBy6C0cWxE5
89nWSR5gf+tKglFGrdC4GehV7iqYzOc/hcj0V/vwBo49Rl0EyM96inTL6URfmInD0s9WrbwrXBaV
qMX/5nsYYi1N84Dpo56CzPVd9ygdrvKwdbY8cEsF3KO9VnR9mF67qGyXHdbsKvUpgdVxKmlRnvOi
mEw+X7LaS2ZzSnOfQhxUO9fjr24rNqe3zt1wL64qGiSc0p8FOOcgrVM1LNLsrT+R9RyDcB7sYNnF
QRbddO7kXs1QsAAeV2baXVfQ9TB4r78BVyzlMcko1FbBj/aI8xMRdqO3F1hRLWuG/4B+hYv3fpKf
FEFpg7zmPVkdnjfdVkAn/3Rn76XB8EiiZ4uV7QQFDzi1ixfS55O7fh39I6JsIH/P7d3YlxpAAGgp
9pOf7eoTeCIJyaX1XjZXg3PnRpb0D/q7FiGWO4LAdVlXcjj5ItCMD9ANIkA8P4yHYCMl6ZimuCmq
jPRK1rN90WPm8ZqadO93iaE6FM7qKuSx8PAgt02Kn8go0YfwYEk0wtuPQ117122hk6CrQA9nmQS6
Getx7Hq1PSvH0Kco/Z34pZgqbN0AVVUe6rXvuVwnY3Wc+dI1Mz5079Oy6CaIm6NcrLHu2Sbn/YWn
LQ7Q8VKq82W231GscJ7UVkyS7f4dinY14EFkobQ4KgUCtFnklM6UT+tNQJyjl33E5KepjCuQKC2b
lGwaITms5ysyql+Wl6O7DslD7LW6o20J6I1/FNPPUqokmnYacv+N298FjjHPVIlmEBDrUJYVYQZ0
16XCJ2rhvZNmBV4xC5HD6h1YPmurTsUWAgzwy7J8+fnofgf9+PYCrHZ3M4anMtZceoMU38w2Yyj8
xdpT67N8DJeHGnHm52MPyU7tX40loepKiqlbe+CTVctZ1kukdbmJs+p2SB4WA9slJU0STg/AhkBv
7MhYEOZqY5y7dnc7LU8t2Eha3hiNbW0nVXMRIxhWIEYWTeTxThEo8/ZWQNaqs7kNcsYRTlYZMMc7
V71s/3uhVxzKwswWcGuEMM1x7r7VgK1yIU/m5OQANlJ+xEyIowgcmmW7zT4xWqMUZSBWfWWxNFDW
IHaQ+6K8mS9gpss7TFNotC4A8XF5eWVeHPFmhCKkL1sxjoipy4GZ3n2vJxBcCDu18qV0BzAAezuW
8dzYkkl/7QR6sb39J7kOYPOy+fhzgh7Hl51Cm80CphExqAm9gfJSmQ7dst+8BSJgIP8c1+8+RUDL
sRlZm6OqD34uWmxApM4HPfOE1GE/d8oKXG+n9yoM09pys4aTuqsytq0fnCz5X7+fwuEl9E4/w+Y7
nrA/E9pQCv0gSBXBwi9aGwWUuo12eTpe/Z894wbeZ0BhHJhSxJRn8wTNvRy83/HcKwFz+gUM62wq
QhIYsDjNRagl+3P8dRmgUPEwPe4KMkXrsBJX7OuiS14ml6tMZM8pfxEQCcf2Ui8+4QKHpdXJyus7
SU/KnQkP0eWoOc3RPzMdg5VoAbNxaY2F3lLX1ZIWAiSl7NfVJfuGRoRFUwzMTIWyD663TSgIb9ab
Aq3nu/j9Fugrtb3OJHIwWja37DU4Ano0N4coMavnzGoeKYm8tc6BGJOiCoR5hoZlRfRteG+9P3X9
HsbXD6ZDzIc7OJO3t32kAHRyeNvp666VdQSw6jpro3TiLEGvwNeehoxazqZpr5AU0kdbnaV9rBeN
ifFkhu//iIekYYPQgZbkIpPskFx63Vlwdh0I/SF4vun/um9wb5OYXAkzYYmfXO/iyCcglDZLNmH7
dGgSgng2IUBvjDikEnsF9dtACs1Z5QpGu+/sNCtB2DtXJiKBpswedjYlBHcLvkL75P6RzZ0K13YF
55u6+KSIZ7Bkmqvddb/jyN4Wja/KShXlQZG0WSdjWgau5oVuRQnRUXzub4F0ec4UePmx1ED6blhw
7Pyl5r/UqptoLfwhG6I9LUaivZje5DyjANJY/nTbc2+iDgcQoLFz96YAR1LBO+nd+SkyZqmMbBq/
qTIcZ9XJFB4wWz1zD+uN0JJis71xgRo25fuJqYowlZP2nMUPv4PaNT1pqxSYsqqXB4nj1ocD1Kmg
B0r3BvBn3DHzI6yOywWvEaROw3cRGR1j4WiT2SYWUyDDVIy20ToCBbeO7FrVaPQqfmdIT51qSLaG
3plf7ezLB2AeZ6VD51nykWkqiDnIFGuaGea0oCvUZwaaL/paABwkM3tucVC45W6KXLs9D9G03PFj
lZqXdZx6rerznNKW2b0lUZ+UgA+vaNOn9dVhRthh1oJEBJ3nUP+edAQLcAOYsHoYMMpIdEk+rFg3
3bs8VsSNWtEZFtnShP4mkBurt+JwvZLfGft62TBy1Dx5ITLo4fMWhIwuCYWc8G9AWpAy6zaIkru+
jCg5O0dlPw05wlrsMTOrWDYNSohQge869glYiAUBwpKVbqpS6mc6ACadfrF68NXEeVIYZwt4Znl5
xuL8RuYJF+ve37AYXQVmaFAbcvA/c6l6NZYG0Xdi3eHpqOP+t7jk+sDHwOzw0zSVooTNCvtxd8BT
wpfbYzX09LS6XD4LUiejonooAeBRdU2OZHK9iOrQIH16Eh0bJb5qchnaMPJoiJPrYfVkeoSiJ19v
Md7CNPT0CVcaZZPvxLf5HrlNPqUpbDQFnTu4ea7H9ImWcdizFmcUkWMh3ne6+iclC91LkktOxLaA
m+jga7c6fTfIxYw7HVK6bhyb8vQ215Iy4MKUzoguDjFYpO499jNeCL2DXehEfM3C5QFG5PVJB2yb
MH9wKCAwmrQyXZsXbdVfu+7XzqyDUs3qRW9IOKWrkZYTfFE0JdoxDhsOvpSJ7FrwWXcV/2CicPo+
zl5wPIg4FDKGwoUcImCrWU36HFVsPuYtF8TlXJNh97QgJwmKrPjgmbHIUVxMCXpoyfwIk3NpVbQ+
2N83a+AlnRvgejINvBOGuq35Nk2x9AE7faLkHMzUMhbXnN/RNgmCTtBzjrth10h2M5uneYiSd+M+
GZ1fhfm09tdNtLcAQt3hnCAktht86fuhEtFr4KmgFL6ncKdu7rF4x9W70hZ1lVWeQ3JeqwoklyaH
QKYot5I1aAIKFpq9cYmkJBXFzLLTNfs2aksPx7pcI/TxMvljBy2NDe4IFRibM23+rWg6fSsni3+S
Pl18Su/pWx1epOPTHc8DDefa21LAgTBIVHBWsDBK+/MjBLHtPRoxtWa8qZJzhU6LSsGtMuSPZZbK
I8u01VAbEmBG2+mUBBXLqBhItV0JA5KrhXR6ffrI5856vYeggT9RNO64xaXDBLGOZ4kUuCTb3yOI
B5DTJ0zHhuWnA/7AP/c4j2RXJsuafLjDpNNTytVqjTeVy62biSRXT8FQa102ANilHvA5ZoOD/aKE
JTbKzWgZuMaH87JTtUjc9eL1cyj0yqY3ruz3ArG5VHw6PaGlX0spXQA2VGFcXOdPe5/cqiEh9Lcb
izsy0vQLfDfelfEQxAFDOmtzRAv7NMZpCalGgmSmQrgIX6dc0hxBE8f9Th+r8twiH0XdqPWt/2sL
//qZ+8GJa18OZ/nojenpo/s2CVw0LnsO4bqKdnm5lxWjq180WCRxdJHs90x7GmmELn/w5Giw8QfG
BmSp91bcCGQfSXJO7pEBLLxlE/vJ2wPC5lMTilrAh6Ti0OBpJr/9kiyDPNo8UVtgG3OLQjqQ2o0w
ZJPAfoHHVZodWvttOFMZ4brNrZV1z1cnryK4fguis15SGXR8ZCXRsUhCtzcd3ENOXgHUWorDhonk
jVwe8j2P9BcIAs24jEEbbo7dOk1bAJEbuQ4AEIFan4VYkADI5nRGQ045DGqWaFtITHNQhDWGcptw
YkfXGwNYQpLZuzelDD+XDlDXv3Is6lNsogvVjUoYN+Ak/1x/eD6VjRIR0iAr7mLQGlv2rzZnRcRd
8YLHxyNm0zECf9N2c7hwQWgTnxM/fNmOEMtVcYT6JBFtcPgZ/WYf3OmLAsj8ntaAG1n7ug0kJ8ZV
bBEMohI2kvUnhjbj+vOUuT1BTGWMUgc80kQO53j8TEfVapyJtTNnw6J4mmxFzmIQgc+aJTG13Z/h
MNrr+P8Ksi3cPEnaF0ZsRda/gCmkAwrHKoHa+Ic4+AI3cBPFd8Ii5198eBYhpeCoxjVRUKJbJ8oP
sQZlvrwjVWSXBqGj6AGnz1lXRINUkJCHvSPKFwuBqfX+XaTzSm3AvQ0MeECwcYWzgqR8QFTh8/LU
CWtrBo36ZMcPYjrfdzRbCUNjUaEzzO3+g9uH08HY48hO0v51A73Rry/7xeKBxpy9YdyfvM9s4XGR
wf8FVz10NLbHKYjB+ngWaYB0tlv5AZUxOiE2BS5IIuYRqGRPXqMi731bcq2E8Au8Sdw843ybkA5p
R4lZFuucrJJigGgYZDjettjCHOGUaTzzpi2/Tj7hmU+6SVX7vqsa0uba3k9Mabb5y2M6kgSUPvu4
zoFQbeJok4VA1PwFv77VI7fs7YpRj7eu7d4M+1ws5H8077sRzzyh7vw2ETDn0hkFMY/mKX2nLndr
lRBFgVSZAAvTMQQ5WTv9OjuVhhgpPNsHyT87htOrL/6Tm962tknHAQSaqDkJXE9xOHAsk3zr9T8p
zIIWqQslVzZTBkLvNQWYW5OQV4hKfThJDmB36leGHraqTCb+e4CO0ybrV8H6jyZIlLsiKYHGvjmt
8ln+Uf7kg0qYJeQmwaUYFO/j7DFL3AOIYlorJOoI6a4/PVAcyaiuXGf0uDenBzAIHDdwhisR4dMX
SzDGG/5UxBhVkCHsBhcFDi8Hpmc4YHKveXiA0UAxPH0Pn7Cd8DX5xt5aaBGAdgCqvEefk4nAIG+j
9cmJ0DzIwf2zu+l2E4m8GLY0KHM0mt0/atrmJBRC8J6YauoHK+pxgo6Oz0CL2RqiiPoPj2HbCjeG
E1PVqcDZ7NBcP6phDi7Oa8jRrk+shGbTsRq7rKrkyb0joB8j2QpYfo4+xZgXGU2kVA40lojCHMRQ
B6nr1Do5DyI99vZ8SedxZkkQKPvZNWl5AzZDhngeU4FA9XQHnpKrYSWmeSTTm92zmHjkvbOQR1gn
vGI3RbdItHiAU/0K0LtdRJdnMwYduk4QWuLDN2cCW/LHD5hrCkSOGwzWmmXxMd0EJv2uhLIhDcyn
hCs1KstCw6/H9Ccz0O5x39Wm32BatFst0v4ZU3DeCmOIR1BbDHHDYVfrzx23oGNEps4cGPi8RR4l
blKAgMmAsGUmoSRaa5z2B2cVrJCVeK592OwKnFlr47ETh5r5nXLnyp6IBBKfJ4lLMbWCu+dwUJbX
Gqa68FLyesJVZ/S+Dvc8wJaZmhnz92mK3MUwshDkEtSFf7+zwVjEQbaZhCulQoLl3IV/Hd+C2/M/
h9/kDALXUDblvlUxRL+hPl7YFY6fXHPAeEublgSKeCadzlTabdrZi2D4FVsMbeXnXA9eupdv+01S
IQA2h+6l1CMJj9eYxgUuL0o1t3x0iD+7ALjannFYcl234XnooNZ61ZhZTMbXDlmloTiC2RaWD9fp
L12fyYFxQ7Sv3YBe6Cdv2F5KCQemMZ0+hs6/3FqGGe1vPii11Un+jF5Rhne5Tl1j5Scu3vGnhVax
9uTfYrsV0whFXXH8toeFgvV/ZWuE8FACB6QATMXKqVnUt1s8AwoRbEC/uM1rrzcdR4OEWleBw49V
FmN06dV0qRxkuoNE3WSulDMyOZ45qRdNKl5l9a8vV8okvT+OSt5bKdf2mzocwDcbpnkztQXh/JmG
X3k4TNsKmGjn1zhr5jR2TMT4c/e0ALMVa53UcbEKiDBXFfEFRuL4uh8ZyhFSVw2Uu+97cZ0og471
uxorXdSGbJa/izsonTrm28CsAoA1dyMRP1NYsAAHJ+479N42QqOlAaeOjq6DTbC7UfA1JGVAsqnY
Tz2UseiKHrkVdEiWU0nywXto67o8clpT2MXPxSCgtTdszYadM2UvPjeUQ3vQekNHSCN0hmzcOZ3A
Ytdrtq2cbahFBvLWF2ChH6Ibn64pBa07WbMOgDut/QkRJbjo2qPDhbhFBWcKB3RLarUHmkt+e89g
qiuC33Vn1W8zEqUAXwHHk+1IH0aOcymscXCwTraxmMvNjk4/TrkTjonTT4l3k7AmaJgoTLA+bnTZ
ggQufLaFT4gCtM1C9bCB2SbJlrgFJ89dMaBlZuhCAyindOxG+mPNdtJO8MuLUl+O1r6Oed567nFw
uzi2wkGfovRW7NblfyrcQpERd0ys5BbPoGRCL+tg0nFTY8SetoWMlBgzi8Ace710fYJ2VUEKNpza
khlEL3SMVvctCpjTJlEifdd32Ki0VXOLe/OZvSMGAFKB8yQ4SDzs+rsdgnIHyzYpyabqT3MslAjU
+ads5hmn4OWbWM+XFbbaqyUyamG2PqQCxJ0JKNK51w72kF7g0fgH8mMp6WZCMxwXG0gquL73vE3E
CkhI3Hexvsb5p4Vo3zym1NYmcgmbLM+6vpclGjobLPET8qNMOkzwIzWJdf9/zSMJaliJa0lM5vRY
xaDIXIubF4RVNUYPi33FGWOTEiHZ7f3vCaTgqYNSYW81TnQNfxzo9wae4l/OOtfbAjCPa3s4E/TD
Cpa7yXfq+C0Wkvs0t/fNvzp63dBgch5dcEIjkasIHKO4JZeDpOgU5GV3gRhlg4WqEVBq3LEewZaF
vKa0PtEgk2eCmqzF0c0SjgQNQpaFTMWq9QUSsq/qe56ufuIijiCk4nmTg7YK3e9oPgpWXROyh5Bd
dbqtXAKAgFHfS1rFmcMwzNTuupz6VgX3RyOiNfj7N9Vf9FLbF/IWcfQWHoaAVog0e82wrPKvzQw2
sNIpmlD5EFRO5gJjLNGS+6U358s2zvbqv5v+N7zNMKhiCtWT6+W25WyyiQe+l45J9csPkDL6vI8s
KF3Qkzxgh4zp4eoq5dF6CVxH2gIrOK3g877LgUwC6CgVCw8lnmQ1316aprdkNiPFcgfL3bvuclvv
3eAbqWZqUtaC9aicxYgl+ncZ7kpwYn/sFocHKbLiPWubexnGtxW2BJPTT0/mKpdhlG9/1OtExDFp
FfbJVBfvhJi3FUJZ7QCzlAg/qerDNahgCZu8guzzYgBD33AjO0jdwB70kF4vLncRJJtxK+7DYnaH
RS5o8QnNNNZXCDcs1mj4q3em+65EKyVpOFw+L7IvtLLWPC8AFn8iB/MMpqPrdrKBx4F3MJXo2pUQ
sGlk6Ne56fpOGM6kyCDNG1bcAUOE23KRWBlhszy6iuGSdChgWNuX1Tuu5xTnNhOt6hDFphi3rKgK
SFpd2mqoBwxu+3Luk9TPD/GRMZg62KrzjU5h11ycieVQ26wwyWdLTr6g7krkOzifzxVi8pXBfco5
UR8VdwSh4VK1oBw1KjLEeiUgF3ybhCJDJwsSv2R2PqiexHtft4kGE9XEsAbvwrypcRzhtn2LL/FF
RcmBMFTL2ai7yxJZJxrb7WDgH2+gDvp/0oN2oslTv4mhM6h8J/WjJFRbxXVeKMRnX2NiUVdvAO/k
L/DEdr7d+Rd95Na0qtHJIaUgiVaeGpE2N+71j1/YxqA8uKA0Hx/1RFsRKbJt23satwunIEWusJ8a
2KlrANngJIzmQFarTERrvRD/9vljy3HCiF39c84Orn/0efjrKIukz1XDZQrjnJ5Toc1SlGvwrPYU
gOXlUcJga3zLkallqQdNuSyzce0oJ/075ah3UE5mDTy4swehdOqxtquzZ3smwxIngPX50Pu1JZan
7U0PFxqcGYRCfdBFpiqNAIz6q2GG4xXy6lPnSPVtohLLnllgx+ybOtRK36wfotGQJKcfmVss2GSl
vpuW/2sOFSUhb9LkQc3AhcaSjdfLwfoAVPqK9W7UuSBYGO2P6fyiegZAnPcgEV9WEY6EOgIhDOwJ
jhyZKwT8ed7vilutqBQt42GrwAQytG7kS99meB/y+S/JEeCcyKXxJb/6Bwp/u1vBgxmUrGNzFgIX
Jl9sTMM3R/LvHRY0f9FZzIl2eOmqHN1UYyGwY5KhaLKH14rs1fJyRE2MPWaqV+cbl9xbJZfP8CSe
KE8+fxqDgEdlGomcfTuIYXO4OE4albq6EoejUF5vLFD/zM1p9geQPgl1kFkJcVBZ57K4WM7Dclot
DWhrYWzznoz4nezcjfF//6WuFHrsFkF6CkazazMD6DXrnvgPscsIrYYWkVdgKSWprApEQCoH4vsd
u7JI92S7KqosvosUM7SYxK2ZCh2YkTuWkls8Vi+f75Nch4go4/bfmrFhCmzBwW6d6QuzISovNF/J
cY1FyVSXFy44c9tdTSD+31a5r580COEM4+ZOGF5EgHf/NQgmqrq/oDxNLo5Y7HH2kY16/G/TieVG
SCMFRrmQh6SXOAzkOKJjVxIcJOx5nm1qmPCXeqPOQCOC+x3XZGgHUUPkk0Jvm/PVCmAD2Y5eOwc7
ton3SMt2PqtObEIPgronCQbTYdVTt4+f6c/IoL1PXZde+kwgRIhOHjaTSQyGutM/TO1n4h2Uh/jy
OSkGaj4wymP93dBYukJAJRWPR4c9lJrVoK3DR+8xhiVjIiayQW6BjLwu42hjzxLiDj3Od3kbiY3h
SlAWBNPeYsmBfppNNnXZ6DMLFpjfftxLhfe1bY2uUvTkLED9fVLih9gR9b46gGEtO+wT1X/5F7uk
/tI8QyajKzgbJuXnvbBR1bFdASbWkJWTvALtWh4x+EAnyFgTlcKKn0a4F0y4IcmR9WnbeEFwhGj5
tuRMZ9utgfyh14sWlk2MR0NiqJuV9ubiUHQ7li6Z1crh0gJElRDLAWT9/R49stOPCeie1/fOm4Gn
vQlWLTTMGx5SKr+pgt1/WFV3yftw24Rc8lK5POS84rljuzbGsyb5rivPA7GBIpUkeoQjvjIpeKhS
VIJOaIcuok10a+FNFQRyn4JpqW1iOGco99Z9FKCx1JtW7uh++hKc78iJzC3eI4X0GYDbAdvjGT+1
Ey36ro2JxeOCAQgfDjMgWSDd4Xy5ulsCsx+lDE4hWLLJFzGzyxhCqbRMHCfvk0aWRbyv1NVlI+y/
vPEIPkWx+/Dx/vxqvTAKq397dg/fH0KCcU0icPxS/zyRrPPMHwpdjRlfvS/AG2c/D7E9vXeKwDd8
vjZlf+6HuwKmjbvQf6HpBoB8Ynv1Wcj7hpkoa/WOBZGQV56oyjB5ZgvpfUu3UCw9tymYl1J6f/e4
b95+KPXfOHWy6MIOg0nniPoHnL2hvw8+ZBpI+/h9SSpht6pp9WSjYYfDS5pxpL2kkq/xBGVXmUrN
3LzLxiaKEom1R89vxUiHkbSrKABhH9MTJ85qsuqjHuMT3B1FSGKxZmEg4y9qwf3KJIZDpLU1Gwg3
nJ/+2QYW2ymjuXjka8tglFUPIR1rDxICCTjt8nY65OnacyHt+i9OyMwf5BGadDpBEhPZsua7L9ur
38JoyFx6KNc3WRdt7xIXGFTmW7YmhpgDtzcATXhp5C9XS15ADFOTpOixmJamfgBzKxMyTJ9s6MkB
WswgTFee/BVIue01RUUD+NyUdNaZ8lu8j63mW3u9mlkTSigMGsRxYqTyncTa+IMFF53rW5b7OlMV
FJ0ntQTLZdHM9BN+G3tmJh5qWhLypRvJEJ7a1WS1ve8voHKMSdQzYYaQrF/mv/QBwEeXu0v+a78m
Bqrt8CS8hVAQkF77AfPxPY+R4Gzh2pNsN6yXXbIpmU2BwaKKzbZYcMd1UZ4cP6Ycuim9AXajonIQ
vecycA2IgFidLEHca77Ykdf/MmV5f012J+1RpHrVwznh1+X1Eb4aZtFcMBEChpUc9jtIBQUq9p51
bQ1QXc9olLftK8KpfIxNjhgXApa9qo5hI+xbW5Qn16QUH0DIV0WNOKDJSiRjaRQYBHLEHClYPawz
2iKAux9gECG/4ciyX+IwaYFWHGcM/ffD9h95uz5jxNNzNJI1qeFE+au0XN902NuITDyEVPN9BRMr
mv6Dwc4nudECFn3ExOQQmMiVWuze40i2xHCbSamyRnL8BMbBR6e3I7gMBH1FmZvvtSsexmkLWIRB
1D2coXPie8HHcDs+IO2F0YE5EhXNhnHZrn7UHROa7HclDQNdviiSltIYkrffj5+lA89rucNprbLF
fRVtoS+Vt1aanIemi+S7W6BBALtCRYo0NlAoWthwkft1GUj4ZJkpyOn+K0CxV7gVcT5rfH1j+kll
9wtuRjMX5UNUreZChYKVllJUFLM1HDkXpEBUpzZhKvjVDzD3tTUZWiIVjvaaFoRQq+DvfwmA8bOu
vr9WXqOhyLdQXqGRXP4/Vt50vkua+1Bj1U55C4wx+qYOJTwLT/bFek6UC9oOSh8va/V6iup9ZPWH
unzFDp9xLWbmZpam4HvW9Vn/5yEj7ucG+k8KLwaVtzN2+UBTglkIrN3szHkIt4aih/P4dOrUPsSk
OWK/NzHyqC6w54uJen+LfVa2lWPO5e2JWr/EtItrYEzHN1oJwzYP+kkocQk+e40CK6ZuGgMG5B4N
FAj/M3PbostOBPsZ0m6B8zkebqteriTRPKt9WVhVDx1l8Ly2RP0SLF93uvzaTkrXvPTS4FyJBPQg
uKGT9JJYDMaZtSwyH8ez7ohqrVDMo+kAaEvAc1RHbcIKsIqaUMcyNL3kS24Ni/85j7SLqZu+iC+M
GGQyDhXFdkNHuWNhVKa4eu91H1AbSpL9GsboameHiWEUIb4OGXgdVGlhjvI6bV+cTIsvvYO1GVvl
kQUdnNmjDEuEuO2qYNbpBgpoIFJbcwl+3rSLBJ/PLuxDGQ/zO7M275W6042ximDsZMsgLTUGYbqN
fU6v5pLy0toUq425ezcZ6JMhX0zFGygviQyk5VZo0hEt2kdy93KvSARLlmudiJHAAEZyckRke/uc
DdAt6GHorRK3QJOMMwijLlPZSJcGnKYk5Wkxqibl8rwKqKrBNXiLdaJXVhoAjdTBO4a4JexXUsqR
IS7y3wynDDQpLxtESk7tTPvsfWXBeJnGpij/B86PAcq8qCwUoYlLaY9O+iX7QUQY8GaAy78KJ/+n
A+1i2QSMMYocHCSpmhPdoI/vOj3O7D+48fzyEP/vgOwurRPd0hYwaxA1lAF1uw+fkXCBgjwnMN2Y
fwB0am4FAKCEY6dWcfCO+Cqc29e1TcDfm6yEGz31aPG9053qiiwk9BNkkQkCcL2Q4VO0cwY2oKb5
qb2mz3EybnXshBKgZ5YoX7jn1ZU+jHZzoqT8TMcMkskqmGkPXcdKHQUo00q3i46IKdfEEdxiq5Wd
Q0r9Rw2PnSoDM/yv4DfH8rIUAkS4JqnWfiQOEX92OZy37Ts7xRvdeOzrv8Pv4gKOpsit4JA14biW
LLZ3qAnWdRJIutaLjYChqINjezNgjOOxBsd3uC2ccGWZXnA7368KCf5mrzDohy1KFs7ZqbgqR85L
RBKez1H7z+InZqioZQSgfrUzVSNfgs6GlSLf3NbACX/bwDro7bQc4ESLc2GdcRBLKfOfznxjCk4D
/W7h0BxKqLZ2XpaD3RHlZRxAZgxhumv6C5HQIPeefEzbwOZ6pdpACb3ECG/AP6dHx0HZBK6ro1Rq
B3ZlDAXYD1LLTjvGJaeAH/Pw9/3Ny/MA6fmgOTstQDjqA7IaeVEgqoqi53yFGkJ0adXTGeESoYnu
lfKI5wCu5KTzN8yqscG7AisXS4/cMFJJEzttkw1gfKvffKdu+SvPz+8YTnzymI8ajNPb2XYypTAM
squwuKcEBXwF7FVcb5IOd6LingBqGqqGVQ6E3vPlLmR9pzicEWQ2tsVNxy/55dAuTQ1AxMVPsEk0
zTCIjpBklhlW6lJPVdqH8WqMEzVDxsZM5DuNH1UW3yzDEH0tQcYYG5lMbmG9OVMeN0ECoKnIZFPu
L3SFCEFQ0HlKeG/xI0aiOZve6Rj247qt2T2toLGD7kh5+5zsvAYQmjccZfYR3Xu3XFB9rSomwnmC
B9l2DQlQhhnzVmMW+OR9csfizddfsEkflFRfLOkomcB3a/0Iv1AejIKJ4GsyRxEBh2qavjG6YI58
KUQuC40oj/eSFnq77f5ZywCLxyu0uGMvB6Nf1HBMjgVho08XzCmixsi4aSUlmg4eNlQ35kY28A3x
DIPM9FAZVk2JMvettygXRLGVLHfnLSShwUFYSmuhA3LnaOT6GG6W3ycb7QWcKbgybnId206PFvet
mYhtinGrU1Q4dJA8qa0VldERPZeI8fnGJ7snXsJcAX5+a84fRgf1Cnq6OS6N++fgxQukyK4kZYar
HSM7dIVDwjMSm859gyxHG38GOFIkDJN/H+obD+yRp9oJCxtHKyFh2RHSYUa1ujRMaDbReZ1t/5iw
oC5gj69qqQLw+Siu0dPWiJLMJxA2ayGY925J7vatpiuyut74IQ66MVwvtBrmwFSYdDtELrzoartN
Vr65ae6oO561Dojl8fGF1f2WvAggG3Ssk63VzOyBfMk6y07sOsFzA5EZK0NNmDBXyo261y7d3Yqq
4GzQXELyIIOTjQ5KK8WtQPurg4QKHPF3cF8OLqEkDFnccCaFVAu9/nuQJqVU0HviR8E1uikHQY6Y
M0iicIuMtRO1HkM1cVSAjwtdxjStyqrpDQEfyIyasUI4ZwawMjPz9tFbX/Qy/QGcfba5QlO8R/nQ
tBQ/425sSDFdc8Ly3CxlmwhdnIg2HH1yT875Q2ZDm/yNWzc2PW/0JjUKxR3Mg0cAYrtpt8EYdl4W
gtDmpUPVsNRvMhA3Qfl6STNUg9rt9Ho79WkDlcyVdOanDAzTsLu1c44ZL9m/B9A80luEToG7ycNu
Po2mmahvLy2ru57PFnk7VyA1iEH44IyPLdIwSyiW48N8GO/VFwZ2eUh/nm0EXNIHCvKg8+zMVNxD
79B6eXQMXejfWQdpEga4qQLLGTwf0+9PqwdhFbMVyYlIYQBVlkyuBzgTcd38TUgLp9MK1JHBbnk3
ELape8IkzoDbm1D7lcJu2LE8lpPdtzJkS+o1IukfzUkjTC27YY7ILp9qKcYP8v1B7FnZbomj0TiQ
PJ94YS1iJ9tVsv45ww3ps5mHSX6x3I95N1Fo4CWN8c+WyocaSbVhaoSw6AXGb0oKtOBHqDWEPvLr
bjhNz/oBK9qc4scFq1g8DbDUHBEWf+MaqUUsho5Mq0AGb+OFOkcaS6DFT7RaZUTSEMoTg66vlF5w
zMwui/R70Qr6p1OPDfrQhnTV4AFCB0F0MNLYCzIS62Da0yC5F8WnFjYe3I4jsik+/3HTRJkA853R
1J9aPkYyuZYeI8s2oCjpoHk35P+aebejWoE52H3yA5zjB8pp4w5vEVXyOOhwGUm6+8kPEOgKDBuV
JLCu1drfvMQMSJ7+CYafsO7xjutIVGZ5JlB8OxnHmiPRs5QFG0pq4CRMc/jEqrvdtUXNKuK+SzqJ
M+EmOjX70P3E9JVk0P4nSlp9XADug1kmtHmuDT6D7VuSCiefmzVmPom5S0rZZ5ajm8KyaSlWRQOL
i0gOS0wrdbD5BgoMu5dzn/FadClA8yH68YPvNupNYpPmxAlXLWGZ/ppNg8nemdKFrQCCmeW0jRgM
4cs8HpZUnH1BZXz9yynveM1dIHtwoNbAAbtyTI0mxgSQYcqJyFYfxmv11HIdaJDg9K5jxOKD9lwn
9u3JfenAZjNA3Jio1BV3kKgxLFIKYxo5J/dQfTjxOn2P+2DeGQiX0XxiOXa2jSUZqn4wpNbbPWtM
i8rMO+SkOc6N362AgvVtt7Ijl2ZBYkBQAnQz9on4KMEzY0MlrjWpS4xnkNDT7A7gIFr+lLSiZekS
N6gXX6qXOZTnGqTxO+04CYAxVwYmKdHVzmMyCvF0wGuEXswfxwRoZsVeYX1WEMbZvP69No/7yhVg
ywiHS9St1dX2qME7of65CmxRGxAJggUwZ4Fnh4yp+kgsOLTq9tFp6TZifS45UjvDKIseQpOwjOsX
C7tSHOLrQMIJLG5lsVnWpXjtK4+o/KwkMEDRwHVJqpca7SKHmo97unQg67ZziqMca0JA2tbZbJw7
X1sfoGvfctD8yDqBCvDEayngBGSaRjrfZTgBFgcpzBccNKWd+KSGERRKEyDwhpuE5PCcv8ivbqla
33drhOlpn9I4zPif+NhREr6Q090xFiG7t3RlpOiuOEDCt0VhPd4Z1/wdYygYI4bzmSn6NVK/nNP7
0jCJBYI++GSbwZ6dcuvi0YOFqFL9X9i5Q0gb+2+anxP4cgVA7lCFUMzs9rlxt1LelhNr0HjbYqFQ
hprz79ZCqIodUUBa4Yim1d4M9aZmTiNJtUJgb7TdyQYxT8Fzpi+a5/L2uajfzLJAsevvY9NE5BTs
ZIPyfCaHlnOvCk6eEgzrtRi+kYn5sKqhScobJcBKFOhGMoJ2up2jXeFdJlxStJhSGREjyPNbWztU
G9CyjctEb9+zZ5tVbsH0178/yZjdBlvAmKDlKI+cPMpwihSuxWiGdecvpZKYPxRDDKmx9NEdD2bE
jAJBWOSgju6/Pr+yx4snv/XIdOk69VJoa4d4mdUFKK3V1bjuu3Cx5HdHwXlfxWcH+NyPM+7yaewf
+NDGQzucrE+UHIzrCgLXARxE82SqcqVJFJKWjcHvlRd4CVt+gOignvbS4wCKTRZ7W3Fsg1yiepfa
SLuOaPT+gsNqvS7QjYpaf81zrUIN/vx6redLheB5+UoF7CjKfQc7J8q1ujBa54ARjyajx6xpKc1Z
ZTbXZR0nt4TPK9LIM50lWnRDWy2rZRw/vRcGmBkLCOLpVMM/lGfqsSBAik022EMVzumcAXHkyLrM
+uv1k2iLpcobyOD0lZqZVJurTIHhIHZWNOJmYPE6MkKSZrKfx6/bRo+5ZHicrc4s0DpQJn9LVPbf
6QWSr+WPcLwXf4IjHOpIi5+86q55tWTtAx19FAzCO9/sNtjUW18k8Xx7IYWOCGTUN0OFTvu3VlGT
6J8Y+FfjtlKD5AK4cn/32h+wjMe3DW4dbEvpiT3ns4MLpN7t4TGczanNFeNSoTSmIiu3p9Ja2nnw
YCRch+so8FeM4HjgO3mVJnFWpACNB0NogDHDfi8wITBpLogDmc+gizXPgDw/4GEbTou27ZzyqcwC
Flg876gc5f5buUFkgH0GpkIJ1SiUgu8bxTo+bSxJpHFAVCxoikW/igjb0cL4cBq2hakeeCorPmwO
hlYFyiShd9N2Va72t+/1lSaw0158ekjoAYq2YB9KV4GNoZY9C9unW8QX1+evNgbY4NAgsmoY2bqt
wztV128ff+1qNczJgOhqmEnUaWn01RgEmypZltLMbPtD2QMY9+Q9ZIwwQGUfoN7VBRn8KjNVkstL
tAHCpFpRCQDwlLFC25UZk9VhVJxTha4BCSCgig5glAZtprpK1iNCNmfD5Iyj9IhekrBi/jpCzCib
pzY6khWPY8p/vVr+1DmNWGazg5LLOl5u+LPogvhtgB9r/H1DTR/dC7LLk7NqgGgaWXDhje8pV8x3
O86dLmVxBvgpDfBBHDHfJOFIDPvVXM9cLEiNZegiJjt2HFluTuK58J1OpiXISIgKsJVKIkPcWo6K
AXVzYesfIx+jAKW72ErG0mDyAlEHlIvyfBh4Xx5r2Zl/wf6Dohwv+iH7R9KsXayTkXZGgM74rFTk
ccgtitJKqOC/xQOQWh1IfIMT1NT38rsXvC1og5HqJD7CgiTaOR8ithXBN6kfdPbwT9g/kicOK435
J1b5gZqXy1WKOAaRMgsZ2zf4oNPawKxy9rLA6VZMNEah6gaEBsiHMh3LN+mP7+swbXbM3AQRhH+D
YwM6dsFdpOWqnoTKi+DxgheUO65JOH7kQ7JMiA38/AoDOnuz42J/IorntlN+ghxTNmrk8pfKc6Nn
rl847gTZEJIhyO21R0ZkYoN0v0kHK71zdfHRmcZ/HyYySPLYG2h+KKRExVdD3tqeGUdcrn5BiIyZ
2XBCpuDSv2+7axylPSrL3+YGWrkVsqx0tiKOLFItep1M6w8esKKeuoaYUi8EoyThc07WHg3mMaQJ
zdWwVsao968qClej2YHPIJU7ev/39eg6z4OGKQrpaxV2IxYVcbbIibKcGRq6yw48Ws1ZNm9mo9PL
b0yNCuBNVMf4Hy4KtDTfOlzrKJMayZCW3trj97Fysc0b7A0XqJ4QyCpM+xZvqReRgddrFuJBvYUb
pzAgpTklpK+6HNi+J2yAY+PuZ1KKUyn0VhyNkuzkrFnD0nSs/1Ug2bWN55+1p4+pN3g0YeLxrKZA
k+3dzd7QE+SOd/Eepw0VgSstDFebqqnT7pzleYJb2/0ESa2h7Z37rctLS8f5g8kJa2uSfM5c9l/i
ZauWmpH1oIKZrMN/+cJPxSZas+DmGlmM8/Dh+Nk3S+5pDgskVMnFA1M7Zq2lMwglV0CrByOh7QZf
S3Dw77uMU7UCU8KDyUhOtDD7pTI/4o/imOvpGtDoX5kD7qC9HfxNJze+E7qrCld2AeNE/drL/s1E
TvmEfjrd6IWdinfLAwFW93XbSF2Z0rYoKuc26VDWARf0b9IANC7YqcjSaDn3N4PnVgMKhpSLOX3T
PniZv19IRQm5fwHSkgrGt9nxdy3hqfEky+fIjULU2jJwUd6psA3fEqiJBSCV0JkF9j3ztdSwfcC7
u1pFXm3KHkBNvekFIwYq1+UGLmZpll5GdO9/OGcVp0RdidUm18IVFxH2J/vLLvAM0PDZmBpVVK0l
XksMkViEjnXk+I/Wt7A7Xb4+b2JAYYrPDdTHmWr12Z5h1BA/JPPMT5ZVDS9LKVQiW9C/ovghn6Cj
rI30csM07W35unIvaJZ/mzj+LXAkIOLVRat3hv5tpyE/qAKgYjfjbVWQftQAUG7RthyZyIpME+eG
/rqJiyzuawKE+Ljm4gxzq96qHM+VOxyUQCw/QwzViKU+rynPrq6/oyVZl03MOuJtDmFQ9F6y43Nh
Qu5pN6cSdF4jJID2ObOAJaCubV3yUHwz+JXjk86O5D+b9M1U8Pj65GbxyH1wgO6zZUObLKTL9Dbp
uNaUCQ3xe9BYtRfAxNg4a9u26cnsp7m03AeW3TzSPL+RT0Yj2exqEY5Z3+rLfxob04s/4eRRPUjs
3JeWcvcLrgrDYwhYmYm59IPlt+4Mjttfb40VYsXjYQcWHsZzTvVtTpmjgPzs9PBnjHIHWHfYSftf
ABU9jq10D2EqEUTGaYaXbMrXo9d0R76vI3cCPH2G1UDpAOw4i7Ou60G/ycrIu4FKchb0Hg2vw64A
JUroWPSz1kEfmbewpC/6eloawTMbwgGb6vR/+juCVZeSD9WxlaTg/sPvCwmT2xvS4xfFclz+qrjK
nf9JcZg+Kq5LH04kSQWnzL8KejrV23J1QOWGM6U9/Eqd+teg3quXgMUfAeYcCrciUAN49tk/tJva
9SS1s6yz31WtnQGmzVYo6V/pvp6dtS3ZZ6YSubpmeZde9+gJVWe7sGVoFZHqwZL3Yknylnh8ZAs8
NioyxwNwIJ9Zovu3pzFpFKjY9mS4vHG1Oi2TxjfCb4gJpW5GB8/dgSE6Kd+l6l0PVn1I2IpvePoN
rMD9clrFnOjg1g5mBV+RIwjE+d16dSR3c6d7hAwVreVmBSCtlCSehRSbskkXyn8FoFfKC80X/9mI
+bGfh5BopQ8Boy8cBj6fuA1MznqgRpoA+/lOMiSLPINns5DlVl7dBBJANda2v2k3B6jp0fiuSH0C
58TG73NDfQs18J2W3lmtS0YY9pig8g4R/3al0mCWj19wmgj1snvaM+COur9c0o8qk5CAMpT8BMgT
fYN3UpksoIeMhfKZig2z6xasXmCmRncyNLoxTugyYJ1oph+MdMceXkY6X/NMcBkZE4HcGfkHKJXn
/YikOY5m5ukyrl3qZKaS4YpMpOQKfJ+n221NkhN88LJRhAl/m/EzwwPV9yVf/5hzOpzRH0h7SK36
HVu3BvaXWjw9Bx7byW07kITnkfsc5Sc9svydmBj2gk198dFWY5y/rwaYGT/pO5jyXd9kITZ9zDWr
hVTDj8wX97Omyr3QHoyJMzIJFqyIqkjFeX7rUWbkRHS/q/AUfAJ7wkYUC9Y/avI3nemaiAc/15cG
oL3EXqm9z8qKyKZvYGJcf+occ475I4hIp5DA0c6a4+M/lXAv2DWMHg+Z334SAnQDgzWe5Il3fD55
18ySHqgOY2jdMgsJmkmS7xTTp9tMcsaFo28wcctDkDabDAdWblAdDE8WDpBDnmNo9h9oF6CoYwiR
MbcE5LWGKQqfEx1dnnmIbI22Wtlyx0D8mzXclJ5vjp8ig2CzvqdJs2sgGN7g6sbn7Dq+E54yHSAA
gYPtaWZSBklNzCaYHPeyJ81lLZazXWaYF7xGHJob9JkVSFGr6jrY1uIZzsuJatVehgJxI14HGhCy
WeEcptEI+TNVGEtxDUgKWnXdxBq6Z9JHnJj/SDy7R+MBg/XxToojRifEunUwYi06wP7KlhCrGgoW
V2E73ruIZkk5FzuVhgGClYSUGzdOG66iRRaaM3pPXwfRh5ZJdEhFmSbQLwd5jQXoJ8aYEl9rZupy
fuL/vVophwb/4cyqvgfeQ4pVK+KVqPRG55bCToPJPJiEpXoKZr72L6W+C54EYlT7ysUGpRXG1gg3
Os5Ea/AvR6bmgOzk3BnAf3xNS/dlJkUcY4829jfpZyrrUIRrPAb8CMSesgTNIVkTOUHH53emYxP7
YzD70fV1+FBdn+APihmWiVV0Jy9SOO1swgiuphkYKE+PA9JncZZR7EPCiMOOrsDNiawPMpThtJex
Yu9WiAmo8+s/b04OG212nFR8jXvNsKp8/+YOKMVUkjDz0lcKWy4iAb4xCwZb5kmEbaJ2anzCblvi
Td0oijqiTzuNGjGw/NSnc1FgDvIOZN12LJI2Dys6seZAXmnRdyoyxQMh6yK8GPPqU/PeprVXWvJZ
7Vk0REHvCabnfUkB/OZQeZNFdrLXArh4JsI2nGcIJqnkjUujCYDDUfSp4LvUXFNIx0Ux+Lxi0/AF
FTRLIlbU23OfyVDINDcS0hyJcDNL2AGtjjA4aboyhsSNVaeoLWTB937EdIqZosTqjvn/lBYKCOQF
wQZlE0cOQg2qxi9fNbnm2rcnojSUWxCiFe9O8Ums1QItlC2v1YqbghlseaorU8hPoN7zj5XKfhtj
tXLOlAxE8hMNgDn4hDUBYSOLOTR83gwVglNdGuCWAERknGuu3+ALC40RGE1oqwnw2c9ekloq+Jlp
ChdMT02r8j0FnwzYcz5yWBQd2NkI+Z9WlzmnahV2VFLDv6l82WlAzwW6U7gTllwpheOurSQN2azv
HU9qZebIyGJme+6qoVnO3LilA0Yhb6c0frHpsR0SXBnFabY/zd7Cxlkh/aMZWZiHVp6n2a1kTtlA
xDXHJyChTGPOGl/tfQ3Xlr6xA86lAEMnMcGVQX2kNtBMc8lRn3UUORP9s3BAAihsZ9b/TabPcZje
oNHk/Byv9NGXut4yXjkiJyU9YyBARG3aSv6qdTZtGzYOB2S2jpKoZwUkVT7t8o70pXIo83KIXTOo
fWuxBTdGcGFZZEMqmwgl/GeSryqzAFBGbh+fJn73wPSlOfnyNlXjoDH7J+rMUI21GFZrUckDxOFL
wpXusglmuNumYRAOOYbR2HpdHflavyVFfuHC1uc4Z3JmzexOvLo1UnqBSJiOid897G1KsYl7vvsW
DkM+Bgon6Yf1P9UCr7ncL/NtH8lBXSiO5qFuNcdEwTg0rK67zaZNSVJQ6SvzxpZgjIyArao7ENht
rUSapfiN/gSf7jlKDXYAX5EjJdkDtLT0nctVfPXyIbcR8JOrFECPDz14airktXcXy6vW1UJDyOVF
KwOK+619/mGfpFYLmpY4kuy/vPZYroAj7xH+OdhZJebdSPZK+k5IWbogJ3ieHWehREaK0TBi4bzJ
5Y9+pxMgvUar8Issv2RwWOt5lISKDTGVvvS95I62IrIm+3ieMxNqqMlHAlQ9wDTpkjs9wh5jkQNE
6Q6ZqKdktSZk7eLg6EG/6SxvrHH6XUnsUI4JE1MVcAfgRl9fhkGRCFG+E+IB05JxR/AwuAZUQXgD
reIaaH33RErSxbZie/fVhkZiMoYqVCrV+IZHFBg9Rz/2H74JOyY8w0OkOHMrZTZvwNPYDzc/fKAZ
mteH/m3XozQm4SQ0Zq/gECQRQN/2XY4B4czD7lgaj7SZ8WgSLFGx7DOKE6nOTS18U7eui49ObjbH
dhUUv2EZtJhpmF5ShLwlQ9Bqf/KaQl/4OeCCXuxudhDRoG0CqTFK/QSq7FtzWkoJ4jovN8ZQJ24c
baX66rIhScBKqnne9Iz2yr7xeuB6ylNh7kDLJqc782F1VE3BMfJze7WNWCFypk6MSTHtzecAl4wF
/uGouqLc8YnoS5aPxffB5YCXtXLZtR+HOiSuSoG8JSh2DnjJG+jdHMwP6zD+3dm3EE9cIuYfqPBQ
BSLAFmsu6LXrAzv2u76vCLyoqrGQ8SPIjyk/MWBrdtbjwzSq76RLwE0xZoRr9eoYC3LwK4LCWMzC
HpAvsk6JUPaqNA8939ouIATMsMh/gx9LIQOovZSgiV4siI/VGnkzcsOuuQ/0IhSFJbTSvMK0yp4Z
NXsvvo7cP/NwfQTCsn2f/4lpjXyNSvivoKzXvhc2ALc9G6Z2DaN6BrPX9cpZdpTsHvAfo4Hy6yhM
CCZXkIb6H4hcUS5Tlr81vRaIdWFvgT4pTTORXUwWvzhvoDO7Z8gHNJJyTuRgLhwmULrKeEqGVCHk
MNwY7y3Yt1xE6Euyiu2gtMsWQatxgkmS+Ioz9A5DptGnjuGQ4460YBz7QQQO5kVlvkWpq1R0bhm7
edApFyeQSuuiTEdI05Eh1aUGR9HyleOk34RrxjrppSVuE2Fvp9OFUQWxsEgTGfhMgT2E49jVICdr
yB2cUyWyK8o6l9YfNMHQGCpT5PcfYbR4eTLv24sm6bMq43olx8LdSahRFeZEGGQ2qp1FDJDNl1MW
wa6hUzwoi9m2Z+n3HUUfLJQ7vUx9qyPZRdcXd2NEP5gQhkgYxrFjXBiK+aUsBXV5CO4Om/CXe5KO
xH2SVO7CkHigUw7+w77r9xJ1rjCNrCDdVuWO26GLJEQGY4bW3k7j6jH7rIWUrd3I8Z7cugAC59Ac
K0FnM96VqxSus2ZWu0N5dEEgVemt3HLn7qwjMC5mfLKM6MOeEIm7smnU01VG7qfAMnWNyeO4c/le
ZUs2zi1fk5lOIp0tPaAwtheL41nV7WG3q5+HOeKT6PmREoHc6/vZHPy/3lXk766IFHwqMfPtWU+4
MmQW3C60Qz6JgO6oWeVdC17kMil73qNbeyIKyPAiTViCtzpVAKnMxpEhe54+wNouiPU/GK8MfHxZ
to8r9Z2SiSh+319etAn4lWtxNVbHlKX9jiMVoP07ePC+kkV5b/J4jhroi/DK7Ov88DbD9ye1V+0a
uOoGibLYsMy2PDpy6/9V5lzO20T6zHUz82Kef5sqAg0A6uPUORgrSYNOcITob2tLciBPVwKmSiOL
xJq5NIOa/1KQmhg68gOqqqrbPL8sYFIOf5NCEWfw7YeUs+Q/xQZZFCVhduhVPNh7+D6GaZ4dfO2O
XRhrTa/itvF9PODrJzjX16zllskME8un/KHRznJ0r05L+gpbQzjjAmgEGjdBxofMRxkNwhSOsrjh
DCcBrWPZCyLPAKR3RypsfRfB0j6LniFuKh7sg/nwtMQ4h79K+CDFToHYiD5wXJHF437YfRkW7Ums
R2hpngL92XBf7cDtxv/zE/hZQ9aj6pqzqv17vRlISR7YaXTrGFpbomLky6aUaj/GsmravTGTjjLf
vWVkZrpJk9CDisdQI0mhvWo1xzGQT59foB0e0sWEADCxfOXTslbYuzTamSuHpTYbM3HkqMiByiey
P8HaL0zK1YbBSP7m4emiYZkYpW2GyYfTWHtFpd0aylWSgI6Hl05IZtZUQhCjbu7YScv7wDG7gNoK
y3oDyG3XCDierQz53m28TLNAghznnB1gyky7Za51YgxGQoOqRHBRJ3pIhegrUZGj0Qc54KfYcr61
BvIcf6em9JlXz3dJ/NmcTKbjRcgtgDTu0hHMPD8aN/Z8uf1PPST0iMm3KMcEb0CdjT+RQ1IBOvfk
qMoaZgiKy1tQJFx4SzwOLNu9jZdhqTaHbt8ylI2u420jnhXPIDILt7boDVVEPqSynokVbdMs2mZr
zEHOlSnVOirMl8NV/rZPjHtbPLm8Hv2TFoTjgbLHWzLfA7eROVBgAo/FI6cC6kUXVUBMl9TSOLTz
sq5EEerjAKINHO1LhuxHZyBqmbBnXROIp+Rkxa6RDF2h8dCtgY60fOkQqN5bUDr811fZxgffqWhS
1VQ1a6vb4l13o5KuUcdFXFcKyKehm6A/QtB6x9oSXkqktKeW5bjJSbBTTkmAaRuKfrNUNB2c3Pfl
fy12G+mntl99v/BXrkUHdrmZX89f4ffnTZBEjE/Pzt3pKZMl8mX9e/YXg/LpdgGTvAmuV+1xji2k
KiKsqPur8zLmmMEVfQ07cr0YRcSFDwzGs0wT+S//kvs1PsX9fQy4/GuGMyp2n7dwM19pL8WyDStj
yul/yQVdI+YSMES/LARbOLV+6nZdzv0b6BMds7s6wku1+PsmRdlouth/NVcfSs6bjIGfWK1454OO
e91ahV+W0rVmR6j/gihHKtWPBINlUrG81IY9ZlXPBcDd4Uuvjh4YDn2Dt6rwFcYWvfHtpQNCnUBA
U/1hN02mB40icYw1xQSdYOdTxm7Vj/FArS0epXq5k512+yJ1yc6ZA4tooApuVUs+Q6KeT6ptyIeV
gGS9SAIHDK+WpbZm52Jq8Ek9dWS6dj9aSADm/603xK11fi2wPaVCYtMhqqY+m4YEtXLfpqfHwd0h
SyCY7dscleBkqNZnNBMt0mNuVyHpUm7vL+QiE1mbYXfwBm55oNFd4R2zzdnZSaTuLhB99YZtwODr
e5dZ38zVZFIYEnyZtjsXNq7DChO+TXNHdZT3r/Ea631/gyW9PHJA0FFHiBV6GpWdLl0Q6z++dqse
1OzAiS6E++DTBfB/uGUAE9A+XiZT3iDdy3y4N/1yUIaaqhw1oRzhXCM4TYhfPkX3KCsW/6uBberl
vnQQ0cP1VH82Ui9Hxh4SrdsDS3hfL6lyRjx9MaGsPjp2KAjJBztr3aKUt8zXTQRmckcayjSn24AT
IUw2cM+M86ayNKoPx6VSVs2zFQ/RV9gGfTehizVQ4Ek6808ll6svOpW9M5H8Ti/0IU8g0UPsE4Hg
ZOnVXQfgDcGi32tmLXAH0KJWRErTpNUCZ7nCf2D3RBfvffdkqexyp2Q/8WqM9O+0XMK8Jz4Z8xwc
SQu6Ajm7gn4KpzN3w0+rVFCHB+thtw4IK8zZ+rIgC5dlUreZorm1sEaNGT1d6q72fUYByNgrDRvb
sqjM4ScaDwBCgTLNewj8I5mVov1NebRGbAW664nPtpZh5Finn0s21N33PJQZwMo8/NFL+//Rnz8M
yXoOuPNf+fjFXBVHw/ySEegbvEvhQIhWmU8GGLEdSnZUDagbxJvpbliWx+bBI/M2MDVXayQwXOS6
DoT0gbFxhxu1bhc2RuvQ6EvhInMhH+npLaKif3rOusZg+NS4+owJU2ZDWr+IVcOq9HUuxe8e5Yu+
VXT6JU0kaYkoTrmCUg0m66KSQbQYHdR09NorwWK2Lu8XoZsbPb/D2H/RHbJngRvFx1AtLSClxnH1
D6rVsz16aVFTwosh0/nnMcRewZiXv5Aw+ZnMX3I6n25d/jiFLBl9+bxuPtJnRtlzI+Vz4TgAqfed
AP9H7eFuir00HscF6XEVAFNftPTOmaBtQXJ1r2R9zgKr+KEXu57MVAa2UvdSlihGlDftKfEP2Y7p
HWRdbibKwKYLE0vOdDj0vE2iQW8v8fuCmrE6v06vWLSGxUDRecNNyhfvbPvsnGFdOk/ezqxeBeiO
NnzuOvaDQLYf1Wkmbj/gPbdwaD/9T9aBelJjNo6P1isuL1sXOooQxcJWpDZIyFOLLyBO380dJ8ir
bolORq9rkXiyz9ssuF/i2X8oKl1uiIBNioYeaENIUIvDuagBjqfqCrELxVQXYf5QikTDS7Pb6+tD
za/lxR7c4GqT7+9XaZbXSVW9ERrSM4stQVYIgc8mePdPraBJHcA1EZf5SW//rMTEV52aF6WB4vqG
/M7hcuIUHom8jewSMZgld/de7Dy2g7iodBsf0BCeTOfljR4GVufHgY1Zq+hm+esl9KwUL5u+tvFC
uzkxnSSp61M+VeqcQ7iV5waGgDUCwOn4R4wdP+Ae5zp1axfLLG/T3UqC1cxkB9pN6DqEcoDjBx69
5Q9JJGZ+XlDKaioR3IX+j8RoXAKmJD4mkB3w3rMALANZNxkwxtbgo8Q173v2eXH5VAkUZF+XylEx
8yA12Z44/iWvse2H1lMASGANVSOspiSBAr4otcFROFhb7XEuSkdGV7NZJsYXl2xrHqQNWabTK0Lm
OrUPhhJvP6lnIdMjQYZBqgfeWe05HbaspxpDa3eOhryOJjv3NdUigxRq4Zdlm4P8+yfOZ5jzl49a
vHFksF27okkXOZL4Su0v6x65J73xJWhltZg+qU1N6mdSlRDn8qpUHbSqskIG7eQv+XC5WNEfqpKP
Ar1Wr7Njskrq5zS7AMha6mQCbCttOb1R1NUp9614lLMF4yAts8XkXw9ugNB9T5IpAoRHWfbvtuPP
L0pG3Oto7qKohufwqm874nyVmYW678opEoY5zgOurruyzWuo30D5hPd+a7fCdZMZUsPWDu4TqVbe
QvH+huT6Ar3TfhKnzU2gVGoBQTFe28C3vn26Z/RLkA9cHSLxVU94WmgMF762uRZ/1l0lv8hhNZwZ
dxo3JzGHhkd8vqx1P8qxsLsN09+KYLNohufQXtSp8SMWydpOM2a/aYQfAv078DEIC8xcTXDhsPAS
uSiUl0A4MWjmHYc8xxGWXyx1JCKFohU1ZiJEVzPjJI23O7YBAnL482O4ldbcFRnh85k0vQDtz6JQ
CjBHGNb2VePw2Rk5/Y+V0tAYp/DMEfA2t9pIgF6F2dtgusw3yCuLqjtO7bvGYUdfvCKeTm3BCBLx
QJrg9hYGu3xMDqr9f2uHOcEJqA5WENhLWKW1XRhszOrOzmWOZ6hPXOBB0qZrt4WMmXh3/Uz6/yOd
CUDrYCUTCmBft8390DyiE4DCSTkLNMj0FqKOA6fKYdpv4oajSvnZJKkX8qmEkkL+86B1xl3fFO3w
7Ubb5hsbB6aj7eftnAnnLJv+VT+9/njQeuAuWNBXnqXwcbjYSqGFvOy+pHTJemEOK1yhq4/mTnvq
J4yWtq7llmWmS4t39bExoIORAPpmoAeJE43Jm4ODyI3pNWOTTdk5qFYer6cVLKAZeoRttW0+4UVY
eLt+w7PLRbJGL5nQGPz9sb+fySH147nbOf0m7+sonb/jcsgEpljoanbNXGKYnQvvvI1qZEkct5sb
tjigd3aEhQaKCUumlQZrbNa2NZGYka/sw861ioX5x0sw0yO3+sgnNUQSTadJAwVR1yzx9zOAs5gb
5MVwWtyULIsg5diqGinraM/q0xQQ6cm0zBr0n+zOR7z8K1Yv0nMXxQpklFVZ5dyVxN6RoKhPeosz
xMOIzdXJAAB4tljmo/XDpLiYdK2YF/qgo4hjOMe5Y3krRDLRRp2VRA8kmI7HRWz3Kz9OPJqfOoA0
cs3SZmrneUiYg8aOiGC7BENT/FTGDCoYC69uV0kyfDcHUpwgYFsQp00KRgk2h7zxdpeBwY2V2gce
xFfpZZY+iq5PThWTtE1BTnjKcUI17w38LY4PpJzL6q5NbkaI4nbIMis7kVAleL5i79FIGlfxrbEb
ImGSfP6f0MtM7n7+f5PG7Pz8C6QYt/NYHoL/M15efbA/wmNFxJ9W0ham3Vbak+luJlPhJaHfQox9
AiJHPd3ljQl/tLQX5Se0wvD6awkzjLn3USn1/pBWekbKnK7lEAbwUkhyVW7Dpd6GPNi5dGaH04bJ
py9/XNk9dhM9BLmaVD0Oc/3K8CnqZl6Q1Bg1KAUB5g9GWzYaO2Zg5k3wuL33eJqwNPt7aBM7U+SQ
t/78mhe8aYAcRrjnp4BL1KxZ+VoW9H+eE0v2jRQ5y6HbqSTLd+i98pEK9ujKGMxCzQeM/6zECLxp
uvXt3mWRiYetKxU7VLhSRuIoxWkFcHRWk99JKdbxQwSr5X3c8UylectJqyGWBQ31e07/UPeA2nAR
rrst/x3CGYGNp7ExVKMG1JIp6OLZFhpIL5gcKrIcus3siqwJFfaT6UvkvfWDLlkd89F4YvQazyGl
ITayujwm7RpjxQRaSJ1WOVGfRfKAZn3zcU7XERCKwt4/ho8gWcHd6I43SfVB1/KB/8CaF8QhZzzh
XMNB+qm/l02yYwzdxfT0Ml52PeYlsN50fE61aqwWNb38BGvCjzDpk0t7T/Mv7GZwARkYFuCXmnUw
yTYBaj+oUTmjXCneWiZQ4x51xhxLmj5ita3NSAd/inY34MyFC1yI832vLiQKrFMYlxiNp8puzfBH
vWE74ihs1UM1+qztl/6zTq3PztbDgyYURfQVn3CF5q0Edlnf0U/1kFFptBhTdaYa9zQP8y9/6Tbo
zsxdU7BFuoL65DyvMPGvd1mfnNwxX3BEOfsPGBvR7H2sgUzr5IJdbLbDphKoTvj0XCTKi0XZaB1r
eJ/SQvsXhb0RfwUbyqRq1tbQiFaaOixxXaVkKqAxuL60yZKHdikJ6iY6dZFnqqNZT3+Wru6Zqxd0
V2XHtph1L89NHuV0czlSQw1toIJsLmrG21GAAJArhqnO/O25vImn72Y+YBUXNMSGxZHbnL6gOe2f
+o1VfylyeC5URGv7VOMq53fnZ1Ck5TXFqmVQBWR+aMvjr8OACcggutCBt0/dnzn5Jat2g/ziBSoj
qOeF00HrXpWr5c3m1l27mxnVqKb+6YB1RATOorbX2P2gZ1qRvgw8Q0FQYX+08yod9A+MmsWrXmTe
IrJuEjnV4hP8x/CakUH681IrqG8sxW5PHRVTBaE6cjr9SGV1lSNscNILzJNv/mBWo+BoxW6VlVGy
9Zp/yKwCH2idPICoTaAnVu/jdkVpFchsJipfw9CIxjTdSs0KyBEy/glMIg8g34jZJzUPUlZTYnyP
0fH3zDe/wUvBP48JgQY+dOrW+a3822j9OLg5L4xe5GgQVtlj1DMWto71dmTog2fL+K1wFzc2PgGC
opa4m1Ld5V8ThA2sEzk0hG4ZZdbca50emn/KsNcv3PfiaLAuhYV0Jcr3YSfsy84YgvEZKNCgTMw1
OKO85hqRmoelVtGoufPC6FdY8RlPlLKJxlw7AscEbRq+uZRmkCtoFT+2c2d/Pd02jIYSAOntYrRu
4i6oHC5iBImnzrTQIg5UKUF+HAZBwViWlOAPy9OgKuktU9uWOhFXm18Pto6JcSLZPcCAObT8Xyxu
6RCqb9UpeLi4NHaLMT/Ha1DxBiB00SWi3p6f2jjQwOsNTWguKUx5iuywn2sVc/eWGFFAipKAN8oQ
KM511YjneTurHslMkXXkPL24NgiBiWktQQtkNv/sOxqwpYSG4uIxFcCmdKWKN2x3YQR7o0WxHaY0
lZ0YGH7O5AARrT2MQa6MhlTt97g9ieDoqKXqcbIb27JpUHc49JeTMLW35jl7ytyJ2eiofGLz30GM
HobJyxaatNe0vxsmOKLfTj3IWd8W4ersugN/zgwi195X2IT9/l5gYMTKv+xrf5/GnXvMWj8T4wwT
HZeQggYnCVR5Z8DD+VYJX5+Hulfc6pJcEXtPWCFWD13hkZsXzcKDCOJtUgWtx9rUIy3jts5qCgfW
Ufk1+Y+5O1DnWTIj/1ziV7o6hdWNIlYwSVfj+8gTjW0fKqhlhjyybaoiIY3/vL/toDDgjlQY6+0M
Xz1Ip4T07vha0C+q6XO7XRkN3boHDDD3nAg8cRyozrL//y5tfPpfW3ufrkP4dOP8Dq+9FpGXRSCH
8asiMdIKM9P5OJ8J2MakkESrCweQj62hLxK5OYMwnNJHBk0p1UFaVs3lJCgPXu4wXpjzLtqk8/3y
xmEyPUXC+Mn8F667Lvw2LK1+vnfI8Nkzvtw10pXRlbmKUGEE7gRUSliQQVdhoyyd7QLVod5b05gf
Ly1RXHGXCmqgamYjhekbdhRFHqbodffGAhfxTTVCDWxYEjBMt/vtgyl5GbretYAec4T01pqEUytG
aNC7vonO2cXbVtoTXyWJjMP2JahQCEZMnECBrBMKni7tDGi8Pf42wTuzIkcfScVDr+2uD6/PVzmh
hp4pDeJ499o0lLfFPkedyz0GO875wft8401osHfG7Dtq2dst2DK6+zofakP3yXVme2Ri2sCxWjQ+
RcnpRiXxnkb3MehBEcdWin70x2AjEdr9UjDUjn6vbY7u1CuXpF2TjR4/OJ5kk2UJk/7Ue2+33K1F
87uF12F0ls3zJlB7acEaHJ8FH6LqFTFbipcev2Tvq8maoFSSW06JbWHgLNKFHmvrpoHPhdSbl5FP
oFtolx130NyeBF0qTS1kzHRhH6UlbX5pS5kxOCmghmaBzOhpCA6tryEz6hMVrEqcKjO3MgAonCSW
ZijdPtfEryY9xGtgQafP+H59tW92eGeJq+GEkLEexrUn3JSThObLHGLWDrXZiNZR0um1WPpkTsmK
qTATOg30ksKFrfUI12kmIPcSwj/l22a6jU7carOG2MUmu42MBJh28aDe/c8CfPJGaekM8wfbgrQP
gFT6DXL7II6PksXcTZRd5WMULr6oYt8STxIRvjCBZq5ISWHHKiCpJfXig897pfnmBdH403d+smRd
GqCfCmsHyJGzj9aDa0B6RXQCvDseGRI2ViBTwOV2A0XEzs8H/lc8RUFqehbUO0f7s+HKB+j1881R
ceAMtj0KE0yKbwxC3McU8g0bLW3isWrEM3DR0n8JUgUPiqC/B66TojrwWXkCkTC1FSGFo15EkhWS
lV+Yk5epKWRUnSFwgXlwqgbKWX/piauyXukniRvsGBNy3hBqovKB19K1sNca7dd0ztbIFjFMJned
CLDFIN33vS/XyLwv8hnJ+mpTMpji15IBB9mqzjFSc1vagEtFEvCDmGzG0pz8e5N0OInOZyLxqHL8
OGLwclEhfGoB4oEfmUJGrTFHL/5sHNDzUq/SVjy1hT98dCLJt+i4tcHnHjApXdLbEG2xXAvVhrOV
hqDwIzz4kJyyeFRROS9po0PCrhj6m4YrjgErV2FzlbJU9GCOzWgr1t6M5ZZgemGVXl8oOj7C9cf0
87u8rCl1sWM2pz+V3qxo3wwcIPBt/U+deQ31ZK5t4Gr8MKpniBFwH8zQroNJQoxx++EUn0pVEMRu
Ma13pdbrJEVmgcXxKMiweMoiVXoTGPPJXUQiZx2rx48ZhoUx/HVZsdfioqAcfrOPCpv/H4LHSW4j
H98d8af6ASETFKTjexgpXVUubC9UblKbfv4O2q0MlWSueQtX65rYg7dyRyH9dcrLYWhi9CmY4uc6
Tl2uesIieXPTsP0f2giY/kJxCduktmKwfZCHXRo/Dq/U0YVINe5Y66qxRxaw0bhUDrrTM70CENMp
6uXDZBfo0EP7/ojtUhZt3QoT6lV5i0JdIH5lLE23F8qlHCVIrw7BU4jCCbzbBTKPRTqZ+W3ugH3B
22JMp0qMI/+arnQDuabjibmYS82UC76osSvmJ9g3r/jywEsC7WqIdY+znelCWmhygeZprjQHsNkx
fykoN45sliIUwFPxZR4uLPsMWe1z37v+43vMnj1I/xfDaIrFDB9gje1UrM6UEL26+2zrveqI0AxA
0uVXYzQtGSU7kPCbq88Zh/jbLcqSPKJZdj73bqJA8T++tzBYlQIOPuWV5V9y8I5Y5+IeZd1mLrvu
T+MnxRzyUKR/IhybBygMbxgQ6L6MI3cFxyMFL67aR+MUIht5U86TWTyer/XqiKHjckGTRnFz9tAt
MEP+SbpPkqDo7xdsjO3pfr1tWvhAW8nVl09Noq2geKorRSq9lkIutwYrCq88D2e6ussOgMr9fU61
5qsnnBBrzOBaYL+zlGykeLq04Kqpn+V01b9OKS5CVzNsoW3N7OgRkG1dY2DJ+WKoAazUIOPxq/r3
Go56mK5WixDtI5NIKIalm91XVpSyuAr61+Ex964A96+Dj2KU/ZCPxEMnreA8kKB8O0TYCzbEzg9g
bNcOPlJwBkbynkIQGjzwAVubLRLW+GLXZ9MvOtdyl/9YpR64OyaHySJ8PRI1Z8UT+2Ufcbvri5VM
yOe2w6kP4xKqwJ6mAVcz52TDYPOP6u4ICODv2uLcPak4lxbU4rBmWvRbWmB9GWuXQuMbFEXpD8zF
nhZjqtkpx0SOF0ZK/0KtkXO8A2OemJMeffsaaikKeCwXWX+4AzhEZ5Js0UZgugFRdTNP1l2kf1Ih
JbxlTPV47E5P8K9sSI98paN17izLrgZFl8JLLAP6nZYVPPrvyhkLpkh8ZZpGXqo/QpL3XSJBBD4I
m/JaA2BEcVR9F2vDUYmuG3vQFqXL4NRZb4ijY/VNWOJONkuEbnzddRztfLxRYI2BESaZmbJEtFth
hWjIDk1kHi9cLRGnb0Nmvjqub4za6MXYNnu1sg7gebYESakV57BqDqug/KFlyGaG6qcTQoqSk3hZ
4jdM94syEzHdY+kAHj1aXMEfpAUsZfC2y7eOCOrIQriQwSjldy9DKTacDsgXJF/AFXUUYfZRtMpT
vEzDCjzJHt3X7M/kDYrwIc+LzTTzyF/NKKV7LBHCy+PVE6To2QZJNEz8/ulpu1c63JoLXYEYmTg1
5Smr6MTx/mhQBYry94qlJR3biqArVgufpD669CX9CXpsn82LJW3jyTJK/vyM8O6V+Ey4otwE6ysq
B6JvkqmhMnt7rEwT5bc8MxZQdYlqI50q0clyIfuQBz1HNKc+hg3zcTehf5jb8LCXdmMv2XIsVGcn
KY54+MFuZ4/f7xbNjMYb/Mn9GqEZjOqm8HN+wP5mdqgc1xgloIF8uYSP1kWH0YhyBRJl1+xOWiNs
pDtuGHWVf/mdVzSUwE3ay8J9c6X181eXDOiGaT3IRwW6Be8d+4QwJCOQePfvl8fWxtd9nS6aXqsX
56AdKptnw7iIq1juXx/3RfZxg2lnLCuD1KPiW5YZCpXkKJe9IMnjSW2o7lVWii/sdNqj+RKjXQDw
4YHS3TY7Me+2rJmU2j7q2mpYXGRqAz4X3/O61B7z4QILUzYfoJJpYeLnhvdplmwooRfW3q8pzGSN
C4Dv+WHZkgYCKEpa1cAOTvmH2M/HvtCCdTG5ABkWNkXQ++YjRmOwGfGL7vvlt6VIO8PF+NDExZD9
BFvavvGb2FEO72BAKOk+2eqVE8vmPEA8791WEvMU3vj4lKyDsXNJeES8KI8xGfQF0ZcR3aNEvJcn
e34tHjIOh08mMZ4E72qjPca0QRGWgyeXF3rruUVEtP1nJSBHQ3Afiok0Gq0sILmEXxJLDKlFdrYZ
CQsZlsDzomuUokhpZMjjignGmTI8DGFJJOmsSArz2Pz9+XRDrBNJqc8yE94VI3dP+M9jQrW2G+4h
uVscAy5gn/x6ZGzUcgXGUhUcBtJQ5O3biLZcXpSA4OZY32YOt5b2XafVnxIFs8OprBuoS3p6ttfa
bxDl2vUSEp2pty9KWlHqB+4opApDck0lPhxKSLkqs5dt3QAdo/iFKU0DowyonXrlGkKcomhA0gd8
+1DE2K3kcAfBUeSi1L2qa86C7iy/Y1QjtIdfg+NBGFGSxKuD1zwBDtIUlVRNa3P07mTuZfvb5v+N
hPkglWwZovNtFAsA1syVq1sr2LO78+lIfUg/ejOVUKbXT+EuoDL3n+LgTa4b3Q41m9aFakDvE1fu
pb3KCPG6rYqEmk2luvRDdLhDo/FqntHzXnbqtuBq1TUXrxU/RIvb7D6hfnJnqFKwidzfWSpobnbq
K8c82EGbh3OZSU4kX/HjvouULC5ahjnhwqKvnM0N3Knqpj8MxywU2DfBX9A84FBpyA4Al/dUpT0c
DkSQh0Vh2iKToRNGH+rhAZAbXWmgrEopiddmPINfhEggjQSv01TUdah8n6/gxxJMcxBTxat+Y+uD
UwfB+aksSmBHEj/Ln8Mnoe659C92rmW6UChDKJfMV5JFLl3R2dAJglfo4VXFUj0V4X7QaDLlpEwj
YBgAv2Gz2N6fJgURogFA/hzsEoBu+zYjmGNeswaFHyO6ZtTCwbizPEoI/oB1FpBzbOefPv26smWR
wrZ1rik4x7MsLHf1A0BGFyiPu8UgVmeodcLJjj9eGojDmyG1m4sfQg3DrM75HDuGMyJu4BFW8i9c
i4kU8ixHQ4B0M1M1UTIwxiBgcr3dVSKSPD4MFYGvspZbIHhTaxahM+I6VBTT3q25n3iqX9PVvH3G
31h3sX55LBEz4l+nFrv2YZ6oleXsbOoNpi2x/SXf6vqSfumNB8mxIAF0jpSL2lsFcabLSVnfAkB5
IbVCKyUvUPPAbJI2LR49EPy9ZKJ6GJxK5qYptoBg60Z/gpq0PJTEMBqfJ+YPi5H4YhXFcZAlNjPV
3xEecQkcPUZ1uvtcwwGZeUrC/2vglsVvnRlR1DFOZ10REiVNf9WshP8h/Qa82VjWtaoNyMURZbk1
eobU1fdAeMnxiuB2nfIZGhKF6Yk/xKHrGcURP+vJGhPosNetlXj4RnYmPEDhZZMmvXgOVTK278at
Bk0+tLt2FGL5E0EQGLrHsa6jcC5ZvnkVEViCi/gX14vTFLArEVHfu9bTq96tX7ZNnKOrkFZF0aKL
vfVb41NnIRetaU+qZky8x+8BIw69/JzQUvUBh1Ahs4zgoEcVdm47Hw6v3RSYTKHTx0McQ2wm/qJM
nW9nF47R6Vhf6d87w6+teXmHGAHGYpipBPJQHYMWgBsBAvX0YWZZQJO6aRWW3KEbUpUEALvxZjXk
d2VBJQxrAE+8vIkRZQI1x9roWm44UvT803PXJaCGXkKfW2QX08xDYQ5GdR1RTI+Kc7xAA0/v3Nyk
0F5EYcY6xYKrBxACwWooLi21QZTnTI3VbGKtn5Vk1EdSBcynCCw1XdnepdxcWRvAaDd1wAXjoi47
NqiUBrx/8e518aT/fwdi6XC/QXOzx2JaOKFf83GsVPlAFvlFIpNA7TZTLWFd9VhiD30eAs6WtLXX
jbQ8XaPqVGBuZPqBnJP4ykBtmsp89doeYhLd0A/P1sBCdUEYF3YXgjlgLGQerqnJngn/K1gsUHME
J3GWduD4EwF6j294RKRs1G9cPSJ7tVWB3RUYlGQRbjnqrYKYdlhiU0luZ50tt8tpV9wP2oHGyFhL
C7tv9MeKiUQshYK5XbaaYmUNZG++2MRXv/yZZRq61iWmO6+xgMTwp5WBi8GA+JcebkGQQAM/fpsc
m7UnPothG/ySpU0SSRLwJOKvPnBMa1SupnmUdacVSYQ/d/+uoU818TdMC1ZbIZkS+WX3H/8dLwIx
2aSgHjC6xggGDHuwKCtu8aXQEDZylIv/TbYQZKSq0bF2DnV6XB/1TbCrjvB8XNA61bDHeiiuOhtM
P/CmSDTJBogksZjaiCHwO9sNc9um3zeLZKCzN1LtsO4tKhgmfb5GxgSYJ+uj+ZXzZaf5mwenadps
ZqU0sNUqUrT2hsT5b2mHPv8Na8rKRnEKk/+qDcY6ssxp90Xp18CnVp4sGwKftYq/qnWF8o/No4pL
qreVJi2wLLrNyApeLPG/EyEReO2JaptljqR8kWLbwr3Pr4TOhICraDLri7uqOm+8cnD8pqyqaAln
nT0y7VIKZnuRB8zc32DpuMGBTr0KJVdH5GwCyFsHvt1Fio9eHIiRVOxBXE9V3jnkgQJ/sjAZYswD
I7HFrmRvwUccfnlrm7hR0N+XHH3gVYeaRvfWRU/IMaQdZsU9jn8E7LJDgb0EfsjKzrG8r57v4xgi
EfFh0oOwyDppRyVyuB+1OUCPL63Eak+nhriG2K5bUB7sEMzcg72J1VR4qlzNUSMu6/q50p82wA5q
Jqrp+BWuUfqxZuWxuNQ21sMFPaKZ5fb/DqvyzJN7q19MWU1Te8uc/ndEs09kDsNwCpxtb6ayj9gA
QrW+krFzbjOETt/DG4RmN5SP18dWxTtzmGblXjs5h5rytwKHuwS4mdoYacXmEABN1nEK/821AHMB
CTeRqP9XoRVTTpg8knMhNJA1r4cL2cxGqmL8oIICf9WIB3t26KcUO59feFFJ3wu4Bv4TnyQcuqlZ
kqiAgaxktfQQ3ow0at2qh32MIO4ni2nyNOVXZ1t+2ydLhFxao3bi50w8pTjwZwOeaf8n6/ifZSWt
Nc4MgOj9Sb1yIPgngQ+6fu3HF8hRYuUOBZHEUklAneOmurrWwhA6EcCYh1iPH5u7quoumAMhbxbz
TB1qrkszo7V8N2dWtPTuP4WclPogP/D8G7Nt4cDCOUmoLbEp5AnuOB2+hisByGm6sH0vEqCJi55x
ad83GVpdgCCyYJzIRQ6nidRdaUZmP0duJhbUbimBRcTnLjnu7G+kfvyOxlM6SOMhAm/6ykelAZkP
dtdZvH/qJBUSDx8XhHvtqjVPOl1XdboQcOn9leT59WOkQyCMlw4lNi9Q7le2/8mJmSEYltOwIhip
pTzAicuHbevpQJuqoQWsuDt08JlzgQiFafki8sYnqFF4cQ8+a/ZngnwTh4mfxuudZnDyMVOn6e2S
LMMJMwndA8Q0ZQdfW+urfDNqGq/scbC50TtsTzNcmFFaeKjVwVdjEYObnDncxcUL0st8aU2C0yLm
RFehfZRx6eZYM8+r1MC3PMWYA4O2KQtNfxrBHkTM8OqSMEXJhnlTiNZUmhY1u/QGBkdZWJ6VADjU
sj1OTJm+Pw/wRjoOXG2K+C1C7T3E5PfBauHblQE9YwpAOzovELjfkzKk8ip/2Dy5Q8w2lJ5mX6C6
zC707ptN/GHQeM+HaM/ZLoWRE6ZZfAVn+RSl2HJNA15MQw79s+KJBd1+ICJOehwDKlp/nsYyU+oW
QYH2J13absKPrYlLNTPotxaP2EFPlyknQL9bKk0Nwws+if6epASCTUWHxgmaWJfJ6xKnWadjA8/k
ankoLKnty5ltZtaxKKFow9S+/D+hqHi0PxNAFmBdQap0/8eoZmeZLKsXSpnr0cjlEe4NkEFC3VuI
9JCm5xO26gb4gbV6z2qLX2bNmyxLWmIi4KHVtQ3iG+rv4sMQuysnU3nvGQbZHmgqiwPY8wkXBt/Q
lDrm9DZSufDTh1rgWxkdnu+nCdp5QvUSem7u4qwNg3/WWAF8NiVjOw60S1ne5pSlGzzZ87J3H4Jd
4RkL91WKos5imZj5akbpjMc5+21xdtEfrQt58baEWK43qFTju4o6enprgBeRxMfj158wvtj5pJlH
mAgpWUo0qBUhvCgMzPyGwXRWRENxSlcuoVOba2TT3w+4kaE1moDwXyfxCxUMbsPUoITbaPtkTnyg
aSrjWZ0lY5B+OwgFGMn4jEYfCRFJ74OnSE7ZjmHk2Tsqg3IiQI5FusOF5NQhmThAnjjRVBkjspl1
jinFD0Zm7PHv1PKezb7BHRF476C7CuYQhO6tcMLgDXzJZDSv+MccRNx/MNc0k+j8JL5YdoE1dN/N
a7Kn8yFNeaxvY45N7TSbSxUbkE1UgDCS7FAAB3mgeTLgO2uI91U+hQkkT8Tse8JzU9RWnKxYjcIy
frCIbdUQ1ROLKhafiL9m0JRJUPFt8/coaDKKF1nrQe3xf/xiRXq+Aa68NSev+spKEKmALsnjZ+w+
NDqsTG8lFGTsrM15uBXY4OCIT4wnL7Cfknf7zyVq+1uFda4IgJpICpxR6hoVSJsxOKVhRXG/ufDX
1FKsO2xLRKiucMJXkgfMXt4iqFIvJfdtheCr7J3eXJJJ/asdkUK6nCw2gAVguVZFK/EniuPEavt5
L5excgM3ZfzCk8g1VNjN8Pcm9J3vLujjKFxHidt1iRutKqj098oyL4r4mM/FNmrxL8mbDUL7Hd+V
YAFy6h4ecE7QYY9JZQ2OPOuVAIkOea/dxhg/eJRvHr5rf0zi1415HjH+3R/XzoWI6IiUeprAwz6Y
xIfI6ADENKQweXQVa+eY2mynoh9laO9g1fIXO9wtnyY5HJI3w+uCIQ88YeSV2NiZFT0y84AwKq6A
O5h1gSLlisxGkY3q+jdiAp24ExaafnWR+E5M3jJRocQLjH0g8YDFAN/EQg0VXaBBGHyVAg8TlpPf
PblaOzcq79fUmmBewwwWUrOoaOaL0q2wVvJu5kYFqdb9kbY4kMm2tp0M7BYv7MicyItr7DyyGYcI
tLjVk6ar+I1PRD5Spt8BSBi7Uh/woim7BWz6akLXFCjKNv+o715rtUfA/mpK9v+xYII6bTGQufi5
dSFot9nvQLeOyNubTCKksAuNOn9VeOv/NO5JBvp4JwR4OARcSRmp/Pvl5ywtVFXe4IzguC9xVJ8o
nJy1olcpbdJZLyT3B9ObTJKY4wFeYp45JCjiK0d58E3+iSp6QVvW9tXHsdLbT5CXadGRox8ChyEW
d5Xfd/yi031FZ8CUCnaLDEAnRJh1FTjLGpCLMdrhWDrVBDm/d32Cslc5M5bUoyE+1duC4RHSxaiu
i8ofDVmjkul1S8OUzU3tGm1r86mwy7U/rklB/QGATxXTbwuQJtq69fWcKjJRzR8qteIw1IIP1Z5M
MoXH7WvA8oSmOAUhMtzXi/gMcTUE6KIWBI13OfWmHnI2H2awqDPuy0DZLZio+tuDuxn5d7hOD6it
gfSZ0pwjCFL1ylRvFdd0NWWWqf+1FNphGpJj+cH1SOIp2ECZRXtJ+K2Peyg8L/UON0dJfotpp5Gv
V68rhaQUmnwc/3noo6yLB+0AhtcE18FI6S6WFHnMbIWCq7l8Us/X4wsb8KhY156idyuGhDpJfu+g
ntQmxHksA3LH38l/L2pEo5WilobXg4KufLq5LZmMcxzD0D9YNzaEAp0i7ajZooEicmjX4z08TROD
DREdBSvZ8WndyGrc3dyLd67Cm/LKzYizNCntwgv5Aq/t9CRKEXDV/SkScuQRMa6WwAS0iuoD6vxh
2fgWRO89ivPIq7QEbb/eU15cguvZYTq452w1TobLnXRdaQg40baYRqZQz15sJnl73KuiNn63lLm2
9TlhBuPCaAYTmcC2mtJoABva21vRC9wo+DwhMFscjHtRVYQ4XSNUgGhOuifeXZexHlnft4o4MvO5
5DqkFwkJ5B3n4ORsJb2ZLPgvZJCIlGeEcE8on192qAFJgnSI5/vo5HffSWggx9k/1ILiXwM+emNB
6jwmJG3hPY+77ixM2ChsCgTebwptO2YatZRIWC1QxQfsef/0QF3f4cYoCbb0rFC6jqXWVcJJ7QMu
famRSFMsXJBoUwxm/ET3AjfXAkre7CoM6dm9pb9098sdfkSivKSLTMVtikZgPCOwfmAC/HQag720
QWKFbJlQEDziglyx/jSf2mKleCfgiRafl7PeDRUtzRr0i/RCCRwI6W+kQ86/tR9q5+Qk27wh+zyY
IRU/ul5sb2ylRAKChjRSHpOY9eGYfUbKQv8yBjXRne2BUH8KusKdL04e7B2uQ6NzB1NfOlBVbdlX
YVCcBaJTk1I9Sz8lN7q8Qf7jf/YaEsIpdtw11ejKT3gJEKZkEmvJxzOwpG9ocwN8ZDaZSw7Y0JnW
badhz0G0xNN+syE37g4GDwxm2K/RlVhH0G5Ic5qvtmhpl5bQMOX4TT9YY3cWnP6gABc9QFCaMTpE
ZV9DBlcD7tXtUdNqW9zy4uh/7zqLZa6OPfiDfdmc57p3hGMgIuO3Cf/EwAV1UraIFmoxMTAE53M6
lNj4V1jwYQrkiXlnHepCfaZcR2zjqXApegu3+oDn28QGrSDZ3PEB2cPikP+nuKlQ2B6j3CQZnKXk
B2HCR45OY2rCHrwtHCsyyiYg3Hx5fOyZJ1BInK2p07CgBdQlrSUv5V1qiGvC410tkkK+56dqhkD+
wPD79shYTAHYwnoXgjE8f+HXT0kkL0jHWhvbP64wqSKWUI64IrnLbTPCXaEexKB8VxelGrnXFLKy
myR5xdFKOCswJMznxGMnagJnwgj5ciJCTpiITrpBMLfv9bEyETUq0HG12tU1dLF508Q7iVwcuaBE
tx2mGkmc/7niv3CEgBY/OY1tlNmUfgQUie2/mEAvrghZVfZntj4rlaR3gUMrwj3m9n0Ce0M81eqv
Ac33245eujyyznQq0cqteSJUAdyc47dfW/iKd33ugEAwBw7heOHBxME9WN8AQp2B2OuPS3FYqakh
mzykd32WjyZHLBDkni0LUz25G4i1SDtxkqZK77pG4LFW+MnnFYdwzGuJOTevZ0MtNCx9+QDR6gdt
WbT5JjBfdXICEVsTf2wDL8lej3Jea/udETqADcnvdg44A0Y1VxEPKtohKvCdoV2mE6UcM+IAnDSQ
K7cdwaVsItzEk78NrxrFsAeuDaxtAbnSEcv1qaACOWLEN4xPon062RJKnSkFiox8gfIyIObnLNiF
3XDfuhhY0+YWase4Zc3RmdnEVWhPI7B3DfQBV+WFrC2lIf40I9lNog0FG59KNvuHQPepZqwljqPC
oGwEf0yMOH/lAjC5dnt3YSUzD5cVAeXe3CImXEl1rWb+M2za/jxapabM++8ASfvkVTy3YKWSWD4v
2TArRuBazfpeYfJQEekIvuoRtkTGp+rkUApaRLFx0OTkXUnMkYJd8ajUwbo3V0Vh2qKtfncIch3+
jjiVnakLuXCs27CXaunyKLRVBMWb3mXL408CZhOn3aEbKWNC6Ac/85cl3sZwfeTKbBoui80su0Lm
zQMPagfB5i8KTMfk+1MKHS5E/a9Du5rsHLclSPCdFI5xfMMariJ3mjA7gDm+B1mbt+RrnLsMgtuI
tA+XH8nOZQz47BYhcZT/4AI12ZVpLiybJxJy82Cb29pK4psJnHclI5f6EANesUEau3vSplRECn/g
FaHIlsPowubUzBQsIWd6ljj5VolVcrG4BZwkeowSrIfj1Ezi7Okz9EsHy5DsjFlzRHrFwDQ9q8mo
CSz7ztCB7EmuCCtzHKFKwFWcy3SPVxh/nOSSXGEogAiWRgcDIwL8dij62C9K+b3egPOrg0VCebyj
a9ErH/V7EEu9nLo/hnD/veWDmMrqyy6g9bVS+0+xAXtww2GBXlA862KinJMLO1oudGsrVtx4mfOt
2h99DsjQzZgDu20eKwq0YJz8LJ1NF4fAf2NLbEw8tS6mzzF9RV9zBY3fC+PCJrBIbcpK4fn09rPD
T8121fsqFq9eSQf/v56HTrVAscNVBji/jZwt//TOOv6J9BFeYpcm6F7N+GSSZWpadsMpoe6AwxFI
BDQOyPuxEo9jlS9uGEOcZo5BUjXEa9OfnDCN5eAnXwWjN6PW1yKBPMPa2zpVTpy6IY1EpcncvDRW
XW3sWrnd1mKCXLs1FpYEmvSZWSdWqMMalqegekoEd8uPTyh+9KECcpl75/jcuROoj8b78+I9oHf/
h+xgmGXqDMCWTN4fSm0oym1FWtoJlLS61A4a8tbygMeTrP3veBIKXJmGW1Dj2ZfdxeP7LsUV98Ff
VVXZilTpJ/2lURibak0T49+In55s/QtxbKn9cDqcxvBOGOzjSsqtveAd6tKQjoVgS0LgC70+pXUc
pzX5eIUIWBdCo3C6xpO+WyHJmzZCKQq5KV9JAmYuQs0izv9t+PwUVUufv48hwWC+I5umWPgLb7XJ
xT4aepS6yxec7pb1f2DeU/RCqKc0GnI1d0AFcEAztNXd6YRi6aQsrTqLg63XuD4pTQ8igBMRfLcr
k4HEeJR2RmQvQBBolep880WWliqLfsEecW+6TfPW/CV8nyS+m86NxS3MgD6Pmpycc58xCRZQP14r
oVjWBemlhtDDYcYR9XU3Rox3F4Y9ywRKXpZlwYPeVBsJf6n6RoAoKruWTRviyw8/h4xArVBKxL7A
mDpSzM3eh8Oh0oMgSywKUaLWerVmCuDqP5WT1rdlPAD8KZUXHl3GjVToR/u/oZJSRO69/7f7Zoqz
acORaw1Q2wR/LdPDim0A280lmlY9vEUO6LU1Bl/Ql9CeasZiDFm2x7ejBlLeNfmZQ/jL/gqXlHli
8P/q/NFwViMwl/Ip9jzwn3VeklRWkp++IPS1obekui3L50bEio7I+B5wRh86C3ilvWFsW9jABT/j
OJuMIrvQaTOcTErbEc41IZeN+c/dnnsVuxYyUOY5SH89QMeyo3uiBHMtqGwvs59DU1PErrHAuaUc
J/LSB0AJ5Tag+dELfOASkQcLaQbcHDDbSs74p/UeCSS5ZRpGEe5zzAUBLUSaGNdRop/toEkNxRwm
F366kyCOXEwERgM8PoVqRNZFWQMz+JNXfIvqVJnZUIHGOxCwMEkILHAoUpd2kWKkwtg0GI48C4GZ
H+6cuYqUQf4kI8NYs59opYKymAjNfx/IXnPHheZLclI8bkQEoO85w8YXzWkgq+wHPfrW8ttDoThl
sXu0w/1LWj3CJkV7s8xCN0e4XTObYlCU5I0rs+sTrD0riioHR6s5tBzMTBbnKnGlxDdLp2+qOoUP
pqVXsiC87ZqafHuBFoaT0Z6+NUJ5EluXMActr7GurazzuO54FUw8CuRZtrIW2VZMtODtSCSzCY3t
P7McEPH/3YUM3+RqgiMy5BElzDTLBuRmGe4M8dN5j7raGkhdNt0nkJaOhV5UtZW/tbd+sBclOC8b
6cp5e7/zapBtfGTWnld+04sSFeSa4S5bbHMo+cGQW8UR3Z73Nor8we8zcSzz6UmTsigTtvnEJvtJ
L8MbEXn9ZaB/frjzUlKx3PRbSCtCpyhOIlcruedj6ia7IpktJk1msWW967D5F6N+wpd4B8JjsUx2
qw8VPnCf5QedgRk4t29Kg4c4W7n0hMYZXLEtiEeNvmvmlUrMVRYxPW7vxuYzKVx9LnG/xh9K2LbP
FRx5qMDgwTpplz4y36EhoGW+1wo6bw1BrRAYNYgLOds/s2kiCu6ZDHutFTsH/lj8CMklzf9AS2C9
7vZTVO4++75z1zVU7DZcROx0/VBM7oMhiUEsEmcrt8hsR3NNKspB+AoFLcD369DT39a/6yAa2aHA
3dfoj3tjPUp4Uv3EFkYia2zFfZSveg5cQvp3vQACyE88GFOkSVRolJR0JqsqrVVcsRtsls6lcZES
NrkDIGQtR6UCADb089L19nojjwGAgMicwp55RWb46a9EQV6RnlzZLhe6NhvxUr7KU5JzAOmP60tW
QyCygG1JtJkUI12iLSupUws4b6VIbM5OGaudIdlGzRSeoNG6va6OzQrXU4VuXGACb7Ef83vuTmI1
NT9OIl0rNi5pO2Y+F1rxQP/QdYvjILTQnG+9YsYA0zjUE8b93LeMYpUHqHEDhaJfmD4NIgrSo13l
shN21N94ywzQc2FHPefYgI5sGUlL8YHAh18gV0cSBnAGU4+pkm41uDgFG6XmFaCM3esr+NamasK1
S9bgjbi5yeWeQePhcp3PzQy5ML8rLIZ8yWLZgQT77vt4EaJZ2pS0lQDlKapxonbw69JTddK4zoo8
qoGqU77TQAmfF0Z4UARBO7LLkYDPcPqp30ahNnXG52c1X+WUwSNa8Ns4npManP778F7MdnflySqD
JpYg3OnqmUqltaJl2o8D618BYleCgOUNSVa7OTjQh1c/ihZUvTr8gXSqSDscwvx8ehTe8CByZYJ1
Srw1YuSA+bUKbVv+L6216/832KnOUIxyElyu+PKh/d4J+H9qxNH0xLJeIlxngTZQY9Xl53iE04jV
5GF9disbFKJsRidt8lVTnRpJ5jlruUrN9WvDG0tXnZceNYgsBmiE8p/8vUSlL7UXb00JBRE2AQun
x8fzTFO2MqDzvl2Gua6z9xXZLr8A1jBJu7l3Q7N0wGZ7UNLpbXiF6OcU11JYj+5HH2PNWlW7WqRR
lTiXK4bmHjGx29NnZuJxb7dIESWiFvOYFcS2WrynDI7Abb1AwNTMTolexnbNTrNbYz1dBn5Etzcc
xMRG7FfllcP/6w8+XwMA1OemsVIT06QbRiHba1ANjTLzJD728IovDN6u0WD0MOjVFr+QznLrKog2
vMUgvgGOPxXwr1oTOnPxdDawr3ClDe4C8UQrzkUmqL6/boQdTLHEsespGYqyb1R/u0qdXN8y4mV1
g2T0rlTKdPl0D9U50IzOwzqRBisZAuhd6jGMAR1roVNAypKOYm9U+zvsRCo7BxubAD+Ogi74Hklx
2HisescmKMWS/B5rcm8gsvBukK/v2HlxJ+xqu3oMXpL2e1FF1WVuUvi05ATJ01ydffWKKX0SXoVI
Hdw4ii9lgegjg7jYiI7VtW/ex/QjraIPTCmMcKwHYtx+u+Pu04naiqpCPeAqzUyG9k7ocM4pqXug
fk2DrYk9syah6DXFi+UeKRgC7NzqDXSS3Y9u7BuYzrJgsMygOX4WQ4IivbE+NOhNxOxAuQ83vlAE
qpGnHYdxGeWzXdHCNTtUzMt8PLeqeqCM0SI7h9ghw/d24zFC5Ve65arsU9mYZHvNb/jHtxtLWTnF
rmxUnpqgAIvsO3xgPfBoNjM71h15s81q5IuKBPkVI3cGbwHR0E1k49Js5Cu2ymY/sm9y0L3ZznP5
Nl6nCd84fOiHKuzsepIVQ2ZdkbDjZcwuMQEjKgnMkTik9q6iYQHm190rsk0Zts6+75lU0BnSfZTE
fM+fjb7ykwbbiTabblePc45NfVbJqQMEfHp0vWNZDcsYBlGBlwiNVuNFQ4t4YB+qZSRwAELRZm1U
JkMZxqhNhwpvdWUGjqP6jTDBf6gp7A1tNFFyU8+xPwBFyhs3u84VpJ5wC+m8pej7q6EKfrGlCTNc
pp6Uv3qnfvjA4AU/ZVlOF7P4inhMB7/TG1BzEzkklqLx2U+00m8QMZ6VLxHdicpXPtq7txY9oq3Z
Jzew45Wga3qg5zTQ7/1zDri6ypcSyeJRCZIYt8FKjL1wqTxAnsy5O4e0BiFQ2zE4fSeCu9Iuq8Fc
cGd34NxPr4ObBv8LapraX1hiKzukkueYUaRB1m98jmj95qWfTM8atECyy4B87sOwruyy2klVm40P
pTl14ErLsJSfJEbsZo+VYYc/qj7Zr5jFcNgzJwWhHUAkWWzOH203xzsRoifNFEMHHPFjWubgh00g
NyodnAiv3czowS5XXIzcC9fDGIoS1Utvw6xo4Cyk8rgpex/btsCcn8hPhEPqNj1Za0zvfVxWaQ7F
huzN5F2GfacIMWTOQEre3qCbZF0+HB1hsXvR5ctaMPnHD2YSN/58E/i0KFAA+rUsXVyQDCOeWioI
q8/r/U5muvF0VWPp/d+IRn3WdaaDDOOgaGJblPBFDGys84krzmHx8RCnU587HAb3E5C3s2Q3iqiy
u5duSU2bh0FBu0Zk84OMQl1k3R8PRuZNE/uTy69f1OBTuxvJZ/0DjVJiwi0B8xh/SNCZI90ePrSZ
HTxdtnCwR9FKMdI05eJk+7aeS+yW6/Gm72bXZpJTFxVk943q6IQNJmP/mE8/3867zZed2oymHfKH
CGO95AdyXmOljF+YMNH3TMWiGsorh54lT+DCDWy8lCR09n4GQs6N8NPy13Kbf7M2cYXtPHftijpl
Wl7Zn+z1ciuSNSe6UQPKz8lvAC8uFCEvifa7K4ccGSetp2MeqsfiN0slUjN2Es/rYd4+pDghUYz0
0DmlqrF8oAaLXcAocfnbXXEMZZfCSXDVhI5qgqXcJ4ZspDdSDQZ24sOjoQUyh5rOEXkMxit5Undy
2nF1mvNhL4BfyHY+9JZ+RPmbInKvAhpjjJG7kMgKbXfxV1iUaQwPkm6OUVIxRkN6aEN1qLixwR0X
xNj9Rv/UImWGZphKE2d3D51UJdn2RdXBVZCdi0os3JcDDl7rYt8BtixNreFjfduFMSKAUnCmOh2Y
TjIZtJtTkTVc4aeTaFi6jBEIobL6qGg2xhq3doEBFsI7eynVwFA27tnHzNEpEio9Pqi7H7iytGY5
qmKv9u64FtrlQb0k+7hB9GztDATCzCibSU/D+9BLz9qDQ3TUIySE4vAIysIiviqz/VWwWEMqOQ5/
UaMEHToeJbeNBhya9n3TtaYq9fJH1ICVJkElGrh0maRx6XIQcspBwH9jkkC0AyI5nh/CSFIWGNhE
wUbgjx9JsJHHz87qaEuLZnOAf6VN1ALIgP/2mfczkwEsqDNWq9Nsk1cXKCKJ6ykQSGL95VEjMpFD
FTGfqxy4jfq1QfELc0Q6jEJ8RXGRThMEf8P7m2ii7kjMIPn1NvEhFJPMOZLmFBpUeUHbQ8WRE8cp
EzdIpjoLRtCO77X/WZavyT5r+QZS+wTnUuFyx5o7/DbnOjSS8H4MUwCMMO+JlP5sQR8NG85Uhgs0
2UFoiscU7/itKbOjuO32zG/eefM5hwzj8DWHMmw3JYYXlu5mOohF1W7KACKR0cG+xNV9AH3Nxwy/
YSri/8olsxVQVFlLACvLHRxn2lEBaUbhZVDhND2UjWbWdYC1WAYNiPb77PWJmkF3eyoThNHCuvho
1wQmAX0Xh11bbMecHyIFaljpgscgwr/edrpuPkDGSZtw/nMAG2rpYSN4PSjKg2r7+yVVaz7/yyzW
JSoSMFCog2NFzMHEHx8auVtli1CCzn41hIiBfTt2HIiBAk5Apj26C60h13O1duxhWVK4bYUptR/M
yFkhj+ggUtYnprTYaan3nKy13v2+wN245mg7uG4YfYtPpV9M/JKPk8tr6Qm6W6LTh2NKO643+9Y0
RgZW6DBPcA/1kmULW1lOuxteFqPSxmAkHTD0ZT0WTdH8wqSUJI9cgoMys++97FvX3UTGN0sGsZDf
Itim549rLULXKvWj+r9K9oVJGKwpAqsQ1SmxgguRASBPcwTEFd6bxQkWkwamqrtoO1c/1J5//zfh
EeQx/z/FVXvcgSsA7ffKRyb0/aO9rw/nkgWNtJ34hEGdCmMiR5sstGxfP1VpkFQftgkEPmhWgQX9
9i6/sIICnYarxZVFEH4Xn6rep3T0cGY4sX1dWxKKMdbjtfUloDC9YcAKQX0wXGGfrlgOiu+YWQEh
tG9T4W/yi5lCX6SBjyvlEOSccLwacYVQcsF4XZVnGQX8hqaA6wd4KsitBDjZLyTDwdxXUIlrBD2Y
uM4BmbvxEX2wZa2sVCODcxSvUYKEYhFRa5zJ5kdBlfwyPMMfM3ocMXsm5J77rGvr4OV98HCo+u4W
sVI/FPqGp1WboWVeV278HZ6EDzNZN811m3aluW9t+iHaalsehasqtC3AG6Uiap6qtORzK0GD8erL
TiyxFU24jOvceuLs2ud9mh6WXUSKgWrwr0KAtl3iO3bHHiqUzJCfzVzrk8XGr8nABlM2Hu0kuv8Z
GLsiEEaYXzui29NCwsSDMcU83W6G7gfqgnZF3SeD1HSAYbW6FSejalpJAiKwTeEtV46maWmh8Ert
lU7IXQ3NA7nFi5SBokdocPButTQsz19kjxuMojXpVyyQE026PbkNLI/IEQvgq+onYHf8i8SGc6ZQ
EFAFfPuFscf1dzLODpTFbjhpM1wHkurQNAJGGmZjs+6j2RZmAhlvqotLp0sC6ofeVZ5SiqGdv25T
qF4xDEPR8RAfG3i4fOsPnh1OS+aa1f9HUnj/tAIxjLeJY+7+n/KJoFltsiKU0+NEf6mbUS+71Uw7
0FHGjkkHo1gu+OJxJ9izpfVpFrAIJVk3JTN899ZKmAaIXqLvPkEYxe4umwFG9Lm3lFMY6r6IClhu
8dJR6mszk9p9Pi4TdoPfNvgm6DhCP2qouKKi7B6Pjft3xwE8FrBJxoLm59vWWiCoc5M19jL/uADG
u3WzLtZKVbR/RK+hLXGgQSBeMh7vaQXAJ9uWI1Pgp9/cMqcy2G5gqD3JqES0wzpndaUQICt+K1D/
WxIqX5AFbcUj9vfL3jsZsfxn372K89qyyBW9VElDCypMR5b8pHRlYdQLaga9Vk6ZVF98TmIZvAeE
ZL+jU0+YZhTw3JeGmR1ay7bSftl87c/Uz2jOoMdehcHjBb6hHseD4A3w+QDHIr+CP3r9cJNmeYFK
vvAOOQxioTmsfecJ4fBZYSGuDzyzCjU5YVCwnedTiE/UgwcB+aW3ko3BJ3rQkhtPKH0RoP1T5zJU
fwvXSU4SMahRFvMmuU2GzpPteqOT+g1rvpyxaBtVu2LVtIsc6K/QSbDWd5NJeaZKUj5skCTyIm8h
qPZdwqji3if6lk1vToZaOj8KqEYnguEF4Z6CXlPwUArNCLAePUkTp4hUwVISnfrKsNCRueyUyWP3
pP+3okBnLvbEaYCjNBk6q+IUQNmK5g9/zvn9BABMdmCEOwQNnek/mev/ILNpvwf0iM0gatXAS57+
uL4ZO8q4gbdt2fNRboAd03agCqUVv2U1eP++rSyGqFck0nauUzHMR7ywM4rGRBc/RspD9loJ2CgM
ot4bq6DMIHg18fWnTKcbxXLtQELbsbsiuhIdUxIVg9d1N4lT816zXdmr06RjzSqM04ss24qapcGp
EQJRu5tiNHmg9Nb28yg663CiJB3h3avKW+MSFL3Bnqpm/B1ycc/YXmIfJ3WuG6+cI2q1aURWQvJT
kHQ26RCBgeeiaysNENzmcynCnXuE5tCXMl+hGNOn/IsFTEIHjslZVKJrfErNcGjlyNgWkxaplPFV
yUkIHc/0xNtnJwwkzEYKe9DNWSstclT03jbsYQ92tvQN1ghjwjBArQGuJYJcD3dtEvCMIhVy2Lap
i/BXc+qVPFtXYXqlc4hkJudcy6ob5wQR8dzty4HKIc4Xs/Jjdza8RRer5FaVvGaV1wNLJ0G/CFIf
rOiTYwbACpwttR+/2VDNcjVG5UZDtNII0JR3EZwWMuPlCNTnUm8If8kIeUWhxrYr6dAEDo8CSHSg
rZeyz7js4OIgj+Ty8DAobRk8/G7vkyVbdEhNDmSneIV43FChVCYsyRNZzmQmsu1U+vmaayri9SHp
3Ib4RYBp1HWwSJVA1SDL4bcxD8Go7BT5FPIEDxbwrPBE+TaRcPMWQgjxtIPbFm3WNQPZ6vPQwf56
gv+4NB0M/S1ixOb9FcgU+qeOPZHqvYrynTLOUBh3MgfNa1ROW6I6h7CxmlWCUITDtOKUgToPeXHZ
3lWMRWBs/tCZYocJiVHMK1uoHFkiSE/9UgHXJ9ffgLawnAEe7Y/RaCu6dm4R7DRRCNtb+G2rrwdS
du7dsx4p4yr2W/UPCmiNlDguPyRrWgPEHxKdFK2SRINc/u1WEbjmRhyDf9o9ExkZ6lgPooRZvvVM
TaXXQyDY5Y+4o4hmq6y+71b5Exq16vmHXHKjfkRlEfVrABCN6di7VJi1hmnkUdPIeSKdRfNu4IQW
Mv0G30ZDB0z9z+1/JzYdd+xc0k2A0Koo5BuHeArf9AZMHM3XUIGGbUOJ+JwPHCrN3LaLP+TRl5P9
fG5KqDfpe2mN+6JliqV0IbMfAVV5so2FMjXYlwTQuDFS3xkybv75InUYfztR/ObHzBekoMKBfuop
Ly+HWfZwsKzVS9AA8e9ly/hpnR6yt7uCUjtI+S7B7tcXFjklcvCglL7u3Pp7P17JEYnH8fZqXQVH
9Ws/pOZ3XYxpUJALAK4LU3bfXrOiKRpjfGNi/69j3CBE7xKS4rjcYU2Y67u8zsAJj2aaenuBVD0x
iWfcrOKy2excothoyvahl/4dC6OQ0z9elAB8eLWAlEbUXjeWuY22Pt8DwWMpk1tEzT4LdKNgjeBR
abbRZ3Y/KVqAgIoX6N1fPJU6rVBX8Z1g+8xXfx6+DcyVRjwIuX2WDq1EkRm3VsXIJCBw/LV4WlTQ
54eUGIOmHGmsA/iyi6R+kSBKjS7w9ryQn6ObYXJpeJzK9BuHV/SDBP9b+hprxOf1lSFZLANTi3pa
VU/+jOD490P/iqedwoFUYKU1TPmKlgBU2xaodZg16ULZGBbI6uEspAK2TRxIAWNCWJCY82UnNnOD
BaCTDDet8BgU6o58vTbsRm8Q+FxTjJGGET3yFV+eYbnpa2mJ8zHlYdCOpGga43zF9X5hcs6wQfau
Gl5kvoSeXS2G+9ygfIVYRWIpXaV+s3+BU5XMRLepUfrHldsU4EL7xMQqw0e3fJwpVmwgiudyZ6yH
u4OS2ykWBM1ZG83yQ8B5rF3sFPrgfebtKTrPJ1FhcMcfqNDvACpHmWKRhj0q9P8f9uKjX0CoBdLV
YgyBcREq4kFEpzPizllHctgAOQRUUyv2dzxbaW+qrlQbpQnZuFhc1A85ObMGCYnFknb1GjroEJFH
de0R7Udl6c8NEFh4mJnPsvUKP2ejZSZvY7Rm5U9O0Rk171K1D5YIP/Nyd4Mt2lipBofDyWRkhGy/
RwMTvW0IOELYCOxOqkdsJoLtjGAXN616URZ0ALJoBWQPyKfRKmchGGCf56+OyKzo2sIg8pdE+mB2
NnKH08sCsWfapqXQfIfDz6e29JJ/wPJT5gbYpVOOE6yyna2Hlv/IAkDcDkGLmO/konOvf/rxv43X
Z+JDKAoGU3M07JtiuYGon9RVipxWYFSaHRDiiZVppN26myiDi901Fard2P+tVek4QY/THjeuSa/7
SU2giBsGyMBAi7CS/vgTU5MJ1nx4jb6sbgBbsXuoXxOcvqNQYe40JhfJnJRf+NMXpLARq/1i5Nzx
3JSt6EjM3hnR3HUh+tJjHtwNwgMMzNMiJuLxo2iwni8ETI/Rc7mq5Iy28D9Ll/rtmjoLMsR7OsNV
AyshYiq+PnVSEKqDWTmkx4HPw/eBTrKVK+3k0O6q6+R2/XpcrJEBSeSRQWlfBFkz1LYMPrLJJ7DR
H6MLcr0DPwV7apaF9gP+9SQpXeYgHzx7iqfYIEmdRd1kNuNEY3QXS+hzo03CAwDyXDQOyXdYs1H4
u8WmfzbMvfJgUocJPCwsxHBAYyHyHUqPsAUZsAtheR1jtdjhvR2LTb7y5Zh2mjjNJJqTCmqfTddl
R6P6s+ind9F/1D8FBqUXtveHvLrbF+8Ksms2CAoxKoPSG0GBMdlZfK1gD1VrJRvUP7YgUzG1vZ53
PoD6+aM5dk6o71yrp/JUP8jN3atuRbgfmPaAjltUTEKckggWm3N2EXBuayBeQpfwnqgK34vMVtiU
l1KShD2T7BfDnXP8YHncZYbyunkf5H6S7F6rg8RmDcpxLOJXDMzCyC4FVebi4nRGu17lMyu8S6/3
H4+n0Ca1PIsnrJPzMzobDj/hw3js17qXo/6GvPDwsJ+1DCjV63i6gWiCPqs7Mb0seu3CN+1uCHWM
w0FqS+FGG8rUEeUVD7JEGkOunLpe5lQbRSG2hRA+euuyE324RV/ntc2hDm0fsnK4eNN0CzwHxUGi
A7OswEEVbMQGQYIIvRMfkOwOycpxignbHA7aOCXjYjVg7L9Iym4H83lGUO3RnP917G2MPWhPBlsY
16i3NEDZjzg8baso1ZmJ5IZ+GplL8Lcpf8Bjpv7ztFEmq1ve01NQNOb7qriX7tjtyhOmOAJ+u4p7
nlnZAPS3XGUBiYGvcwlulURrIV9szBkdEAHAn8cOOs0YeO6kIE3r8ZfWHrokdMlsNEVjYJbNzx2X
ijZ2U7gql7eHmrWpLL0PBPC5mDc3Qm3+M4dZZ/2HBk6A4fbdS2Y4MT+sQxNTNLAW7eR1HKgVTi7D
Zzfpir/jsirwo5OomCQomCoZypBHklkY2u6c4KMPbwjeUP4cF00fcpMi/BJ5UjqhL1KYAWKLV5GM
Iu/T8edNAJ/B9F+sLuopBI4S2zdzae7nM7co8UTsj2jlGHsvo/mTgFRmPDXYvwrNP9jZQAei+d7F
2hq0UiMiur/09d9GhHMQbPL4Mtpdlkhr5XIJwL6UnttwaBRiundEJrajAn12SMygHHJbfSikEX7D
5x7Ksi1A/xt2ZQDifSaSbSGd7sYw7/c9LepySJrFvciZEg9lR/J+UN9866IvHZ2BNZNeK+iMwdUD
mqkW/1NTvDBBJ1RKrGaLXmWl95kFl81COyPUBHLUK/KFk03owHfL4ivF7NDJuWJ37GsSZN1uNv22
EuJisFiN4Fif7vaVSJL1QM2wjq9OKqltRr+onHiymJMMttSKL4vvvdnrpIu/3nQSDF9lCOVfUYhk
BXp/iOHWa7gC3DFWbkehZEPeqoUhFULkIMCRfNMnQ1qDSe79mPFqAsGMmExgBkyIHcWJoo7oyKrt
67+x+3YhVxOCx6kZfrQz2pCm9VvDLGDOpZcyuU+mH5xXaPa3zDZLa9mZR4wepModw2FFgrrs/uC5
BJQLdmV5D7+eg6myXTUMueoHn8H9YLv8a5lIogNYurPtNdWNEiarioCs5I0YYri7IpeEB9Vt6MLh
mCzKiyUwhKZzyysMJ9Z1ea9ALjSsLfHRMdH26ySbi73G32dcOh3Dm+f1i67ENBrcXphYfOZPtAxk
tlPmj1GDL4E8FPfu4K3QuPurVR51e2AOugOaShKROjj4IHn6ewYZKJaX9lDGyurxaXGB2luvYZbP
bQu9fYwiWoEw6zzGjWNNZxGj2T0il+6T6e3S0U9oJ8EtNpgqgKA2IXIWT1U+5G7eB55vmludTcvF
gT3esUiWm/sVjsWONhmNp/zPSGcWPLYdFbDu87lYmALCIb3jkwFVNEuOXdFpZWfdW3QORrfbxpIR
HR/3U6ei68ai4IWodrwWhZvDr62qBBF3QA+u0UN5igsgK6h6og+nCaULGk2Qa0DRleRTyDIc18mn
eyu5ricqb1epp5yzaKZ6uPQAhOBJLbGFKq+2TkGftDdE378tppa1Lc0o1bZUuQKiSBt+gdXRYxiZ
8cZRnxuVAbFdKhrHYD45Mpvqp3renMdSQ13WLCupopazE7NwqnN0d6O/KWHAnJTaKn4fN82hSoJZ
uVVZ33oPDQ1bHilhTKFk8mW4Il7eQCyLEV7ROtDpIQWaiPIEpd1Ixbc8O20hq3R+kOXaF3bKqICx
lWoR9t0R203W0i0A3LoAYIxlUjgcDxGb8UWyZRcjG30GV77eZE9cWIibdueIdZLvWA4ibnPkJ9Co
hhkG0wJ/bTlqooZ4gIwAPVMJ7ZyM2DaFu/PHlFiJakIchlEn79WolXB7Rvd2TLLWk6t5S1ZmG3A6
JffvTVFRayhZ+IDzQt3LihTfaJX8WnG7dWbyoZcidCnnD0oveRPTI6K7ZuK4YG6ks+z2QvWmFiLE
MPl3a4TpyQgMDnfz6AlhkhrfgWRRavsnP/LYyUvVQ34DYi5k+KfXPBC67L2jV+h4MlxquHHXgZVx
7Yy3CsxizUGTLhqlh9zTG0hk47CgaHdZRRde10xp065AeYzDspm18mT4Zq3B/2Wd8+G3QmVlqLGC
H2xSyKUDhSIIqQDcobH2ZiLZJZx1cF23SFW23hVooITj/bzTfDe3/JgblgvYzByKVasL7YCgPKvH
evwuu5oUBAzZWHMPN6eErsAIuqPBTuoQ7loOKH0wQ8qQz+hywDfFpRgbmyieP7F9GocnuPp56Nic
ajK6eJp8EsYm6l0rXnmA/yNeHDMGRTO/7ofuit//eZbaToXQI+MYtZ+8VrE2lsKhndC6jbjKpBfW
Gxabr4ZV6NkAjpkVESXC31vtckzk0Ckr0NwZvtNJAUp0pFK5OCJr/Kkf1tFVSe4x+d1+gDGi/2Hi
agevyz/WTpM9v2gddDhxJvAdO7nbtZW7zYIG9kVf4jXB816g1yVOyEiayQpEUS09OL3nqlfegknt
BQ2kzhb2XeYze7MdurByzA2AHDYq1AXYw1ZIzbf51qR8w0VVvLKVjb3Q5ENk24sAKjhK4DXYPurX
wEZzUOJw4CvGk0VZdOy9ycbQf23DquTeDS2I3E4d7i/MVDYri9glGNLFX8XVYDoNgbhiwZML6uiS
aG/4jTN/jiyqXqX2+0LL5EB5E4JTb91d24uIbcDqSilJ1azlYlfED00ck6WzxfCB0tP/UzxgC8gf
mqy/GNu2o4/EjgpAKZ32fdJw8A2Ey+kR1LOvcRTVi+9FJe7tVf8AoRv9Kh8vtEVKVikLDRDTtji2
4qHnH5VMEl6Y0ko6BNFTztSnIBbev5/RjQQ3P07HpRqEK8Z6TZXLd/IkMVEV1zVHMYlvhwU3BOnm
vOfRS3OZmoRQGWKA0KHWsuAoduof+IHcw53MG5bnjhfCsUpBj09u2y6K6CyHUx2Clb9My+SpCNyt
gYQp3khJPj1ITlZCDvB/N7Ph4/vjxUX7mKSqpv5c71UhgT+wMDy2q/T5u1jzGQS5OFJyas3+hYsu
AYUDzoiqTajhs/XxYr7Q6O9S/WprByLgO//+oMOHqgxSiK+OhTGaxes5FubsmADTTSwi07xKhmkh
9Me24uzKg8mgMsYDQinHmfUJihsrhR1nlX0ibsEk0LGMiXYbZQzB2GpCuT3wyfo6OaJ+Sf0Uhrci
ocuH/ZCgcQ4y1gF14GcP5kR3yaCr5Bgybcv/9/Y8NkNcVEqFjqiL011Tvw7je546XG/opdDoQkYu
PJiFLDdSh5793L0qF4j8g38JrkrgSR3C2fdS/jlK9+vifDI5NwUbwRnijYuvIfcm2wl0wugXM0di
1qsITvEfFjJYflz/UjI4n3RpByEoGUBERXS9b7l3c5ZojzjG59hcuPj+NT+xtIKzxIO4C0GL3d0q
aMkbfP/bIu8xjR7QvSVLqIF/Qho8uYYM1Dvwafe6AK9Mk6N974dxZI3lv9vCDmRMaA3ygZXTAcqd
qATmn4LPUo2ioEvetJF9QtNbxgLh0vjk1KzV7elDPDFcEtKdLbj0Udv/GrQyuTjSK6gdbAsBSSO7
rX4O870cmeNujP0+r69M/0gXqDBBOttuwiK4sw0kU8mcS6ar/mtshXcPdRvurTPvAyhOynVYwcEh
JWCfHqwjs4QpDooyPtngrj87MSgoC4ctj748gtS9qkcQBM8nMyrWlZf19YCvfoMaDjyhKkQcZLEy
9c2vZPZ8RykxygVAePF3JJNL7uCA9mdUW1yuVI99+tbQurdDevfMe2zQHF5xjzK6jzH6FDSXFAGh
G6hFLpsUiXgQVbkTSnq3+gmvxkepYcqzhrkGYAzROBa7k4WcK7GexXQEuoY6RHcPOEbwr9DiDE+w
eA0hyjx3CB3VITOua0Ra25gI//MLJ17gU6rs38qJvVxud1i/qGP8DmCuvuTMKnamp8rvVwM3jCio
9EtAFuBpr+fVKadVlpFX6jQXdye0TnZ1CnoLaZpXgvEluI6kF3SxHUR62ubUuzINMWxZ2o2s75wK
igQrq104PLSn+aEoEk4K0nilCJsTfxUe+fKSUZPAO2Hg5Xv338JpWiexmO24ZdMD38lsXxjIhZkE
wVY7eDKSq5OpLruV0er8AdusRCgiYHhTI8ZWIZlPpK6WpEK8PNPrlb0mFIpdHefQJcED84f2mfRz
moHjRGDWVrKscGovXRaePommY8GKNMak0qatCStt9H39Pw6FoNE/N2pA35MCebvy3E8MsanqAuNv
rFJTh+3z1vY0q8651FdIqMFN6OY8ALMbBL+f13pU9+6qNLziRU+NJgbKIbU5yf0JAC5+l0dMH9RA
3ZF7dXUn/iBF8iKpvtNKKZjVWr4R77GCXKFr3ey9ZDFwOoC2SZg8fC7HtcaVM7ZRxhDsfUHjm1D0
2+85dumrqh3b10DuwQmtvhW8nxfihx/tnFExcuuT8+swvfYR0iDcK38N4qyprlJ803u6GYBfQI5R
OE8b+u9nI+X6TQQ5kaBNXfReBHpW/Y4cs8/oxkPorypbpuppllJNQWFJTIGd6lUDm8AusqJj0wLF
PHDbScsNRIutStS3wqCTsJUJgIppDvprs+rFRNyNjJrfuX/wkR9teX7tzzlj4YIL5VvYZ7Ugy8d2
1EMFcmO68MSmIRO9eIh4LGm7cIFjFdnfRU9VnKqeOLnMm1Gf3H553fM8aY6hkyCU1etelOwNdI5f
ILMX7Gbq1bwIH3OpBpYlENUhZQY45qw3+z18bjSHAT1Y3OzEXpYMaAaLu6nRM/7GH0GOnk+eZ7MA
XsIQgZLeygSC9gnJNP4gRERzzTljhj+E0xocChYHACV7aoYGORYd3jLQGdMQlz2ZxwXt3+v9zmAE
rK8yNduMW/R/Gq2ZmyuLNyrBrTf564ZlqVoGL8P9kmPBvdMrTF9l8spfOoZTFleomd0TIsE7R6/z
nUTKWilRluEIyhnlGA1pMWACaFmhJHvfthfYuRm2S07QQY5t3zUWK2bCKAgfOxMf84uUEcH6lAB/
6AsLUaqD9UyKSIk6XZfSsAdhQeh7V9adWHdHzKNUKCxCCxfm8a3EtT9ehzvSRa4zNMIvBlxW+3Ln
80MWsN2o6uMWKuSrrgQ/pOXBGtIcpMZoUhhdRW6Uv8IzkvKSlrxiLKDWbDYRTZL+YdvlJ1dgHWJm
EMH7DIL/NRnB7U6Nwgtbl87ushD9TAwWRlvZGL7glicuUxAWapV/AQWxhyuaodu5Uaki9VV15ZIq
SEeZsMVVvqoshZjNxHuNrcHPJsVwBw0sLnPBmQQ8OZwrxUf/NZ13Ihpj0RYUly6s/N7GjkrYxP5D
AtRjD4q9KYBZsnoMUB6ic8jZ6dgj7krpee4ELKUpKEKpKDHqWFKqHXVu8Uw4Ik41ZyoqkcfPYjZV
WuxUrVWaNJwtZH4m2DaTbBH4N4Drja9u4MgG+T3xltjhHzHjSGNaiazm43OWL9rHJxhbwjL/trxa
m3luiDX5L/8wgsLaged5HyUQjydMlkTBsBj9z8xlClmS1t5Rr5X5nHUV1BX2TIgp0seJBZqRd8N3
QZEtzRQVxYHOqVa+b4mYevgPo2ju22x+diajxr5G2hO1OjILh2UQeFOVHRNlKWICFAG4z1cuanb3
yCTv3tFmiBQrJ9tD31cABHsYeZE+jIKr3pxTPGoa+PogTLBlYCRGyhY6hMxlIRycHdaKGbDNMXCn
/Ibq5LLhw56FhizhfEz7lOck51gmq2Rt1S2q0UIYyqVAfLVCUZx5qIrkJOmXXEJVXhP8tnc8djFg
/4JycXe0vBuTw+F73Finij6bz5oIf4uwF67fVC4FuZKdYC6XJIvcr/trBo9Rt7W8x+F6XmNEYc4O
LHyw+Xi9mQ/l0QreVczVk0hcrqLmydBLK/uJaCB2VkywFb5F0odgj4VAsEV8Vh04iH1hNjYAxH36
tTlbaYug+LY5bfTkZBXf+J7d5b6uDkwcjAxDqhHmQaMru6+B8yMfaTdQCLytCQYaW+QUygzafpyn
ncyH/r0uZ0Djl3irrh86tim99vuY0Cy6IvdcG60Yv4udQrQ8zekztD722gvR17c8V9gs+3dx+n4z
vFIywKZEkldpJg5hWYJbtVwesLdkD+dB/cCUGb6AgypkWckMUmsvd32a/uRsZE+/zpCFI/YEskQO
7qyafzxvEpVpg7JCYumKN7lBvsXl5LCKyKcMAm66eBgyZ4QNv9pf9o2fLI4bgPxFbq44HZTQpP9n
QObaMgLLLTYuAKrHah7UwAV/IRZWSWETbuY4rej5u5m0XIlXcjU1XD99MBJJEkrkISMcuXw298Xb
LfPpYPhMAjxijy4M+wB7X1UAfii6Be4lesj+AK8mVWrx9QXokk2/t9+W7M0Tj4w09gljG2uNyq6l
tbGpW2n/+Ro7ngEXTrjolGRaZfUcP+UIS76iN3cP+naPQPd0ZsRYFfd5j7nSyrweHyfMKHQAVv56
fxt7TeIwWPjUX73K1a0AhwyLK7q8rngq/VrZ4o42iw68UlzHBEIQtVbeaJphNodYzNk3Vae5b9EL
QiOU/DBZ9pQIwvznUJAw3g/VbjnI2pYVFUetO159F7dxNUY3PVCnnwccUEIZcimN862w8KPUxB3b
aoFX225waj9Mxl893B45DXlRf3XpJb9ksS2AO5RWOjzih79wXWMcHNGmFqXnk0YUjkHvNGuT4x2G
RBi+7H754GvLayndkKGn5yGT4BInkb3HU+9DkH0bWszUJjSfirpYku0RUdK7Hx0NpYt2Ud9U0e38
GWK3WOaYyLBk4my+i43UUfxuUjkLkaOxKt5wmcZreAduBCI8qtGyxamxPdK2wMCtE4/3loeRmuYU
hOy2tqO3N5yPdOdQMsZbwaS2HbtLZs6VtrfO13Dyook+PbIMWhZvWlPdgkyJCHcNI1uBrXfMmidl
D1Bzmye9Mv+dIP1zl/tJF0Re9qZULTbeSJYfmJtMkUUMVrcBRnUh6wV4815cjFfKD6Yy5Uo3F14D
pOhcxm+bBGLVNM4FMmQqqpoi69MC8evHMCwL2PkuYJikvNTnpqSUeOKrsXXoXXsFhWK7p4Wf/7wr
iGgoy2mM9nK1rjanO2HNjvOLuikm93j/IlkxvFVelipoz8oq+bL66I2tWmWj42Dt5iKg+QUf/lmy
e4REl0NM/oP+Dtn7RKRosZd6rDOQD+5E5tNQq3yPhStl/+X3RdzMn4AnBw8dVwgFGk02Nyh46sNY
V4AqHaTiUpk1ScnBZ6aY4w1uUJymz8GvNrhaQgsrqfwBq2gt8eG3xZ4pgWuW/WMho5pioUoZTnsE
nDP9mxmJne2lLZcZ9P6JnMg/5K0w0BQl9WTI+LU9KA1kziCiKjYxdFZIGw9kUPQPFP0iBgvR1YrT
5y/zwQPJnMHqvvjMaWqTzC42T1GjSGF0kfPrDS6/fYQjgd1lYWCe2hm/rPpubojCQI39h3kUM9RG
A/64pjwvu4AlmBYdxj8rpkz9Vl17aj3hLZ1WgaDjfoGWFI+c3o/1mtxiNO2KbJsIZKGoR232xRPz
Or/QZ9WZONHKWI+L8fZOJk3FgfqPiMTgSx/dpgWnqtm+3KdJ5igUS22DJd3k1RS1ixjE569eZTcM
RHREkjwisMGW8U/mWv0L93mZ3DyH4nAxi+QU3DJNBfcw+dvS6BBwmxpZAN2XxbZq/74Ex2OR8KA3
3y4kwxit40NES/vgGsbWWDXCcz+p1HxfT58LQRyck0HpVETnNQPjjgeXPIK7Y96IYZfXKihBBeit
3PNXwHZ1YuI7zJhjsQs+hNL/f5/tDsAq8gpv52AuxxzCN/BCnSqY43HCQnirgGroSrXocks2wyOy
/5+7DOBw/Z6o7BRngcmvciAjELsaptL548Jt0XIPczeqYOfQMIVo95cAYazfdHJzp8R/iqGJO6sj
7zmGpHoQMT5bTBXwWPpD1tk7tDeQEXg0tl9rN9LuSAIf9UmMFNZjV1MC/uNGfT3HHencSUaXeqHb
qSnime19h4cg/Kl5iqPDStnPyyCSMXDfpxNo+5UaZDbr5oUkW8CfsHd/jvq4obzdPzF2agxoMUgy
o0h6MN/wO64lHAkLV9PAMuj9+H4ISwAMPoFpDq6R0mzEYoc6Lnyg2THwyAE5pFa21Vz+BZnGNhEf
vkerFtCwCRtntTjdhQgGFZV26calKklHBjX5DaRAyp27HVu1/DJos5i8ZLG/JquKe4CaM45+ElXf
jWsBEdCJMHDGvdhGIbz5ymbjS97TDGefibW46lvrTU7mRF2X7qJ0CjK8dTAXM8itaQ2ni7XMBP0m
9pqVJDY3OZpzB/hPidz51ERQVCNhsJxX9XA+81x8cPeQkPAfiV1sqUmd0ZR1T528EgJ4GwktgjhP
ZTg48FhO4PAs7MbSTjSaOTQo5rQaCn/WMtDdvzw5YeT92HHHmVVIycgSJbFIcMK3Jxp6EfQLItab
Oc3bap2AfOfvMbovkiIj9nHjtM+K93vIYwgfn9J2p6nzNDu2DLitcWpcDxDIjfumMb57td7ZRhxW
lyPTCMI3dS7Ydclo1F0APrq+DU+LnwgMES1618/LzA7YYPLu+i9A9d0XNEBI+B/GCXCNU5ZNvnrh
LyKvXGEI+GMvGeTvBK8jqZeYwPFCPvFLYkP5csr+Ig8ee3Ne7mRBFE7C7nxLY87R0jXWIS5oj1RM
gXuSl8UBoKAhvW61aMx4w5lve7T8hplaFKCRXBsccc0S01m3HVkNIlIX04NyjHbMAuiNlrOZrK2W
Csz/DN+hOwzrPzhyNbSwXU1nGpPiDqb0yiu7eDGMO8Xlmzuw0mQ3eNtFXF5084TgysmOXlRa7u4J
e04J+Y8Zrb0+C52zAk9B3s76eXqoQSbvG1O8Q4A8l3JvpThKgdrkCSep7FspIbuTHGo0c9ryYSJx
RAbWOngJLCrD6MOtw26VQNalVG7kVMrZF0Pyiq4Dy8gm1mGxm3kgbtefimnTyDCSc/+/URvBISQY
cbFXJi52/0T53jtdwsB7Bz76KFkoBTRH7TvQ6bHxl/Aey3GvrZW6upBcFy64V3ucH+R4Sfq7w4dL
BvU1xDu2VBFR7hnYGR3+Gg0p4TZGpngq59vGvCh+JoUHC5P64w0dkD93ZEkul42QYz2j7LG4TETK
RwkoZuzI0Xeum+Xhf31vkrqiH9bVxFAtucb5xMbigCbNjRHeZ75M/sMIklMEbB6/Sf25rjXRyzMv
dzkv8EXd0HOYjl92oo3eu1WVnxzqVnlN+y7P39r+fRE5FswB6PlaqNduCj7UAFg1bygjsxo9xced
hI0Mt68gqmriU++mCCZSGLTvLJTiFhu0ifxIf597TEzr5AQdQQTKN9MqkB80KfCPplCsnfcpbF7h
5Mgjg5pUAcC/FSiwbIk+uWhbpahBMjpt0dDFfYlJklkRrcSdRhBHm9xIYbLlbgo7IX0CmzibxFzX
Kh5u4m94/lCeal7lmgY+9+eATclvRY2W5Hii6/sWLcebXvjyE90/+Ei0Aly3hHS2yyO4NY8IQtum
aRf4f0AKor/+HZwDojjTe1jsL2GvUZISTSBp2Nn05xlIUm6nsDLXRMj8Dl4l0ot7GdxVtuZ0hD4Z
7yh+A8THGXG899FmsZz8v2dJo46moxE0SBY+q8VCDdQNsjOIAoE/dItUmO7qWSZIdNFxZq++aEZv
A8/GT19iAC6l66ff2nsLvZk/3B+4bpTOympxhBrIdnhFAPP6XNdPZTqFsMTm0dnjseNuc2Mxsmaf
A6IOPbk6eiq2vu3oW0Arr8hl7iP3PC/OcATknsXhGzbiXNi/+FDkbPzAUI79SB9ULrZcQj+z2uiq
LQfODg9Tzd6zeQzJrIrLq75GFCVpeSKnn5PPX8tY86NNp7ZPjcLdXzz1ReYEK/t7nEsIKP03QwBb
2Zpy69whtvIFI290VZKjVUTnz5WSUhcP3XhQnq4rU/luo14yXZ6VKtBwov//9GxQ9qXKi9JAhcAK
HtM6wv+CgCVqJLuVLTLN1Y/JFYWMJ7ikpC2l2wmrTtUxxR61Mt1eQ8sqstTPjKkX2Tbv6DFi6oCa
FE22PgkpVPXyCzgaKSr6ulhaWWFcBDVd8NR2u1h7SYU17y5OKqUBiqPjIqqy/bCG1eTyG+J8KAuU
9L74uQViJIKv2pMUon7WCdQPZj5UQMcJnOnxETFDHLBm+HxfLSqlnZwTzlux+w+gn+eKwZFAeGxz
eHiRADD+4TxHKpsm6BjaJgfRKvFYQZQWPUeljUTr6TdOW7ljsEP5MaABEBH5ES4wffqhqdmwEup3
CF+lZFjwetv4MDkpC8t/8ERwj2eZ4soGUpEGzNeGV1zU6229pT+qZWJAcU7F0Y8BWPgo9FVzFeBs
RPBkP34PiI5XfU/YDswqy1qCKHTpX5QsOJwRajnkYVSiBtHB6VtUTbgeYIWFpkXKR5Ylyjaw8o7v
xqAgYJCiGZ1doYznJ1/CZuTZUnmMCuZeesRrMu4Zpapftoz1XYGJc7PDnHVxWUseWkZn8QGuE/io
dXx4pcpqKxLRTzBZ9kRtrUkJYjuvhmcWnjmBuPDq6i0v3TlluJ9ITgCqqiZ4NQSbyTM8ocFfIspt
M3OM0XHgUKCjFvCZTArvCEoxs6kuqOXCKHobWvllICM05HBm7JxN9tiP/KctTuvL53UL4yNDOgpL
WYVlnc4ncbi1jV6J5y4kIr+FjfkZYWYNWi547+lqRj1DMUuxXf5ZQTQbOB+scJ0tXBrC+J/4Hgdc
jYP3xZs/rwjHix3B0FUbsxzqsXz5q7qxNNR6T59lynz4IKxubP6CTZ5DnZWnvGl1hhil71ZIF6P+
tO5V/75Scc6v0owwlG4KwwNQKvMyABsuFxZ8bqf6Go6ogFK7xrZTSu11e+eEzs7kTc5/wv7O4vLv
TsqPr5bFi54m9jEqdMWWkGnz1L9klJluw9P9PJ3gVrH1X0HoABNCn0b8RJS82xg64IOcGvPOLJKq
DHmpsHqeKIR6xg5fRGKyijNMVfDXHvDIzWbek2iKBX4T2RCX0UU07GXTkDhalGBp/U1dErbs7pKL
j+e++wx77cHINVNnXVsmWCOB09VvrKbgIWWsHqFNkClDyxZq9/vjaYKkOfvxyGlRHm75pk9YnGA3
xhQEQV57wqicHa+aGn0YeZ9XU77I3b/M7WYppjJP8wm2hX/w/iGygqmTK2xtSUGvxwDeTtkroQ31
SxESIZa8alcpkpVOG2+ih7l71TRIZRfq3WhDDxBtEmMaIEwxGhyA3gJKQyMGq13K+VP2ARkRbN2T
WQ8fe3th8p87cSRHx+GfaXJ4KfqYvS7hh3XKVwqR4XzpIhU5MUFqNu7CsGrbitxJt6t5Lu/fyI+F
rRN36LpI9meqBzOqR1N+IZZbHa8X5VVtgBa3SC5zSZ9WEYloxhdGgH8+t4IW+jwoFRxSRtEOhV1Z
5xztAwbgfNxMOmsycSTmb/hVRNU6+DYamRgBOgWsd+Hu/odaWbgLTny31LWZm5RJP2dS52wdzo2d
05ydIoxsv3KL+wzKz69EATKY7PAeZvE2NCJlpSn8jIC3FA74mBhdnhHJN58dVsoQHSyzLudjUdZ0
yuUQqSF9VNLzbkNNEUKyJ/KVZKTQpPtQ8E1dqtWs9UvUyDJyjlGjwuuclpVO1kmWVToA+BbhGeRH
mPuFEqB9HnXpS2uOGo1p+l+vwofmUHE0oxy4PFlYPBLb+Fg3n4nxkE+QWcQG+6DOMSLM0g4/opBC
WPEQxtEwPq511j7gHhTd60iNrBJ74v9svrVTh51k04+zl7O+FiOFzV5D0rhUynZe0mdlgzZA+/1m
WCRZDaGg+F+vv/SWdqqV0ZbLvSejsK/3O5cHl4O9qGtCtdW+XRxw0XF/7YnxmiqwWxK11ELJ6UP5
PMhHgM1LZUP472lbJz7Z6R7q2mBBz6gwdXgzImHpmZwO+GJw5uOn7SDHNZu/R36oeG3vuorcoi5f
OJ7Q2ovQPAcibbRQE96SmSJE9cQPOrdnGZ03AWQIxnyW0ul+RTV0602fsFg2sei/70qyX4bZSsbR
FW5oXYd3X1FTsV0IOhl8g7sajA8ZaQrHikhUhVFP41tYl34vY4YgpwKwvPWuBmceqf0aAKcZGmHv
Y29Ep8pc0rsSOsn603NHJdDIkhw00nEcyjk2UjznB8ecRgeoCdsFbWzVQsKQw9mE74E4RUgKqJhX
NkOsxMWGZOjPdfa1v6yd2OuROwtoJRbUjtXXz7PXPh/TBr1sIaH01HqhjKaj76IdQKNrT7QgACF+
U6aEtNKW0h3aRfLWCVjPglh+FRp9HIog7GJHveRae1n6Q+JFQ+1LDWFFXRpqev/0cOrEBJBZYnb7
FEay7IWDOxBoWw+ihTwzPt3IRbV0tQHIfhuCjsW3osdDxoFUhT1nFNm/gspYDWtsF185b79yDokR
0iP3WCe5D5igHkj66qnWkuBveqJ96jkbU7Axr3WPbp3Ce/RkJsomaz4y9JlCwMNIZN0XYBdrlCRH
0HmEwCm73llI9KHL2LIHE8RyY11ATLFg4zoC84yF227kjFP0AyVVr2YFjRb4CBGlIayACiWyfHwe
7FA29TmjBhBl0s1/AfKpfmE0NiyLu91QvoRMlvToffaSgKDgNQinSN2eKhHMNxfSVMIWwopAV25+
a6QiuzcjxU0rSMqJjfgz30Hm7MU3fNEYQlQYWbEsjeWHyBiacmqZ2hX10L2xoV/bV61kzBcaBo/v
7il7aTc+o4gLMuvvzAwiF9zWqvjLwPICVtJhIThfBl7KopcXkVLGWKQbza6TSImOb79N+C8K81cd
XAtMwP61YYse6iZ8RxccfNxgt9O8+yjlawsdb7RCbWTJlIPPCh9vLGPM4YzVHsKPRlHPnnuT+ng6
7S5fGyuL0wqMS2HtC7QlkhgT4wX8+91l7Vuv5e95fFPKi6dqDqffqD3LB4q57nHoq9YN3P0GRXFz
PdXa35CPm+7dcQbPyJX5RsoHgS+QxQ3GNYLfYHjrDwGZ0RVB5kdXGWKCSaHFmxkk41CNnG1xXTpw
YHnEQTSKcuaLkKdQO/JUR5vnhb+6dPrIMlxZ1WwbwW2FapOk4ouKDGRYDwlz7/BUAO+e3/FryVHe
7IG1ZnPneqyw+9zUavcFclIdXo3uyYSE4WEkfDq97NpZ87gdAAIWDpWUmpu/81l7BMGlcoL153YY
NHHTElC8K5/2J9DQAChW9pJywy15+v9JPpszYCr2BDCfzedpRF4q80O8bshlO9TyuatOHKGPgZnh
D74YeFBnXZs59hFS9u8qoxH/FNRGbNZXKx8v9fzA4kYwCeZdXel4+CyegdAHdenlsNtBOoNjsCmx
WBwQqAcZSJdTicxlDmlMkAs+k9LXol0BQ1N8h/Y2NCx7ADzsF25RbUXxCCp6/Q9lmRZoaBhG0DT/
FnqCJMPa6gbPBO1ckJiYWhmwsUiYbWSdgmTs7kLsVImJutr6KwNK+hUy4BnY1S612uyAG4J7gctu
+ujq8pn1zjUR7yQU9vjNVQmO6IKyTkCNPHggVSS8SFUVeGt0TYiJPdXsQIFQRDVbQuSR/VL6T0nE
ceIrF+h6BV11rFL9iwuJld5/6DQYfeVrVU3RuDmY8xsmC5+cVoeguboK844d0zP3f+2uNDLWeFV9
dtyLusNvxxmrJxRrx06KsYEU60jlAtc3sZs2/lyfyZ2R4IGsLwX93ZpQkbrrGZ5Zgs8IsecHtCiL
iV7vGCJ+oriV9WiTvKqrkFKzAyRcWwHYrGLMNUTLg7MZrmCriWsdyRn2Yo6BDGVuIR0TGpMRFTAq
SQEOnCkaaYD6NbBzpxH6mEZYh/0TSUh5SmZ0gfJyF3JV35PWqFgR0dIaQaY1sAx7fpIYSuKdnDYs
WTTR97LVx2neOdNCtBMM6AQRQPbHvl86WSAOTGR94OAVVSQxys4ldGgbx2z2/mawz7zodw2GuUoj
dxxGC4A1pzZBZwl3eQv+YwvlDuf0D/WSyzHjWrJ5rTXjxhGY1P9mcbJPYbm8kfrW8YZ8vbNfI+bN
4QStWW5tRFeGBZNHPxc4ToGaB4D2RwT998E32ZZdaCD6daf3entwd6D2y+Y7b0AAHE+KLUjqfIBG
Yt/Zo52BjZf+2ChqgpEl8k1LZ1RL+P22VHI7Ge7NNV37pxCboRSE4yoaX/Y23/3MLozC/T/VeaO5
d2r+YiBnkgI8yjMteIjvFzJbP6l43g0toGaeoqM3QGeg4YUOfuqyanaiStIv4DjhbV8E7lgEDXZA
OsKmxyO6KPgy9UqM7jdLyXjdTBQS0c97/OFkBWYfH6Xq2Qr7INYM88UQQkSMS14Zvs+eK+yhoDdf
4JHB6AvuBNFj21kQS0BuS9K5zMEYwIY5sbcaEZWR4Q6djmew5YyW6IYB9081WV//11tTq33efNXi
y4sW3LfVU+NAvmkCFhJ9xF7Z1gXH0KVGHTKC19+wGqudcJg/B7nhvezMMYl1EKQbe15MHxaRNzkf
B1+K92lZlQpFsEYNT3TNFBkyMB+g0AWsDzWBz2jbMGtFwac8OK1KBE9X3m8Mhv1p7C1ehb7rCDTT
/1rbeQAKTV6ef7ANiMmDQDuYxIALwTFR1kBCPAiKI3cK0seDNMVcrJHsOiyHHiaI4S95DiANBnLJ
pGk8YrA4BYtGUYyw+1sldEPjBytn8JZHDo4TYqxlndFnvtPFHp1ysUZaQi/9LKbXaZnTDrTM9u5N
KMvzD5kNbZocaXrlhPPHRw61kqPgAUpjG3noaAFBxgMwVTKkSo/3pghRbn99y+Z2m6OqEb3SIL5f
uys/JFgBMJsXQzLaMu2f+rURiML/ooGa7GMGfakJo5LaYqMcCFn1stm9/SUq3aPjHO3Xef0Q0vz3
jAVzJFdfUFyMrxpHHCCDX4alJ3pNolcW45If2lfbw/PsPW1bNLqr3gzTBweYhQAywRm2MCe82dtb
01Nst5PAfHjuXnCB58eqwvjTepf2J9heeSPB8wXv0mobJih8rDOnz9WydG1LfctbUuSkDiCu2ZqZ
XIcY8JzCNi+RQtPQndjYxqOGoqwaAHn0s3lIGfS/HU61JqMdw/Pne54bw2yq0mO/WRfQLJ1WCTMb
9/mQXjFZtOxa1jfzNqzHQanm/1AixXrol3gAiJIxJ2WgYkrVmp9heOVT+wlH95w56B5FEwxQIRGp
yUDs8vIjdjdYUXwsJ54wdBTnQNdgL+EBqrQ7jNgS4787YDW4R/54hzh9up3HHoyjvqcaBFB0n9PR
iO4eoWu1h8IRmbH8nvdh74zNY1AIzVxC2kPXVPotWzyO3Q+jXuGt2xsupuaHcOEn3TSj69lBHrQn
CbBGkjXzEkVRGuyPHhSUQYwKDcDJU5KWuHe2uR1dEDkXQt9fhpRbTMQ98593BvWoi3VqXQD+Suf4
2WvV/xfefR2NlTU6fHZJ2uZJIecPC2BKUStlI3omUm6WSvH6VYWKtDUo2oRlgByVKmtoVlLTejms
KGpHL0S0LsKtUII9tIElYS/0FJiuX/c6sLWgJGzNR3Q5ndGlFb8P5Y2RyOniN7rbG8QOsdenuFHT
Y8h2e5g0s82TdFyz7YePIVEFD94mPZoftsZr1T9t0xmL7H+Z3dulSLDhplPOCYZTh1T8v3+UltgK
CM8XkIEVRoKDDVbEPlemudeAFG5DJIPidtJY+ETlLbkn3mLQxuZrPvC7FSU4HLYmbuEV99BUJIBp
f/q21KfYtM7BRh7FSNxpbVvpH4FPQqUxCDxemD1wGO4AV+q4Dw/Ug0q43Zb0xX7ID3cdbW6ZXEya
zrdKWgjzXlM/Gbz2p8BGUN9Sxd8iB8FD8NIioMj4L8en+NcQVy4mdA0H+Zno//xY/yLdN6w7bDMy
mr3z/V3XSXbZ7sHPu/obPGIMNDzs9Jz5BZo38jI1Y8UAe9yrBHZs6qZgTldbpw9JcuyJ7vd4HQjg
p6oz4ch4FFwwQhcgz7Zm+fzmHUrhGoeKO9ccSrcOl8WQG6NctiWV3D257iKRfCP1lADRav9t5ZQ7
zFX6DMQhO1Gr9/PoHqSFous+XVVfEunLzv2lJu4oErr4ah7X/nxp8e9BuIfNhkdtrKXcXViNmzUR
R4gvOYcwSE8/zv3ztg77RdivC+m6q3T4rxnRylmbgKTbWpbGi3GQk99nlmb9ZWIeUzS0IiWXoLx+
y97+qUDgwjMGVl22m79uRUvRwlwoEB1J/dzTcjBuSl9LHyRyXq5E1hUe50uhki/SS2+NRjoccZlr
2JsQLYsGYbhX1Wr4UP+oWtjXPvRHF2RdzceR/Hh/etZ9ziQA7mvD9kYNizuyu2hGrjvQgNWFaKtQ
uDawqTuB+d5o+M1R+f4agSdDWonnlRt3XLaheI0+pIix8P+GdmxESJtH8uDoIHN+V2/ffG2aumwn
raJ8iIZ/42NRf+03uxWV+0QoQYB0hnRwAyafGF1XOo4k8vCQ4S0ecTkMAK6brTjmxQ+lVY8hzWQ5
lC5OiuvbbM0f3v2FsFQQCPpDTuBDAzmfo4uhYLOqRZfnhRA2qwvMhpb01nedsLYwlxTD3G8MBsB7
vcmCWxwqnQZSkLCQL2Qc87W8iX398UGyQ/kV5zYq+Ho6j8mAnrfAybopW3XSdQ5Vn1NEvD/u35ms
NkRrMfvTaqwz2+g1tE5DEMgViQlBny8AMv0+pFEsKzSiBtG878Ab2PTOmxQo4SMfKDb1xt+CZLvZ
LBg8Bv7dFCUcAaQWXsj4+B2BDKFlKB6JCnYtMmZsjYeab4tP79XHBHX9t7BJMuR5QwA1RCNaiYv8
M4/4BUV3AGdPtlaSfC6oifqKfsKAgMjswwGcO9EZApbR89TS++A7ygJglgShkL7zJBJrSHdzRhQi
JKodB1Idrj2gPAZ/ZRX9t4NBSEHX5mwqDZk+MQpT0zY7qZjiy91uYYy3pUZw/gDZCyl1UKdkzVbY
SHlOu0vFrF9MSmJbZtCTALn6okblkeiVxfKiP0OAKysHLsCgSAjNyMdvUoYNgu8i9vQLKGMR4+vn
EZ1wRexN+eGBb44jywuVfcooJQFOC5rqzHbAjQ8f9g4WwyYbA+PLJtF9NVm6+dkw4ewm8WhuoQ6J
6y8sRgzQa2AHBux4lKufI+5SehTPGTXvwOr2KBs71GOLZYS9ceR44/QBXUqJyhjzoxhZhSgy6l6r
Gq9jZ91telcy0dpML5AL2G8FiQ6zwPk7SqjsncwPIeGRNS/mYm1uJj9UFgXfdtAM9ryiSaYt2L/2
4EbsT9Tktr5AQazjmyaeRlUpX+EirFQQloaaAlHcIxEzqoAvd++sq4ZadVZ2DBvirB+rKAkIRZu/
LlDrvMvl7YbB+pklTUFCSVD+/HXxQPQI+aofG33MlwZTI5KGzAArMbYZZkfPgZCwJhMS55NQ7nD2
oXMuE4J/VFkYVxcjGSWGBFCDDzu0YFv1XmIMM4tQe2kSnqf4aiC6B3EqHAQ54x45H/6DXhTR1nfu
6k7fxbLUaY6sK6Y8aipGPOyiOU955uxyAbpeO8sJ6szOfqeZXpxQSxci6JHIAtk746jR5/Hn2fFD
vZhmNhIDXYSUxBM5kqT3oCmIToQTPnA//nA6e9QslQKf9I2JP562fAcAqQb4yOXQa2mo6mYUZCgz
m7DtiOrV1sl3huOGTPl4osHTT8DijpA8Y2uWWbrXcABOXXZhfzAkoCeXXL5BkmU4kSc26JQeej4Y
ncDWxo5sD1tZhfkqocIo5GgV6xlcxqSwk+OHlXTwDW+4IC7y6Pr2FFJ3LqVHtSsgm6RAn7ExNkhv
0FkDO248EfOGSarGcov0RHtJtLUGtYnn35mQWNT1x1/2vmuVWkRQy/dlS945ZXPCPaGSCSsIyxW8
v1MIqZSJYoBtETX6orK5gxVFCXEjm40p6FGFn20voTAQWvfMyb0bdu2Xok4pwwzhaePEARuaF6Hh
PT7kc6NR4DUKrafO/qEeZ2rFVzIV/3cco9hQA3fxn5FYAzsWZw0968xtbX5Q9DupuwlUJ5I7j0EP
4c7hNGuhvsi6pr2Pz2INdM04WvoQd0hUhFj7TDRvqq6df3WADfLeN7BhpuCP6hobWJutmh6M6n92
6KhoxCtuP0nQD4oYPVsWalP0+Zi2/JxVE4vNmNu6theuWZxenETtdu1Sdw0FZJkEzNxgrGmNiAuf
MHvn5jfWTGHG2NQbwnLpSb6ONMd1Iu1qn/LtUsnnqDXjIg16dzkUYq4U+irISVQmHFC9hxC7SIqb
7DJW3lde07Ef7c0PdnfTF51uvNYpnF2WpMSIuw8AvkYIYa69o7U/IZgrCOPcHsosV2ua7Gbv3YnQ
ZaTy1KmynWHW4kKB5Vjl1b+93K2HYLWqHz+CCNn61Z0AIlL8X98D/u1tJN/PDWud1Ly45oB7V4ke
kGFns3RV5dbKg2CFLSJ4DPVzvt5j43qlgqOv+x/u/kyDUb9oHtsefcRo2K6Kx/PIp7GKxZWMDK6Q
tE4F5Va4EoXdE44FSjjw2VbPHh2vj4YPwokVKC/tNSZHgLx4ffHNbnSTfh71vQKH516L+2kgeNtj
JPH1278g64MXuirUAsEP6RIixMMXRK0l17C81yIMGXsYyWHvz4LWyGp00OpsEO+OmnZfw4CO2QKR
Iif354xJD/1baVyHKZ+G2Pxq7gcPRwEITJjGAlyNlGwOPtSTvPnAh+En89dgPwrVjirh9/EVm+Od
6+64RMtmXoi5Gx7HMK2HfgHbkh+EC2MC9KE5ndrJue30G4IxBmmaPGZRFWKDTR4WIsfr64rr9RCn
QwerBL7l9bs8Era6DaxrEnsnoOCR4eaW4gU3jvcNkB7ttjbJdT1N+oT4G6XdcH5/r2AwqfoPQU3G
RCzU1Fd4U5g6QOcj+mg27rl+OOEMpbky/v9n5fgq5TArEdSrL0irfte3qJSoz9W6fyVcOW7C+Odj
ADX3oW8PZlFiVIigtC0GKY+lOKDzP6/F+nLWbNISECe1AbKlYpHdMA7BDg2x6S1nFDTpBVObNL/R
rKDg9z9tkbloCJHPPBjSpRvCYhIhmEX81451nCR5Frh4AZfrzPU9DKYl5Dgt2N4VYFHGr4MCvGEj
lWQIsQq8KFyK00a3yIYoVRoQcnjgCNVyWPvap0zppLYmo+mg/N5tkIcOmHPPacf0cQWVDzbJFXYd
3HPQsjMpwQYI6RM3pSyyi5pLR6bPm/IsBseMqvkXIOlsuiqu7U9cnn48g6nYno9+XktvxiyjoJVV
DYnkPXydCfPyaLwldYF5tJHUs1KxwF7tFoeasMLxBF4ALVXy5gEk8PF1cp7hpGNK02eovOoNRBw5
JH7ijpfsRCAMPFhoO3isoNfRnG9OHBtPFT2hOF07RDEfAb4IkoFthrTTJKgKLqhR+84jJkI/Oi6D
sdH7Ym+EBdAO7ukbvQDcQUfUVENQ0jcaTNbuGBA4AVM05c1x9HQx6VObggByLrYeRvWpoNMJEcEz
BJbfRsLrLv1HXj3OSqmFZSvY0bKgEkoOiZGFd7a29HXNIbpxVMUGOupd4QaK9X+vdWfiFUs1MbqK
HFWEXaOf3RjSKR1YMq2Jvqb8QpRBXWoMtuA5tizdtXfHZKBfvDXsVX2iWjxVI04q4zaxeHZ+Df9Q
pqGzf/Taoe2LLFrQfGi2NQyD4U3PbClEBRQbSN4xCXytb8V5bYIK8XjfgpFReVQFhMRgCYcoSo3A
EvnywyYMO7GNAcGnAN11TEIe6MlGqY4cy545sB8JQCzmhtxl2xX+Bspndly6bjp/0jG04F1f0/7P
ZbKQlbhGcKlnZLjMeEhnRw2wNpumwW+PcYE2qOj3+hZV+qJQFpEZIykUP5xx7g1uLLN/cVn6x9W7
garz9JPkrXLyYyBVA2l7pG+bmdbP/giNwu9uNrolBm0kXa57cC+nJlyAWCQh12S3nU6Cl/11E86X
LEAR1HNozLJKU8tjSHZcUMZc4fAshRR3PQ0S5Xk9Nx6gTqzI3xLY4UZlXw6WG3dDcvB52Ia4L2NQ
IOjNjCzN8HMD0pkvrPVauzjzfwZmdqNtoFr4UkXbY3Bv6AEFsWAwCVxTNCgm0bhX37xmWcmv25uN
pyyvq65Y8YKTAvp8LIOjkC4j3FDuViJorJib4M8QiYG0Mp5MR/9/REAqTRR9Ovo7S7eEfwpq2W2o
hP9j3NrFIhwAgKw5ciZx2332ofk9P0MJStcrfDFiDmUdJ5uq4ZZ5EECkg4Xy8HeUOU8K/AYD8JGD
FScOYPKyqxyrEfAIW/Jby17Msq8lQE6vqylpJlz70SzPjHmWezh8JR+woCBttw00Dj7pd+08Vfrq
6zDTmm0b+oOV7OHKZgSfKMnRv9PwVnElaIAXFotb6vhw5MSaQIHEfgHnitpwRD0TNEYv+FQAuHoe
wntrSaqD2CvdF0rzENiCVp+JVbm7A4Kd49N4D9p4btGfUui9EKreLeu4OFN5ENieKY/+i28t7C/E
8Lecaf06Z+BGmG12DeKIb94zQpdbiujc7WtEUpFL/tk0UL9LXFa20FrFxVoAQccQ8WlZ/0W6t5H6
z0Ykl8EZbGImn367orWrZQKMm6ipiDunHx7iDmthPKfPkVfrfr0uPF5GWXQAcyQ0sjn3kygeGIUG
BuUuZ+ayDtDUf6XVewmtsTXXqXzKFD5secMmB3ZOuQk7q9bEs4saJNbMe2r6tj6rtFeSNRETqHtM
lhVdqkqdFPkf+UZop528i8FKRV2APmWL3qZ3f9F/t+nqcuosWldlSuCl5vO3h8k7nHwyOgeUpiw9
/51aD+tdiCazhyP4r59aBYY1l4Qetfw1XBiWtXaaUIczQ15+9KR+WczxW+ufY1DJ02e5dG8hNV4J
4L/oeGKf7IWuZrpAWQcOZBuloVQ8m5kShAFGE9L/SWOq5LfcX/fAi+NyUYQwEVMh6mdaNeyHkHeu
n5tjxzq6GuflPwkx2cNohKymOXlla8gMXnobDHO6WRnwHB6qWeloofb+OizL7rhS1aLnhOxUiud7
Xsm2DFCG680WUwfBLsPU5N2TMvREmxNFvuxhqV/ygwMZNM6Xgtsx6bAIOykPhuqzAGarFWxu9EgQ
hRujPdD90SDRUav3dSK0gF2Lduhn5mq8ZSudzyusDWSrVtN/LvZ8ULqF+uA45xBGGIDtUv6d/ptZ
YrfLXjn58cbceWkuIwQHKrGuWsLDrhKqDKhXVtlIuOwALSNznz0iG/9Ick4KQCJYwGIXS3YvE3Lh
wzsBM3hrI4zGvTS4z0iCFq4bJdHNdnljyTJEYtbJcndJejj3LOSm6zSdk4X8kzLxuUg97Lz/dqA4
pTjNgyotmzGyvrDiRgYNoU/MCdiKWwvZP5VeSwEJYyYRGsG6ub5CD/Q7CoXXD+y8bk4DwPAbKf0g
eRA4iKj57OZI+jpWFl5qvh2tdzyUvTNKNDFGhxjBxWgymr9CADmwLjQMJ83dXWlZ6gEELoUKSifG
GAiD0tzovTtquDbLAdTbNBETvPYHFuCcQ4CpsTRvfglx8pFZxrmcXqMZHAVLJhTXnYryOIcJb7gc
YL3fGMc351XhI5pF28NKi/RKzAKNeBkUMGWAu/2wOb3hsLrY0SbmVva3+GGDt6XOai3NqkjiieIx
xu1w43dOMNd1d3L8L6fyl6g4Q/Bl+HKoAW+YG4wUimP0B0I96uuJQDKocd7rWByVZL3JWxG3PZNh
vC9B4DMTP0HuGmyrjXqjtySjfMR43eFkam70Dm0+JfhycxzPLd0Fgt92lXRc/OrLG5tX0YezJQgY
Zgms4dKo2WJshagvzTF53cNxFj+VbOS2ndwgn1QXdEl84wBREdp6kz4=
`protect end_protected
